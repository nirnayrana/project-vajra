module riscv_pipeline_top (M_AXI_ARREADY,
    M_AXI_ARVALID,
    M_AXI_AWREADY,
    M_AXI_AWVALID,
    M_AXI_BREADY,
    M_AXI_BVALID,
    M_AXI_RREADY,
    M_AXI_RVALID,
    M_AXI_WREADY,
    M_AXI_WVALID,
    clk,
    rst_n,
    M_AXI_ARADDR,
    M_AXI_AWADDR,
    M_AXI_BRESP,
    M_AXI_RDATA,
    M_AXI_RRESP,
    M_AXI_WDATA,
    M_AXI_WSTRB,
    led);
 input M_AXI_ARREADY;
 output M_AXI_ARVALID;
 input M_AXI_AWREADY;
 output M_AXI_AWVALID;
 output M_AXI_BREADY;
 input M_AXI_BVALID;
 output M_AXI_RREADY;
 input M_AXI_RVALID;
 input M_AXI_WREADY;
 output M_AXI_WVALID;
 input clk;
 input rst_n;
 output [31:0] M_AXI_ARADDR;
 output [31:0] M_AXI_AWADDR;
 input [1:0] M_AXI_BRESP;
 input [31:0] M_AXI_RDATA;
 input [1:0] M_AXI_RRESP;
 output [31:0] M_AXI_WDATA;
 output [3:0] M_AXI_WSTRB;
 output [9:0] led;

 wire \AXI_BRIDGE.clk ;
 wire \AXI_BRIDGE.state[0] ;
 wire \AXI_BRIDGE.state[1] ;
 wire \AXI_BRIDGE.state[2] ;
 wire \AXI_BRIDGE.state[3] ;
 wire \AXI_BRIDGE.state[4] ;
 wire \AXI_BRIDGE.state[5] ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire \counter[0] ;
 wire \counter[10] ;
 wire \counter[11] ;
 wire \counter[12] ;
 wire \counter[13] ;
 wire \counter[14] ;
 wire \counter[15] ;
 wire \counter[16] ;
 wire \counter[17] ;
 wire \counter[18] ;
 wire \counter[19] ;
 wire \counter[1] ;
 wire \counter[20] ;
 wire \counter[21] ;
 wire \counter[22] ;
 wire \counter[23] ;
 wire \counter[24] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;

 sky130_fd_sc_hd__a221o_2 _093_ (.A1(M_AXI_BVALID),
    .A2(\AXI_BRIDGE.state[5] ),
    .B1(M_AXI_RVALID),
    .B2(\AXI_BRIDGE.state[4] ),
    .C1(\AXI_BRIDGE.state[0] ),
    .X(_002_));
 sky130_fd_sc_hd__and2b_2 _094_ (.A_N(M_AXI_WREADY),
    .B(\AXI_BRIDGE.state[2] ),
    .X(_079_));
 sky130_fd_sc_hd__a21o_2 _095_ (.A1(M_AXI_AWREADY),
    .A2(\AXI_BRIDGE.state[3] ),
    .B1(_079_),
    .X(_003_));
 sky130_fd_sc_hd__and2b_2 _096_ (.A_N(M_AXI_ARREADY),
    .B(\AXI_BRIDGE.state[1] ),
    .X(_080_));
 sky130_fd_sc_hd__buf_1 _097_ (.A(_080_),
    .X(_000_));
 sky130_fd_sc_hd__and2b_2 _098_ (.A_N(M_AXI_RVALID),
    .B(\AXI_BRIDGE.state[4] ),
    .X(_081_));
 sky130_fd_sc_hd__a21o_2 _099_ (.A1(\AXI_BRIDGE.state[1] ),
    .A2(M_AXI_ARREADY),
    .B1(_081_),
    .X(_004_));
 sky130_fd_sc_hd__inv_2 _100_ (.A(\AXI_BRIDGE.state[5] ),
    .Y(_082_));
 sky130_fd_sc_hd__nor2_2 _101_ (.A(M_AXI_BVALID),
    .B(_082_),
    .Y(_083_));
 sky130_fd_sc_hd__a21o_2 _102_ (.A1(\AXI_BRIDGE.state[2] ),
    .A2(M_AXI_WREADY),
    .B1(_083_),
    .X(_005_));
 sky130_fd_sc_hd__and2b_2 _103_ (.A_N(M_AXI_AWREADY),
    .B(\AXI_BRIDGE.state[3] ),
    .X(_084_));
 sky130_fd_sc_hd__buf_1 _104_ (.A(_084_),
    .X(_001_));
 sky130_fd_sc_hd__nand2_2 _105_ (.A(\counter[1] ),
    .B(\counter[0] ),
    .Y(_085_));
 sky130_fd_sc_hd__or2_2 _106_ (.A(\counter[1] ),
    .B(\counter[0] ),
    .X(_086_));
 sky130_fd_sc_hd__and2_2 _107_ (.A(_085_),
    .B(_086_),
    .X(_087_));
 sky130_fd_sc_hd__buf_1 _108_ (.A(_087_),
    .X(_017_));
 sky130_fd_sc_hd__xnor2_2 _109_ (.A(\counter[2] ),
    .B(_085_),
    .Y(_024_));
 sky130_fd_sc_hd__and4_2 _110_ (.A(\counter[1] ),
    .B(\counter[0] ),
    .C(\counter[2] ),
    .D(\counter[3] ),
    .X(_088_));
 sky130_fd_sc_hd__buf_1 _111_ (.A(_088_),
    .X(_089_));
 sky130_fd_sc_hd__a31o_2 _112_ (.A1(\counter[1] ),
    .A2(\counter[0] ),
    .A3(\counter[2] ),
    .B1(\counter[3] ),
    .X(_090_));
 sky130_fd_sc_hd__and2b_2 _113_ (.A_N(_089_),
    .B(_090_),
    .X(_091_));
 sky130_fd_sc_hd__buf_1 _114_ (.A(_091_),
    .X(_025_));
 sky130_fd_sc_hd__xor2_2 _115_ (.A(\counter[4] ),
    .B(_089_),
    .X(_026_));
 sky130_fd_sc_hd__nand3_2 _116_ (.A(\counter[4] ),
    .B(\counter[5] ),
    .C(_089_),
    .Y(_092_));
 sky130_fd_sc_hd__a21o_2 _117_ (.A1(\counter[4] ),
    .A2(_089_),
    .B1(\counter[5] ),
    .X(_035_));
 sky130_fd_sc_hd__and2_2 _118_ (.A(_092_),
    .B(_035_),
    .X(_036_));
 sky130_fd_sc_hd__buf_1 _119_ (.A(_036_),
    .X(_027_));
 sky130_fd_sc_hd__xnor2_2 _120_ (.A(\counter[6] ),
    .B(_092_),
    .Y(_028_));
 sky130_fd_sc_hd__a41o_2 _121_ (.A1(\counter[4] ),
    .A2(\counter[5] ),
    .A3(\counter[6] ),
    .A4(_089_),
    .B1(\counter[7] ),
    .X(_037_));
 sky130_fd_sc_hd__and4_2 _122_ (.A(\counter[4] ),
    .B(\counter[5] ),
    .C(\counter[6] ),
    .D(\counter[7] ),
    .X(_038_));
 sky130_fd_sc_hd__nand2_2 _123_ (.A(_089_),
    .B(_038_),
    .Y(_039_));
 sky130_fd_sc_hd__and2_2 _124_ (.A(_037_),
    .B(_039_),
    .X(_040_));
 sky130_fd_sc_hd__buf_1 _125_ (.A(_040_),
    .X(_029_));
 sky130_fd_sc_hd__xnor2_2 _126_ (.A(\counter[8] ),
    .B(_039_),
    .Y(_030_));
 sky130_fd_sc_hd__and2_2 _127_ (.A(_089_),
    .B(_038_),
    .X(_041_));
 sky130_fd_sc_hd__and3_2 _128_ (.A(\counter[8] ),
    .B(\counter[9] ),
    .C(_041_),
    .X(_042_));
 sky130_fd_sc_hd__a31o_2 _129_ (.A1(\counter[8] ),
    .A2(_089_),
    .A3(_038_),
    .B1(\counter[9] ),
    .X(_043_));
 sky130_fd_sc_hd__and2b_2 _130_ (.A_N(_042_),
    .B(_043_),
    .X(_044_));
 sky130_fd_sc_hd__buf_1 _131_ (.A(_044_),
    .X(_031_));
 sky130_fd_sc_hd__xor2_2 _132_ (.A(\counter[10] ),
    .B(_042_),
    .X(_007_));
 sky130_fd_sc_hd__and4_2 _133_ (.A(\counter[8] ),
    .B(\counter[9] ),
    .C(\counter[10] ),
    .D(_041_),
    .X(_045_));
 sky130_fd_sc_hd__and4_2 _134_ (.A(\counter[8] ),
    .B(\counter[9] ),
    .C(\counter[10] ),
    .D(\counter[11] ),
    .X(_046_));
 sky130_fd_sc_hd__and3_2 _135_ (.A(_089_),
    .B(_038_),
    .C(_046_),
    .X(_047_));
 sky130_fd_sc_hd__o21ba_2 _136_ (.A1(\counter[11] ),
    .A2(_045_),
    .B1_N(_047_),
    .X(_008_));
 sky130_fd_sc_hd__and2_2 _137_ (.A(\counter[12] ),
    .B(_047_),
    .X(_048_));
 sky130_fd_sc_hd__nor2_2 _138_ (.A(\counter[12] ),
    .B(_047_),
    .Y(_049_));
 sky130_fd_sc_hd__nor2_2 _139_ (.A(_048_),
    .B(_049_),
    .Y(_009_));
 sky130_fd_sc_hd__and3_2 _140_ (.A(\counter[12] ),
    .B(\counter[13] ),
    .C(_047_),
    .X(_050_));
 sky130_fd_sc_hd__o21ba_2 _141_ (.A1(\counter[13] ),
    .A2(_048_),
    .B1_N(_050_),
    .X(_010_));
 sky130_fd_sc_hd__xor2_2 _142_ (.A(\counter[14] ),
    .B(_050_),
    .X(_011_));
 sky130_fd_sc_hd__and4_2 _143_ (.A(\counter[12] ),
    .B(\counter[13] ),
    .C(\counter[14] ),
    .D(_047_),
    .X(_051_));
 sky130_fd_sc_hd__and4_2 _144_ (.A(\counter[12] ),
    .B(\counter[13] ),
    .C(\counter[14] ),
    .D(\counter[15] ),
    .X(_052_));
 sky130_fd_sc_hd__and4_2 _145_ (.A(_089_),
    .B(_038_),
    .C(_046_),
    .D(_052_),
    .X(_053_));
 sky130_fd_sc_hd__buf_1 _146_ (.A(_053_),
    .X(_054_));
 sky130_fd_sc_hd__o21ba_2 _147_ (.A1(\counter[15] ),
    .A2(_051_),
    .B1_N(_054_),
    .X(_012_));
 sky130_fd_sc_hd__xor2_2 _148_ (.A(\counter[16] ),
    .B(_054_),
    .X(_013_));
 sky130_fd_sc_hd__nand3_2 _149_ (.A(\counter[16] ),
    .B(\counter[17] ),
    .C(_054_),
    .Y(_055_));
 sky130_fd_sc_hd__a21o_2 _150_ (.A1(\counter[16] ),
    .A2(_054_),
    .B1(\counter[17] ),
    .X(_056_));
 sky130_fd_sc_hd__and2_2 _151_ (.A(_055_),
    .B(_056_),
    .X(_057_));
 sky130_fd_sc_hd__buf_1 _152_ (.A(_057_),
    .X(_014_));
 sky130_fd_sc_hd__xnor2_2 _153_ (.A(\counter[18] ),
    .B(_055_),
    .Y(_015_));
 sky130_fd_sc_hd__a41o_2 _154_ (.A1(\counter[16] ),
    .A2(\counter[17] ),
    .A3(\counter[18] ),
    .A4(_054_),
    .B1(\counter[19] ),
    .X(_058_));
 sky130_fd_sc_hd__and4_2 _155_ (.A(\counter[16] ),
    .B(\counter[17] ),
    .C(\counter[18] ),
    .D(\counter[19] ),
    .X(_059_));
 sky130_fd_sc_hd__nand2_2 _156_ (.A(_054_),
    .B(_059_),
    .Y(_060_));
 sky130_fd_sc_hd__and2_2 _157_ (.A(_058_),
    .B(_060_),
    .X(_061_));
 sky130_fd_sc_hd__buf_1 _158_ (.A(_061_),
    .X(_016_));
 sky130_fd_sc_hd__xnor2_2 _159_ (.A(\counter[20] ),
    .B(_060_),
    .Y(_018_));
 sky130_fd_sc_hd__and2_2 _160_ (.A(\counter[20] ),
    .B(\counter[21] ),
    .X(_062_));
 sky130_fd_sc_hd__and3_2 _161_ (.A(_054_),
    .B(_059_),
    .C(_062_),
    .X(_063_));
 sky130_fd_sc_hd__a31o_2 _162_ (.A1(\counter[20] ),
    .A2(_054_),
    .A3(_059_),
    .B1(\counter[21] ),
    .X(_064_));
 sky130_fd_sc_hd__and2b_2 _163_ (.A_N(_063_),
    .B(_064_),
    .X(_065_));
 sky130_fd_sc_hd__buf_1 _164_ (.A(_065_),
    .X(_019_));
 sky130_fd_sc_hd__xor2_2 _165_ (.A(\counter[22] ),
    .B(_063_),
    .X(_020_));
 sky130_fd_sc_hd__and3_2 _166_ (.A(\counter[22] ),
    .B(\counter[23] ),
    .C(_062_),
    .X(_066_));
 sky130_fd_sc_hd__and3_2 _167_ (.A(_053_),
    .B(_059_),
    .C(_066_),
    .X(_067_));
 sky130_fd_sc_hd__a41o_2 _168_ (.A1(\counter[22] ),
    .A2(_054_),
    .A3(_059_),
    .A4(_062_),
    .B1(\counter[23] ),
    .X(_068_));
 sky130_fd_sc_hd__and2b_2 _169_ (.A_N(_067_),
    .B(_068_),
    .X(_069_));
 sky130_fd_sc_hd__buf_1 _170_ (.A(_069_),
    .X(_021_));
 sky130_fd_sc_hd__xor2_2 _171_ (.A(\counter[24] ),
    .B(_067_),
    .X(_022_));
 sky130_fd_sc_hd__and4_2 _172_ (.A(\counter[24] ),
    .B(_054_),
    .C(_059_),
    .D(_066_),
    .X(_070_));
 sky130_fd_sc_hd__xor2_2 _173_ (.A(\AXI_BRIDGE.clk ),
    .B(_070_),
    .X(_023_));
 sky130_fd_sc_hd__inv_2 _174_ (.A(\counter[0] ),
    .Y(_006_));
 sky130_fd_sc_hd__inv_2 _175_ (.A(_081_),
    .Y(_071_));
 sky130_fd_sc_hd__or3_2 _176_ (.A(\AXI_BRIDGE.state[0] ),
    .B(\AXI_BRIDGE.state[4] ),
    .C(\AXI_BRIDGE.state[1] ),
    .X(_072_));
 sky130_fd_sc_hd__or3b_2 _177_ (.A(_000_),
    .B(_081_),
    .C_N(_072_),
    .X(_073_));
 sky130_fd_sc_hd__a32o_2 _178_ (.A1(\AXI_BRIDGE.state[1] ),
    .A2(M_AXI_ARREADY),
    .A3(_071_),
    .B1(_073_),
    .B2(M_AXI_RREADY),
    .X(_032_));
 sky130_fd_sc_hd__inv_2 _179_ (.A(_083_),
    .Y(_074_));
 sky130_fd_sc_hd__nor2_2 _180_ (.A(\AXI_BRIDGE.state[0] ),
    .B(\AXI_BRIDGE.state[2] ),
    .Y(_075_));
 sky130_fd_sc_hd__a211o_2 _181_ (.A1(_082_),
    .A2(_075_),
    .B1(_083_),
    .C1(_079_),
    .X(_076_));
 sky130_fd_sc_hd__a32o_2 _182_ (.A1(\AXI_BRIDGE.state[2] ),
    .A2(M_AXI_WREADY),
    .A3(_074_),
    .B1(_076_),
    .B2(M_AXI_BREADY),
    .X(_033_));
 sky130_fd_sc_hd__inv_2 _183_ (.A(_079_),
    .Y(_077_));
 sky130_fd_sc_hd__o31a_2 _184_ (.A1(_079_),
    .A2(_001_),
    .A3(_075_),
    .B1(M_AXI_WVALID),
    .X(_078_));
 sky130_fd_sc_hd__a31o_2 _185_ (.A1(M_AXI_AWREADY),
    .A2(\AXI_BRIDGE.state[3] ),
    .A3(_077_),
    .B1(_078_),
    .X(_034_));
 sky130_fd_sc_hd__dfrtp_2 _186_ (.CLK(clk),
    .D(_006_),
    .RESET_B(rst_n),
    .Q(\counter[0] ));
 sky130_fd_sc_hd__dfrtp_2 _187_ (.CLK(clk),
    .D(_017_),
    .RESET_B(rst_n),
    .Q(\counter[1] ));
 sky130_fd_sc_hd__dfrtp_2 _188_ (.CLK(clk),
    .D(_024_),
    .RESET_B(rst_n),
    .Q(\counter[2] ));
 sky130_fd_sc_hd__dfrtp_2 _189_ (.CLK(clk),
    .D(_025_),
    .RESET_B(rst_n),
    .Q(\counter[3] ));
 sky130_fd_sc_hd__dfrtp_2 _190_ (.CLK(clk),
    .D(_026_),
    .RESET_B(rst_n),
    .Q(\counter[4] ));
 sky130_fd_sc_hd__dfrtp_2 _191_ (.CLK(clk),
    .D(_027_),
    .RESET_B(rst_n),
    .Q(\counter[5] ));
 sky130_fd_sc_hd__dfrtp_2 _192_ (.CLK(clk),
    .D(_028_),
    .RESET_B(rst_n),
    .Q(\counter[6] ));
 sky130_fd_sc_hd__dfrtp_2 _193_ (.CLK(clk),
    .D(_029_),
    .RESET_B(rst_n),
    .Q(\counter[7] ));
 sky130_fd_sc_hd__dfrtp_2 _194_ (.CLK(clk),
    .D(_030_),
    .RESET_B(rst_n),
    .Q(\counter[8] ));
 sky130_fd_sc_hd__dfrtp_2 _195_ (.CLK(clk),
    .D(_031_),
    .RESET_B(rst_n),
    .Q(\counter[9] ));
 sky130_fd_sc_hd__dfrtp_2 _196_ (.CLK(clk),
    .D(_007_),
    .RESET_B(rst_n),
    .Q(\counter[10] ));
 sky130_fd_sc_hd__dfrtp_2 _197_ (.CLK(clk),
    .D(_008_),
    .RESET_B(rst_n),
    .Q(\counter[11] ));
 sky130_fd_sc_hd__dfrtp_2 _198_ (.CLK(clk),
    .D(_009_),
    .RESET_B(rst_n),
    .Q(\counter[12] ));
 sky130_fd_sc_hd__dfrtp_2 _199_ (.CLK(clk),
    .D(_010_),
    .RESET_B(rst_n),
    .Q(\counter[13] ));
 sky130_fd_sc_hd__dfrtp_2 _200_ (.CLK(clk),
    .D(_011_),
    .RESET_B(rst_n),
    .Q(\counter[14] ));
 sky130_fd_sc_hd__dfrtp_2 _201_ (.CLK(clk),
    .D(_012_),
    .RESET_B(rst_n),
    .Q(\counter[15] ));
 sky130_fd_sc_hd__dfrtp_2 _202_ (.CLK(clk),
    .D(_013_),
    .RESET_B(rst_n),
    .Q(\counter[16] ));
 sky130_fd_sc_hd__dfrtp_2 _203_ (.CLK(clk),
    .D(_014_),
    .RESET_B(rst_n),
    .Q(\counter[17] ));
 sky130_fd_sc_hd__dfrtp_2 _204_ (.CLK(clk),
    .D(_015_),
    .RESET_B(rst_n),
    .Q(\counter[18] ));
 sky130_fd_sc_hd__dfrtp_2 _205_ (.CLK(clk),
    .D(_016_),
    .RESET_B(rst_n),
    .Q(\counter[19] ));
 sky130_fd_sc_hd__dfrtp_2 _206_ (.CLK(clk),
    .D(_018_),
    .RESET_B(rst_n),
    .Q(\counter[20] ));
 sky130_fd_sc_hd__dfrtp_2 _207_ (.CLK(clk),
    .D(_019_),
    .RESET_B(rst_n),
    .Q(\counter[21] ));
 sky130_fd_sc_hd__dfrtp_2 _208_ (.CLK(clk),
    .D(_020_),
    .RESET_B(rst_n),
    .Q(\counter[22] ));
 sky130_fd_sc_hd__dfrtp_2 _209_ (.CLK(clk),
    .D(_021_),
    .RESET_B(rst_n),
    .Q(\counter[23] ));
 sky130_fd_sc_hd__dfrtp_2 _210_ (.CLK(clk),
    .D(_022_),
    .RESET_B(rst_n),
    .Q(\counter[24] ));
 sky130_fd_sc_hd__dfrtp_2 _211_ (.CLK(clk),
    .D(_023_),
    .RESET_B(rst_n),
    .Q(\AXI_BRIDGE.clk ));
 sky130_fd_sc_hd__dfstp_2 _212_ (.CLK(\AXI_BRIDGE.clk ),
    .D(_002_),
    .SET_B(rst_n),
    .Q(\AXI_BRIDGE.state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _213_ (.CLK(\AXI_BRIDGE.clk ),
    .D(_000_),
    .RESET_B(rst_n),
    .Q(\AXI_BRIDGE.state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _214_ (.CLK(\AXI_BRIDGE.clk ),
    .D(_003_),
    .RESET_B(rst_n),
    .Q(\AXI_BRIDGE.state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _215_ (.CLK(\AXI_BRIDGE.clk ),
    .D(_001_),
    .RESET_B(rst_n),
    .Q(\AXI_BRIDGE.state[3] ));
 sky130_fd_sc_hd__dfrtp_2 _216_ (.CLK(\AXI_BRIDGE.clk ),
    .D(_004_),
    .RESET_B(rst_n),
    .Q(\AXI_BRIDGE.state[4] ));
 sky130_fd_sc_hd__dfrtp_2 _217_ (.CLK(\AXI_BRIDGE.clk ),
    .D(_005_),
    .RESET_B(rst_n),
    .Q(\AXI_BRIDGE.state[5] ));
 sky130_fd_sc_hd__dfrtp_2 _218_ (.CLK(\AXI_BRIDGE.clk ),
    .D(_032_),
    .RESET_B(rst_n),
    .Q(M_AXI_RREADY));
 sky130_fd_sc_hd__dfrtp_2 _219_ (.CLK(\AXI_BRIDGE.clk ),
    .D(_033_),
    .RESET_B(rst_n),
    .Q(M_AXI_BREADY));
 sky130_fd_sc_hd__dfrtp_2 _220_ (.CLK(\AXI_BRIDGE.clk ),
    .D(_034_),
    .RESET_B(rst_n),
    .Q(M_AXI_WVALID));
 sky130_fd_sc_hd__conb_1 _221_ (.HI(M_AXI_WSTRB[0]));
 sky130_fd_sc_hd__conb_1 _222_ (.LO(M_AXI_ARADDR[0]));
 sky130_fd_sc_hd__conb_1 _223_ (.LO(M_AXI_ARADDR[1]));
 sky130_fd_sc_hd__conb_1 _224_ (.LO(M_AXI_ARADDR[2]));
 sky130_fd_sc_hd__conb_1 _225_ (.LO(M_AXI_ARADDR[3]));
 sky130_fd_sc_hd__conb_1 _226_ (.LO(M_AXI_ARADDR[4]));
 sky130_fd_sc_hd__conb_1 _227_ (.LO(M_AXI_ARADDR[5]));
 sky130_fd_sc_hd__conb_1 _228_ (.LO(M_AXI_ARADDR[6]));
 sky130_fd_sc_hd__conb_1 _229_ (.LO(M_AXI_ARADDR[7]));
 sky130_fd_sc_hd__conb_1 _230_ (.LO(M_AXI_ARADDR[8]));
 sky130_fd_sc_hd__conb_1 _231_ (.LO(M_AXI_ARADDR[9]));
 sky130_fd_sc_hd__conb_1 _232_ (.LO(M_AXI_ARADDR[10]));
 sky130_fd_sc_hd__conb_1 _233_ (.LO(M_AXI_ARADDR[11]));
 sky130_fd_sc_hd__conb_1 _234_ (.LO(M_AXI_ARADDR[12]));
 sky130_fd_sc_hd__conb_1 _235_ (.LO(M_AXI_ARADDR[13]));
 sky130_fd_sc_hd__conb_1 _236_ (.LO(M_AXI_ARADDR[14]));
 sky130_fd_sc_hd__conb_1 _237_ (.LO(M_AXI_ARADDR[15]));
 sky130_fd_sc_hd__conb_1 _238_ (.LO(M_AXI_ARADDR[16]));
 sky130_fd_sc_hd__conb_1 _239_ (.LO(M_AXI_ARADDR[17]));
 sky130_fd_sc_hd__conb_1 _240_ (.LO(M_AXI_ARADDR[18]));
 sky130_fd_sc_hd__conb_1 _241_ (.LO(M_AXI_ARADDR[19]));
 sky130_fd_sc_hd__conb_1 _242_ (.LO(M_AXI_ARADDR[20]));
 sky130_fd_sc_hd__conb_1 _243_ (.LO(M_AXI_ARADDR[21]));
 sky130_fd_sc_hd__conb_1 _244_ (.LO(M_AXI_ARADDR[22]));
 sky130_fd_sc_hd__conb_1 _245_ (.LO(M_AXI_ARADDR[23]));
 sky130_fd_sc_hd__conb_1 _246_ (.LO(M_AXI_ARADDR[24]));
 sky130_fd_sc_hd__conb_1 _247_ (.LO(M_AXI_ARADDR[25]));
 sky130_fd_sc_hd__conb_1 _248_ (.LO(M_AXI_ARADDR[26]));
 sky130_fd_sc_hd__conb_1 _249_ (.LO(M_AXI_ARADDR[27]));
 sky130_fd_sc_hd__conb_1 _250_ (.LO(M_AXI_ARADDR[28]));
 sky130_fd_sc_hd__conb_1 _251_ (.LO(M_AXI_ARADDR[29]));
 sky130_fd_sc_hd__conb_1 _252_ (.LO(M_AXI_ARADDR[30]));
 sky130_fd_sc_hd__conb_1 _253_ (.LO(M_AXI_ARADDR[31]));
 sky130_fd_sc_hd__conb_1 _254_ (.LO(M_AXI_ARVALID));
 sky130_fd_sc_hd__conb_1 _255_ (.LO(M_AXI_AWADDR[0]));
 sky130_fd_sc_hd__conb_1 _256_ (.LO(M_AXI_AWADDR[1]));
 sky130_fd_sc_hd__conb_1 _257_ (.LO(M_AXI_AWADDR[2]));
 sky130_fd_sc_hd__conb_1 _258_ (.LO(M_AXI_AWADDR[3]));
 sky130_fd_sc_hd__conb_1 _259_ (.LO(M_AXI_AWADDR[4]));
 sky130_fd_sc_hd__conb_1 _260_ (.LO(M_AXI_AWADDR[5]));
 sky130_fd_sc_hd__conb_1 _261_ (.LO(M_AXI_AWADDR[6]));
 sky130_fd_sc_hd__conb_1 _262_ (.LO(M_AXI_AWADDR[7]));
 sky130_fd_sc_hd__conb_1 _263_ (.LO(M_AXI_AWADDR[8]));
 sky130_fd_sc_hd__conb_1 _264_ (.LO(M_AXI_AWADDR[9]));
 sky130_fd_sc_hd__conb_1 _265_ (.LO(M_AXI_AWADDR[10]));
 sky130_fd_sc_hd__conb_1 _266_ (.LO(M_AXI_AWADDR[11]));
 sky130_fd_sc_hd__conb_1 _267_ (.LO(M_AXI_AWADDR[12]));
 sky130_fd_sc_hd__conb_1 _268_ (.LO(M_AXI_AWADDR[13]));
 sky130_fd_sc_hd__conb_1 _269_ (.LO(M_AXI_AWADDR[14]));
 sky130_fd_sc_hd__conb_1 _270_ (.LO(M_AXI_AWADDR[15]));
 sky130_fd_sc_hd__conb_1 _271_ (.LO(M_AXI_AWADDR[16]));
 sky130_fd_sc_hd__conb_1 _272_ (.LO(M_AXI_AWADDR[17]));
 sky130_fd_sc_hd__conb_1 _273_ (.LO(M_AXI_AWADDR[18]));
 sky130_fd_sc_hd__conb_1 _274_ (.LO(M_AXI_AWADDR[19]));
 sky130_fd_sc_hd__conb_1 _275_ (.LO(M_AXI_AWADDR[20]));
 sky130_fd_sc_hd__conb_1 _276_ (.LO(M_AXI_AWADDR[21]));
 sky130_fd_sc_hd__conb_1 _277_ (.LO(M_AXI_AWADDR[22]));
 sky130_fd_sc_hd__conb_1 _278_ (.LO(M_AXI_AWADDR[23]));
 sky130_fd_sc_hd__conb_1 _279_ (.LO(M_AXI_AWADDR[24]));
 sky130_fd_sc_hd__conb_1 _280_ (.LO(M_AXI_AWADDR[25]));
 sky130_fd_sc_hd__conb_1 _281_ (.LO(M_AXI_AWADDR[26]));
 sky130_fd_sc_hd__conb_1 _282_ (.LO(M_AXI_AWADDR[27]));
 sky130_fd_sc_hd__conb_1 _283_ (.LO(M_AXI_AWADDR[28]));
 sky130_fd_sc_hd__conb_1 _284_ (.LO(M_AXI_AWADDR[29]));
 sky130_fd_sc_hd__conb_1 _285_ (.LO(M_AXI_AWADDR[30]));
 sky130_fd_sc_hd__conb_1 _286_ (.LO(M_AXI_AWADDR[31]));
 sky130_fd_sc_hd__conb_1 _287_ (.LO(M_AXI_AWVALID));
 sky130_fd_sc_hd__conb_1 _288_ (.LO(M_AXI_WDATA[0]));
 sky130_fd_sc_hd__conb_1 _289_ (.LO(M_AXI_WDATA[1]));
 sky130_fd_sc_hd__conb_1 _290_ (.LO(M_AXI_WDATA[2]));
 sky130_fd_sc_hd__conb_1 _291_ (.LO(M_AXI_WDATA[3]));
 sky130_fd_sc_hd__conb_1 _292_ (.LO(M_AXI_WDATA[4]));
 sky130_fd_sc_hd__conb_1 _293_ (.LO(M_AXI_WDATA[5]));
 sky130_fd_sc_hd__conb_1 _294_ (.LO(M_AXI_WDATA[6]));
 sky130_fd_sc_hd__conb_1 _295_ (.LO(M_AXI_WDATA[7]));
 sky130_fd_sc_hd__conb_1 _296_ (.LO(M_AXI_WDATA[8]));
 sky130_fd_sc_hd__conb_1 _297_ (.LO(M_AXI_WDATA[9]));
 sky130_fd_sc_hd__conb_1 _298_ (.LO(M_AXI_WDATA[10]));
 sky130_fd_sc_hd__conb_1 _299_ (.LO(M_AXI_WDATA[11]));
 sky130_fd_sc_hd__conb_1 _300_ (.LO(M_AXI_WDATA[12]));
 sky130_fd_sc_hd__conb_1 _301_ (.LO(M_AXI_WDATA[13]));
 sky130_fd_sc_hd__conb_1 _302_ (.LO(M_AXI_WDATA[14]));
 sky130_fd_sc_hd__conb_1 _303_ (.LO(M_AXI_WDATA[15]));
 sky130_fd_sc_hd__conb_1 _304_ (.LO(M_AXI_WDATA[16]));
 sky130_fd_sc_hd__conb_1 _305_ (.LO(M_AXI_WDATA[17]));
 sky130_fd_sc_hd__conb_1 _306_ (.LO(M_AXI_WDATA[18]));
 sky130_fd_sc_hd__conb_1 _307_ (.LO(M_AXI_WDATA[19]));
 sky130_fd_sc_hd__conb_1 _308_ (.LO(M_AXI_WDATA[20]));
 sky130_fd_sc_hd__conb_1 _309_ (.LO(M_AXI_WDATA[21]));
 sky130_fd_sc_hd__conb_1 _310_ (.LO(M_AXI_WDATA[22]));
 sky130_fd_sc_hd__conb_1 _311_ (.LO(M_AXI_WDATA[23]));
 sky130_fd_sc_hd__conb_1 _312_ (.LO(M_AXI_WDATA[24]));
 sky130_fd_sc_hd__conb_1 _313_ (.LO(M_AXI_WDATA[25]));
 sky130_fd_sc_hd__conb_1 _314_ (.LO(M_AXI_WDATA[26]));
 sky130_fd_sc_hd__conb_1 _315_ (.LO(M_AXI_WDATA[27]));
 sky130_fd_sc_hd__conb_1 _316_ (.LO(M_AXI_WDATA[28]));
 sky130_fd_sc_hd__conb_1 _317_ (.LO(M_AXI_WDATA[29]));
 sky130_fd_sc_hd__conb_1 _318_ (.LO(M_AXI_WDATA[30]));
 sky130_fd_sc_hd__conb_1 _319_ (.LO(M_AXI_WDATA[31]));
 sky130_fd_sc_hd__conb_1 _320_ (.LO(M_AXI_WSTRB[1]));
 sky130_fd_sc_hd__conb_1 _321_ (.LO(M_AXI_WSTRB[2]));
 sky130_fd_sc_hd__conb_1 _322_ (.LO(M_AXI_WSTRB[3]));
 sky130_fd_sc_hd__conb_1 _323_ (.LO(led[0]));
 sky130_fd_sc_hd__conb_1 _324_ (.LO(led[1]));
 sky130_fd_sc_hd__conb_1 _325_ (.LO(led[2]));
 sky130_fd_sc_hd__conb_1 _326_ (.LO(led[3]));
 sky130_fd_sc_hd__conb_1 _327_ (.LO(led[4]));
 sky130_fd_sc_hd__conb_1 _328_ (.LO(led[5]));
 sky130_fd_sc_hd__conb_1 _329_ (.LO(led[6]));
 sky130_fd_sc_hd__conb_1 _330_ (.LO(led[7]));
 sky130_fd_sc_hd__conb_1 _331_ (.LO(led[8]));
 sky130_fd_sc_hd__conb_1 _332_ (.LO(led[9]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
endmodule
