VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO riscv_pipeline_top
  CLASS BLOCK ;
  FOREIGN riscv_pipeline_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN M_AXI_ARADDR[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 496.000 180.690 500.000 ;
    END
  END M_AXI_ARADDR[0]
  PIN M_AXI_ARADDR[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 496.000 216.110 500.000 ;
    END
  END M_AXI_ARADDR[10]
  PIN M_AXI_ARADDR[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END M_AXI_ARADDR[11]
  PIN M_AXI_ARADDR[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 353.640 500.000 354.240 ;
    END
  END M_AXI_ARADDR[12]
  PIN M_AXI_ARADDR[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END M_AXI_ARADDR[13]
  PIN M_AXI_ARADDR[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 445.440 500.000 446.040 ;
    END
  END M_AXI_ARADDR[14]
  PIN M_AXI_ARADDR[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END M_AXI_ARADDR[15]
  PIN M_AXI_ARADDR[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 496.000 67.990 500.000 ;
    END
  END M_AXI_ARADDR[16]
  PIN M_AXI_ARADDR[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 496.000 303.050 500.000 ;
    END
  END M_AXI_ARADDR[17]
  PIN M_AXI_ARADDR[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 173.440 500.000 174.040 ;
    END
  END M_AXI_ARADDR[18]
  PIN M_AXI_ARADDR[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 418.240 500.000 418.840 ;
    END
  END M_AXI_ARADDR[19]
  PIN M_AXI_ARADDR[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 210.840 500.000 211.440 ;
    END
  END M_AXI_ARADDR[1]
  PIN M_AXI_ARADDR[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 261.840 500.000 262.440 ;
    END
  END M_AXI_ARADDR[20]
  PIN M_AXI_ARADDR[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END M_AXI_ARADDR[21]
  PIN M_AXI_ARADDR[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 340.040 500.000 340.640 ;
    END
  END M_AXI_ARADDR[22]
  PIN M_AXI_ARADDR[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 496.000 315.930 500.000 ;
    END
  END M_AXI_ARADDR[23]
  PIN M_AXI_ARADDR[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 496.000 328.810 500.000 ;
    END
  END M_AXI_ARADDR[24]
  PIN M_AXI_ARADDR[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 496.000 193.570 500.000 ;
    END
  END M_AXI_ARADDR[25]
  PIN M_AXI_ARADDR[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END M_AXI_ARADDR[26]
  PIN M_AXI_ARADDR[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END M_AXI_ARADDR[27]
  PIN M_AXI_ARADDR[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END M_AXI_ARADDR[28]
  PIN M_AXI_ARADDR[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END M_AXI_ARADDR[29]
  PIN M_AXI_ARADDR[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END M_AXI_ARADDR[2]
  PIN M_AXI_ARADDR[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END M_AXI_ARADDR[30]
  PIN M_AXI_ARADDR[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END M_AXI_ARADDR[31]
  PIN M_AXI_ARADDR[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END M_AXI_ARADDR[3]
  PIN M_AXI_ARADDR[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END M_AXI_ARADDR[4]
  PIN M_AXI_ARADDR[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 132.640 500.000 133.240 ;
    END
  END M_AXI_ARADDR[5]
  PIN M_AXI_ARADDR[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END M_AXI_ARADDR[6]
  PIN M_AXI_ARADDR[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 183.640 500.000 184.240 ;
    END
  END M_AXI_ARADDR[7]
  PIN M_AXI_ARADDR[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 105.440 500.000 106.040 ;
    END
  END M_AXI_ARADDR[8]
  PIN M_AXI_ARADDR[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END M_AXI_ARADDR[9]
  PIN M_AXI_ARREADY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 489.530 496.000 489.810 500.000 ;
    END
  END M_AXI_ARREADY
  PIN M_AXI_ARVALID
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END M_AXI_ARVALID
  PIN M_AXI_AWADDR[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 367.240 500.000 367.840 ;
    END
  END M_AXI_AWADDR[0]
  PIN M_AXI_AWADDR[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 472.640 500.000 473.240 ;
    END
  END M_AXI_AWADDR[10]
  PIN M_AXI_AWADDR[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 302.640 500.000 303.240 ;
    END
  END M_AXI_AWADDR[11]
  PIN M_AXI_AWADDR[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END M_AXI_AWADDR[12]
  PIN M_AXI_AWADDR[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END M_AXI_AWADDR[13]
  PIN M_AXI_AWADDR[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 431.840 500.000 432.440 ;
    END
  END M_AXI_AWADDR[14]
  PIN M_AXI_AWADDR[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END M_AXI_AWADDR[15]
  PIN M_AXI_AWADDR[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 224.440 500.000 225.040 ;
    END
  END M_AXI_AWADDR[16]
  PIN M_AXI_AWADDR[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END M_AXI_AWADDR[17]
  PIN M_AXI_AWADDR[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 496.000 451.170 500.000 ;
    END
  END M_AXI_AWADDR[18]
  PIN M_AXI_AWADDR[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END M_AXI_AWADDR[19]
  PIN M_AXI_AWADDR[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END M_AXI_AWADDR[1]
  PIN M_AXI_AWADDR[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END M_AXI_AWADDR[20]
  PIN M_AXI_AWADDR[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 40.840 500.000 41.440 ;
    END
  END M_AXI_AWADDR[21]
  PIN M_AXI_AWADDR[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 496.000 499.470 500.000 ;
    END
  END M_AXI_AWADDR[22]
  PIN M_AXI_AWADDR[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END M_AXI_AWADDR[23]
  PIN M_AXI_AWADDR[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 496.000 241.870 500.000 ;
    END
  END M_AXI_AWADDR[24]
  PIN M_AXI_AWADDR[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END M_AXI_AWADDR[25]
  PIN M_AXI_AWADDR[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 496.000 351.350 500.000 ;
    END
  END M_AXI_AWADDR[26]
  PIN M_AXI_AWADDR[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 496.000 167.810 500.000 ;
    END
  END M_AXI_AWADDR[27]
  PIN M_AXI_AWADDR[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END M_AXI_AWADDR[28]
  PIN M_AXI_AWADDR[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 27.240 500.000 27.840 ;
    END
  END M_AXI_AWADDR[29]
  PIN M_AXI_AWADDR[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 95.240 500.000 95.840 ;
    END
  END M_AXI_AWADDR[2]
  PIN M_AXI_AWADDR[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 496.000 476.930 500.000 ;
    END
  END M_AXI_AWADDR[30]
  PIN M_AXI_AWADDR[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 496.000 154.930 500.000 ;
    END
  END M_AXI_AWADDR[31]
  PIN M_AXI_AWADDR[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END M_AXI_AWADDR[3]
  PIN M_AXI_AWADDR[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END M_AXI_AWADDR[4]
  PIN M_AXI_AWADDR[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 289.040 500.000 289.640 ;
    END
  END M_AXI_AWADDR[5]
  PIN M_AXI_AWADDR[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END M_AXI_AWADDR[6]
  PIN M_AXI_AWADDR[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 496.000 377.110 500.000 ;
    END
  END M_AXI_AWADDR[7]
  PIN M_AXI_AWADDR[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 380.840 500.000 381.440 ;
    END
  END M_AXI_AWADDR[8]
  PIN M_AXI_AWADDR[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END M_AXI_AWADDR[9]
  PIN M_AXI_AWREADY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 389.710 496.000 389.990 500.000 ;
    END
  END M_AXI_AWREADY
  PIN M_AXI_AWVALID
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 54.440 500.000 55.040 ;
    END
  END M_AXI_AWVALID
  PIN M_AXI_BREADY
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 32.290 496.000 32.570 500.000 ;
    END
  END M_AXI_BREADY
  PIN M_AXI_BRESP[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END M_AXI_BRESP[0]
  PIN M_AXI_BRESP[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END M_AXI_BRESP[1]
  PIN M_AXI_BVALID
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 289.890 496.000 290.170 500.000 ;
    END
  END M_AXI_BVALID
  PIN M_AXI_RDATA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END M_AXI_RDATA[0]
  PIN M_AXI_RDATA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END M_AXI_RDATA[10]
  PIN M_AXI_RDATA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 496.000 19.690 500.000 ;
    END
  END M_AXI_RDATA[11]
  PIN M_AXI_RDATA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END M_AXI_RDATA[12]
  PIN M_AXI_RDATA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 496.000 45.450 500.000 ;
    END
  END M_AXI_RDATA[13]
  PIN M_AXI_RDATA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 496.000 142.050 500.000 ;
    END
  END M_AXI_RDATA[14]
  PIN M_AXI_RDATA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 496.000 203.230 500.000 ;
    END
  END M_AXI_RDATA[15]
  PIN M_AXI_RDATA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END M_AXI_RDATA[16]
  PIN M_AXI_RDATA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 496.000 464.050 500.000 ;
    END
  END M_AXI_RDATA[17]
  PIN M_AXI_RDATA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 197.240 500.000 197.840 ;
    END
  END M_AXI_RDATA[18]
  PIN M_AXI_RDATA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END M_AXI_RDATA[19]
  PIN M_AXI_RDATA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END M_AXI_RDATA[1]
  PIN M_AXI_RDATA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 496.000 341.690 500.000 ;
    END
  END M_AXI_RDATA[20]
  PIN M_AXI_RDATA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END M_AXI_RDATA[21]
  PIN M_AXI_RDATA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 496.000 80.870 500.000 ;
    END
  END M_AXI_RDATA[22]
  PIN M_AXI_RDATA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 394.440 500.000 395.040 ;
    END
  END M_AXI_RDATA[23]
  PIN M_AXI_RDATA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 496.000 129.170 500.000 ;
    END
  END M_AXI_RDATA[24]
  PIN M_AXI_RDATA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 496.000 415.750 500.000 ;
    END
  END M_AXI_RDATA[25]
  PIN M_AXI_RDATA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 496.000 267.630 500.000 ;
    END
  END M_AXI_RDATA[26]
  PIN M_AXI_RDATA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 496.000 402.870 500.000 ;
    END
  END M_AXI_RDATA[27]
  PIN M_AXI_RDATA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END M_AXI_RDATA[28]
  PIN M_AXI_RDATA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END M_AXI_RDATA[29]
  PIN M_AXI_RDATA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 17.040 500.000 17.640 ;
    END
  END M_AXI_RDATA[2]
  PIN M_AXI_RDATA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 496.000 55.110 500.000 ;
    END
  END M_AXI_RDATA[30]
  PIN M_AXI_RDATA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END M_AXI_RDATA[31]
  PIN M_AXI_RDATA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END M_AXI_RDATA[3]
  PIN M_AXI_RDATA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END M_AXI_RDATA[4]
  PIN M_AXI_RDATA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END M_AXI_RDATA[5]
  PIN M_AXI_RDATA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END M_AXI_RDATA[6]
  PIN M_AXI_RDATA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 251.640 500.000 252.240 ;
    END
  END M_AXI_RDATA[7]
  PIN M_AXI_RDATA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 496.000 228.990 500.000 ;
    END
  END M_AXI_RDATA[8]
  PIN M_AXI_RDATA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 159.840 500.000 160.440 ;
    END
  END M_AXI_RDATA[9]
  PIN M_AXI_RREADY
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END M_AXI_RREADY
  PIN M_AXI_RRESP[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END M_AXI_RRESP[0]
  PIN M_AXI_RRESP[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END M_AXI_RRESP[1]
  PIN M_AXI_RVALID
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 438.010 496.000 438.290 500.000 ;
    END
  END M_AXI_RVALID
  PIN M_AXI_WDATA[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END M_AXI_WDATA[0]
  PIN M_AXI_WDATA[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 119.040 500.000 119.640 ;
    END
  END M_AXI_WDATA[10]
  PIN M_AXI_WDATA[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END M_AXI_WDATA[11]
  PIN M_AXI_WDATA[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 3.440 500.000 4.040 ;
    END
  END M_AXI_WDATA[12]
  PIN M_AXI_WDATA[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 496.000 119.510 500.000 ;
    END
  END M_AXI_WDATA[13]
  PIN M_AXI_WDATA[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END M_AXI_WDATA[14]
  PIN M_AXI_WDATA[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END M_AXI_WDATA[15]
  PIN M_AXI_WDATA[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END M_AXI_WDATA[16]
  PIN M_AXI_WDATA[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 68.040 500.000 68.640 ;
    END
  END M_AXI_WDATA[17]
  PIN M_AXI_WDATA[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 408.040 500.000 408.640 ;
    END
  END M_AXI_WDATA[18]
  PIN M_AXI_WDATA[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 275.440 500.000 276.040 ;
    END
  END M_AXI_WDATA[19]
  PIN M_AXI_WDATA[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END M_AXI_WDATA[1]
  PIN M_AXI_WDATA[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END M_AXI_WDATA[20]
  PIN M_AXI_WDATA[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 146.240 500.000 146.840 ;
    END
  END M_AXI_WDATA[21]
  PIN M_AXI_WDATA[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END M_AXI_WDATA[22]
  PIN M_AXI_WDATA[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 316.240 500.000 316.840 ;
    END
  END M_AXI_WDATA[23]
  PIN M_AXI_WDATA[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 459.040 500.000 459.640 ;
    END
  END M_AXI_WDATA[24]
  PIN M_AXI_WDATA[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END M_AXI_WDATA[25]
  PIN M_AXI_WDATA[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 486.240 500.000 486.840 ;
    END
  END M_AXI_WDATA[26]
  PIN M_AXI_WDATA[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END M_AXI_WDATA[27]
  PIN M_AXI_WDATA[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END M_AXI_WDATA[28]
  PIN M_AXI_WDATA[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END M_AXI_WDATA[29]
  PIN M_AXI_WDATA[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END M_AXI_WDATA[2]
  PIN M_AXI_WDATA[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END M_AXI_WDATA[30]
  PIN M_AXI_WDATA[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END M_AXI_WDATA[31]
  PIN M_AXI_WDATA[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 496.000 106.630 500.000 ;
    END
  END M_AXI_WDATA[3]
  PIN M_AXI_WDATA[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 496.000 277.290 500.000 ;
    END
  END M_AXI_WDATA[4]
  PIN M_AXI_WDATA[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END M_AXI_WDATA[5]
  PIN M_AXI_WDATA[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END M_AXI_WDATA[6]
  PIN M_AXI_WDATA[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END M_AXI_WDATA[7]
  PIN M_AXI_WDATA[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END M_AXI_WDATA[8]
  PIN M_AXI_WDATA[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 496.000 254.750 500.000 ;
    END
  END M_AXI_WDATA[9]
  PIN M_AXI_WREADY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END M_AXI_WREADY
  PIN M_AXI_WSTRB[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 496.000 425.410 500.000 ;
    END
  END M_AXI_WSTRB[0]
  PIN M_AXI_WSTRB[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 81.640 500.000 82.240 ;
    END
  END M_AXI_WSTRB[1]
  PIN M_AXI_WSTRB[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END M_AXI_WSTRB[2]
  PIN M_AXI_WSTRB[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END M_AXI_WSTRB[3]
  PIN M_AXI_WVALID
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END M_AXI_WVALID
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 487.120 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 494.280 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 494.280 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 494.280 337.990 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 494.280 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 494.280 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 494.280 334.690 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END clk
  PIN led[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END led[0]
  PIN led[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 329.840 500.000 330.440 ;
    END
  END led[1]
  PIN led[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END led[2]
  PIN led[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END led[3]
  PIN led[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 496.000 364.230 500.000 ;
    END
  END led[4]
  PIN led[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 496.000 6.810 500.000 ;
    END
  END led[5]
  PIN led[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 496.000 93.750 500.000 ;
    END
  END led[6]
  PIN led[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END led[7]
  PIN led[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END led[8]
  PIN led[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END led[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 238.040 500.000 238.640 ;
    END
  END rst_n
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 0.070 10.640 499.490 487.120 ;
      LAYER met2 ;
        RECT 0.100 495.720 6.250 496.810 ;
        RECT 7.090 495.720 19.130 496.810 ;
        RECT 19.970 495.720 32.010 496.810 ;
        RECT 32.850 495.720 44.890 496.810 ;
        RECT 45.730 495.720 54.550 496.810 ;
        RECT 55.390 495.720 67.430 496.810 ;
        RECT 68.270 495.720 80.310 496.810 ;
        RECT 81.150 495.720 93.190 496.810 ;
        RECT 94.030 495.720 106.070 496.810 ;
        RECT 106.910 495.720 118.950 496.810 ;
        RECT 119.790 495.720 128.610 496.810 ;
        RECT 129.450 495.720 141.490 496.810 ;
        RECT 142.330 495.720 154.370 496.810 ;
        RECT 155.210 495.720 167.250 496.810 ;
        RECT 168.090 495.720 180.130 496.810 ;
        RECT 180.970 495.720 193.010 496.810 ;
        RECT 193.850 495.720 202.670 496.810 ;
        RECT 203.510 495.720 215.550 496.810 ;
        RECT 216.390 495.720 228.430 496.810 ;
        RECT 229.270 495.720 241.310 496.810 ;
        RECT 242.150 495.720 254.190 496.810 ;
        RECT 255.030 495.720 267.070 496.810 ;
        RECT 267.910 495.720 276.730 496.810 ;
        RECT 277.570 495.720 289.610 496.810 ;
        RECT 290.450 495.720 302.490 496.810 ;
        RECT 303.330 495.720 315.370 496.810 ;
        RECT 316.210 495.720 328.250 496.810 ;
        RECT 329.090 495.720 341.130 496.810 ;
        RECT 341.970 495.720 350.790 496.810 ;
        RECT 351.630 495.720 363.670 496.810 ;
        RECT 364.510 495.720 376.550 496.810 ;
        RECT 377.390 495.720 389.430 496.810 ;
        RECT 390.270 495.720 402.310 496.810 ;
        RECT 403.150 495.720 415.190 496.810 ;
        RECT 416.030 495.720 424.850 496.810 ;
        RECT 425.690 495.720 437.730 496.810 ;
        RECT 438.570 495.720 450.610 496.810 ;
        RECT 451.450 495.720 463.490 496.810 ;
        RECT 464.330 495.720 476.370 496.810 ;
        RECT 477.210 495.720 489.250 496.810 ;
        RECT 490.090 495.720 498.910 496.810 ;
        RECT 0.100 4.280 499.460 495.720 ;
        RECT 0.650 3.555 9.470 4.280 ;
        RECT 10.310 3.555 22.350 4.280 ;
        RECT 23.190 3.555 35.230 4.280 ;
        RECT 36.070 3.555 48.110 4.280 ;
        RECT 48.950 3.555 60.990 4.280 ;
        RECT 61.830 3.555 73.870 4.280 ;
        RECT 74.710 3.555 83.530 4.280 ;
        RECT 84.370 3.555 96.410 4.280 ;
        RECT 97.250 3.555 109.290 4.280 ;
        RECT 110.130 3.555 122.170 4.280 ;
        RECT 123.010 3.555 135.050 4.280 ;
        RECT 135.890 3.555 147.930 4.280 ;
        RECT 148.770 3.555 157.590 4.280 ;
        RECT 158.430 3.555 170.470 4.280 ;
        RECT 171.310 3.555 183.350 4.280 ;
        RECT 184.190 3.555 196.230 4.280 ;
        RECT 197.070 3.555 209.110 4.280 ;
        RECT 209.950 3.555 221.990 4.280 ;
        RECT 222.830 3.555 231.650 4.280 ;
        RECT 232.490 3.555 244.530 4.280 ;
        RECT 245.370 3.555 257.410 4.280 ;
        RECT 258.250 3.555 270.290 4.280 ;
        RECT 271.130 3.555 283.170 4.280 ;
        RECT 284.010 3.555 296.050 4.280 ;
        RECT 296.890 3.555 305.710 4.280 ;
        RECT 306.550 3.555 318.590 4.280 ;
        RECT 319.430 3.555 331.470 4.280 ;
        RECT 332.310 3.555 344.350 4.280 ;
        RECT 345.190 3.555 357.230 4.280 ;
        RECT 358.070 3.555 370.110 4.280 ;
        RECT 370.950 3.555 379.770 4.280 ;
        RECT 380.610 3.555 392.650 4.280 ;
        RECT 393.490 3.555 405.530 4.280 ;
        RECT 406.370 3.555 418.410 4.280 ;
        RECT 419.250 3.555 431.290 4.280 ;
        RECT 432.130 3.555 444.170 4.280 ;
        RECT 445.010 3.555 453.830 4.280 ;
        RECT 454.670 3.555 466.710 4.280 ;
        RECT 467.550 3.555 479.590 4.280 ;
        RECT 480.430 3.555 492.470 4.280 ;
        RECT 493.310 3.555 499.460 4.280 ;
      LAYER met3 ;
        RECT 3.990 485.840 495.600 487.045 ;
        RECT 3.990 480.440 496.000 485.840 ;
        RECT 4.400 479.040 496.000 480.440 ;
        RECT 3.990 473.640 496.000 479.040 ;
        RECT 3.990 472.240 495.600 473.640 ;
        RECT 3.990 470.240 496.000 472.240 ;
        RECT 4.400 468.840 496.000 470.240 ;
        RECT 3.990 460.040 496.000 468.840 ;
        RECT 3.990 458.640 495.600 460.040 ;
        RECT 3.990 456.640 496.000 458.640 ;
        RECT 4.400 455.240 496.000 456.640 ;
        RECT 3.990 446.440 496.000 455.240 ;
        RECT 3.990 445.040 495.600 446.440 ;
        RECT 3.990 443.040 496.000 445.040 ;
        RECT 4.400 441.640 496.000 443.040 ;
        RECT 3.990 432.840 496.000 441.640 ;
        RECT 3.990 431.440 495.600 432.840 ;
        RECT 3.990 429.440 496.000 431.440 ;
        RECT 4.400 428.040 496.000 429.440 ;
        RECT 3.990 419.240 496.000 428.040 ;
        RECT 3.990 417.840 495.600 419.240 ;
        RECT 3.990 415.840 496.000 417.840 ;
        RECT 4.400 414.440 496.000 415.840 ;
        RECT 3.990 409.040 496.000 414.440 ;
        RECT 3.990 407.640 495.600 409.040 ;
        RECT 3.990 402.240 496.000 407.640 ;
        RECT 4.400 400.840 496.000 402.240 ;
        RECT 3.990 395.440 496.000 400.840 ;
        RECT 3.990 394.040 495.600 395.440 ;
        RECT 3.990 392.040 496.000 394.040 ;
        RECT 4.400 390.640 496.000 392.040 ;
        RECT 3.990 381.840 496.000 390.640 ;
        RECT 3.990 380.440 495.600 381.840 ;
        RECT 3.990 378.440 496.000 380.440 ;
        RECT 4.400 377.040 496.000 378.440 ;
        RECT 3.990 368.240 496.000 377.040 ;
        RECT 3.990 366.840 495.600 368.240 ;
        RECT 3.990 364.840 496.000 366.840 ;
        RECT 4.400 363.440 496.000 364.840 ;
        RECT 3.990 354.640 496.000 363.440 ;
        RECT 3.990 353.240 495.600 354.640 ;
        RECT 3.990 351.240 496.000 353.240 ;
        RECT 4.400 349.840 496.000 351.240 ;
        RECT 3.990 341.040 496.000 349.840 ;
        RECT 3.990 339.640 495.600 341.040 ;
        RECT 3.990 337.640 496.000 339.640 ;
        RECT 4.400 336.240 496.000 337.640 ;
        RECT 3.990 330.840 496.000 336.240 ;
        RECT 3.990 329.440 495.600 330.840 ;
        RECT 3.990 324.040 496.000 329.440 ;
        RECT 4.400 322.640 496.000 324.040 ;
        RECT 3.990 317.240 496.000 322.640 ;
        RECT 3.990 315.840 495.600 317.240 ;
        RECT 3.990 313.840 496.000 315.840 ;
        RECT 4.400 312.440 496.000 313.840 ;
        RECT 3.990 303.640 496.000 312.440 ;
        RECT 3.990 302.240 495.600 303.640 ;
        RECT 3.990 300.240 496.000 302.240 ;
        RECT 4.400 298.840 496.000 300.240 ;
        RECT 3.990 290.040 496.000 298.840 ;
        RECT 3.990 288.640 495.600 290.040 ;
        RECT 3.990 286.640 496.000 288.640 ;
        RECT 4.400 285.240 496.000 286.640 ;
        RECT 3.990 276.440 496.000 285.240 ;
        RECT 3.990 275.040 495.600 276.440 ;
        RECT 3.990 273.040 496.000 275.040 ;
        RECT 4.400 271.640 496.000 273.040 ;
        RECT 3.990 262.840 496.000 271.640 ;
        RECT 3.990 261.440 495.600 262.840 ;
        RECT 3.990 259.440 496.000 261.440 ;
        RECT 4.400 258.040 496.000 259.440 ;
        RECT 3.990 252.640 496.000 258.040 ;
        RECT 3.990 251.240 495.600 252.640 ;
        RECT 3.990 245.840 496.000 251.240 ;
        RECT 4.400 244.440 496.000 245.840 ;
        RECT 3.990 239.040 496.000 244.440 ;
        RECT 3.990 237.640 495.600 239.040 ;
        RECT 3.990 235.640 496.000 237.640 ;
        RECT 4.400 234.240 496.000 235.640 ;
        RECT 3.990 225.440 496.000 234.240 ;
        RECT 3.990 224.040 495.600 225.440 ;
        RECT 3.990 222.040 496.000 224.040 ;
        RECT 4.400 220.640 496.000 222.040 ;
        RECT 3.990 211.840 496.000 220.640 ;
        RECT 3.990 210.440 495.600 211.840 ;
        RECT 3.990 208.440 496.000 210.440 ;
        RECT 4.400 207.040 496.000 208.440 ;
        RECT 3.990 198.240 496.000 207.040 ;
        RECT 3.990 196.840 495.600 198.240 ;
        RECT 3.990 194.840 496.000 196.840 ;
        RECT 4.400 193.440 496.000 194.840 ;
        RECT 3.990 184.640 496.000 193.440 ;
        RECT 3.990 183.240 495.600 184.640 ;
        RECT 3.990 181.240 496.000 183.240 ;
        RECT 4.400 179.840 496.000 181.240 ;
        RECT 3.990 174.440 496.000 179.840 ;
        RECT 3.990 173.040 495.600 174.440 ;
        RECT 3.990 167.640 496.000 173.040 ;
        RECT 4.400 166.240 496.000 167.640 ;
        RECT 3.990 160.840 496.000 166.240 ;
        RECT 3.990 159.440 495.600 160.840 ;
        RECT 3.990 157.440 496.000 159.440 ;
        RECT 4.400 156.040 496.000 157.440 ;
        RECT 3.990 147.240 496.000 156.040 ;
        RECT 3.990 145.840 495.600 147.240 ;
        RECT 3.990 143.840 496.000 145.840 ;
        RECT 4.400 142.440 496.000 143.840 ;
        RECT 3.990 133.640 496.000 142.440 ;
        RECT 3.990 132.240 495.600 133.640 ;
        RECT 3.990 130.240 496.000 132.240 ;
        RECT 4.400 128.840 496.000 130.240 ;
        RECT 3.990 120.040 496.000 128.840 ;
        RECT 3.990 118.640 495.600 120.040 ;
        RECT 3.990 116.640 496.000 118.640 ;
        RECT 4.400 115.240 496.000 116.640 ;
        RECT 3.990 106.440 496.000 115.240 ;
        RECT 3.990 105.040 495.600 106.440 ;
        RECT 3.990 103.040 496.000 105.040 ;
        RECT 4.400 101.640 496.000 103.040 ;
        RECT 3.990 96.240 496.000 101.640 ;
        RECT 3.990 94.840 495.600 96.240 ;
        RECT 3.990 89.440 496.000 94.840 ;
        RECT 4.400 88.040 496.000 89.440 ;
        RECT 3.990 82.640 496.000 88.040 ;
        RECT 3.990 81.240 495.600 82.640 ;
        RECT 3.990 79.240 496.000 81.240 ;
        RECT 4.400 77.840 496.000 79.240 ;
        RECT 3.990 69.040 496.000 77.840 ;
        RECT 3.990 67.640 495.600 69.040 ;
        RECT 3.990 65.640 496.000 67.640 ;
        RECT 4.400 64.240 496.000 65.640 ;
        RECT 3.990 55.440 496.000 64.240 ;
        RECT 3.990 54.040 495.600 55.440 ;
        RECT 3.990 52.040 496.000 54.040 ;
        RECT 4.400 50.640 496.000 52.040 ;
        RECT 3.990 41.840 496.000 50.640 ;
        RECT 3.990 40.440 495.600 41.840 ;
        RECT 3.990 38.440 496.000 40.440 ;
        RECT 4.400 37.040 496.000 38.440 ;
        RECT 3.990 28.240 496.000 37.040 ;
        RECT 3.990 26.840 495.600 28.240 ;
        RECT 3.990 24.840 496.000 26.840 ;
        RECT 4.400 23.440 496.000 24.840 ;
        RECT 3.990 18.040 496.000 23.440 ;
        RECT 3.990 16.640 495.600 18.040 ;
        RECT 3.990 11.240 496.000 16.640 ;
        RECT 4.400 9.840 496.000 11.240 ;
        RECT 3.990 4.440 496.000 9.840 ;
        RECT 3.990 3.575 495.600 4.440 ;
  END
END riscv_pipeline_top
END LIBRARY

