module vajra_caravel_soc (wb_clk_i,
    wb_rst_i,
    io_in,
    io_oeb,
    io_out);
 input wb_clk_i;
 input wb_rst_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire \u_cpu.ALUResult_E[0] ;
 wire \u_cpu.ALUResult_E[10] ;
 wire \u_cpu.ALUResult_E[11] ;
 wire \u_cpu.ALUResult_E[12] ;
 wire \u_cpu.ALUResult_E[13] ;
 wire \u_cpu.ALUResult_E[14] ;
 wire \u_cpu.ALUResult_E[15] ;
 wire \u_cpu.ALUResult_E[16] ;
 wire \u_cpu.ALUResult_E[17] ;
 wire \u_cpu.ALUResult_E[18] ;
 wire \u_cpu.ALUResult_E[19] ;
 wire \u_cpu.ALUResult_E[1] ;
 wire \u_cpu.ALUResult_E[20] ;
 wire \u_cpu.ALUResult_E[21] ;
 wire \u_cpu.ALUResult_E[22] ;
 wire \u_cpu.ALUResult_E[23] ;
 wire \u_cpu.ALUResult_E[24] ;
 wire \u_cpu.ALUResult_E[25] ;
 wire \u_cpu.ALUResult_E[26] ;
 wire \u_cpu.ALUResult_E[27] ;
 wire \u_cpu.ALUResult_E[28] ;
 wire \u_cpu.ALUResult_E[29] ;
 wire \u_cpu.ALUResult_E[2] ;
 wire \u_cpu.ALUResult_E[30] ;
 wire \u_cpu.ALUResult_E[31] ;
 wire \u_cpu.ALUResult_E[3] ;
 wire \u_cpu.ALUResult_E[4] ;
 wire \u_cpu.ALUResult_E[5] ;
 wire \u_cpu.ALUResult_E[6] ;
 wire \u_cpu.ALUResult_E[7] ;
 wire \u_cpu.ALUResult_E[8] ;
 wire \u_cpu.ALUResult_E[9] ;
 wire \u_cpu.Instr_D[0] ;
 wire \u_cpu.Instr_D[10] ;
 wire \u_cpu.Instr_D[11] ;
 wire \u_cpu.Instr_D[12] ;
 wire \u_cpu.Instr_D[13] ;
 wire \u_cpu.Instr_D[14] ;
 wire \u_cpu.Instr_D[15] ;
 wire \u_cpu.Instr_D[16] ;
 wire \u_cpu.Instr_D[17] ;
 wire \u_cpu.Instr_D[18] ;
 wire \u_cpu.Instr_D[19] ;
 wire \u_cpu.Instr_D[1] ;
 wire \u_cpu.Instr_D[20] ;
 wire \u_cpu.Instr_D[21] ;
 wire \u_cpu.Instr_D[22] ;
 wire \u_cpu.Instr_D[23] ;
 wire \u_cpu.Instr_D[24] ;
 wire \u_cpu.Instr_D[25] ;
 wire \u_cpu.Instr_D[26] ;
 wire \u_cpu.Instr_D[27] ;
 wire \u_cpu.Instr_D[28] ;
 wire \u_cpu.Instr_D[29] ;
 wire \u_cpu.Instr_D[2] ;
 wire \u_cpu.Instr_D[30] ;
 wire \u_cpu.Instr_D[31] ;
 wire \u_cpu.Instr_D[3] ;
 wire \u_cpu.Instr_D[4] ;
 wire \u_cpu.Instr_D[5] ;
 wire \u_cpu.Instr_D[6] ;
 wire \u_cpu.Instr_D[7] ;
 wire \u_cpu.Instr_D[8] ;
 wire \u_cpu.Instr_D[9] ;
 wire \u_cpu.Instr_F[0] ;
 wire \u_cpu.Instr_F[10] ;
 wire \u_cpu.Instr_F[11] ;
 wire \u_cpu.Instr_F[12] ;
 wire \u_cpu.Instr_F[13] ;
 wire \u_cpu.Instr_F[14] ;
 wire \u_cpu.Instr_F[15] ;
 wire \u_cpu.Instr_F[16] ;
 wire \u_cpu.Instr_F[17] ;
 wire \u_cpu.Instr_F[18] ;
 wire \u_cpu.Instr_F[19] ;
 wire \u_cpu.Instr_F[1] ;
 wire \u_cpu.Instr_F[20] ;
 wire \u_cpu.Instr_F[21] ;
 wire \u_cpu.Instr_F[22] ;
 wire \u_cpu.Instr_F[23] ;
 wire \u_cpu.Instr_F[24] ;
 wire \u_cpu.Instr_F[25] ;
 wire \u_cpu.Instr_F[26] ;
 wire \u_cpu.Instr_F[27] ;
 wire \u_cpu.Instr_F[28] ;
 wire \u_cpu.Instr_F[29] ;
 wire \u_cpu.Instr_F[2] ;
 wire \u_cpu.Instr_F[30] ;
 wire \u_cpu.Instr_F[31] ;
 wire \u_cpu.Instr_F[3] ;
 wire \u_cpu.Instr_F[4] ;
 wire \u_cpu.Instr_F[5] ;
 wire \u_cpu.Instr_F[6] ;
 wire \u_cpu.Instr_F[7] ;
 wire \u_cpu.Instr_F[8] ;
 wire \u_cpu.Instr_F[9] ;
 wire \u_cpu.PC_F[0] ;
 wire \u_cpu.PC_F[10] ;
 wire \u_cpu.PC_F[11] ;
 wire \u_cpu.PC_F[12] ;
 wire \u_cpu.PC_F[13] ;
 wire \u_cpu.PC_F[14] ;
 wire \u_cpu.PC_F[15] ;
 wire \u_cpu.PC_F[16] ;
 wire \u_cpu.PC_F[17] ;
 wire \u_cpu.PC_F[18] ;
 wire \u_cpu.PC_F[19] ;
 wire \u_cpu.PC_F[1] ;
 wire \u_cpu.PC_F[20] ;
 wire \u_cpu.PC_F[21] ;
 wire \u_cpu.PC_F[22] ;
 wire \u_cpu.PC_F[23] ;
 wire \u_cpu.PC_F[24] ;
 wire \u_cpu.PC_F[25] ;
 wire \u_cpu.PC_F[26] ;
 wire \u_cpu.PC_F[27] ;
 wire \u_cpu.PC_F[28] ;
 wire \u_cpu.PC_F[29] ;
 wire \u_cpu.PC_F[2] ;
 wire \u_cpu.PC_F[30] ;
 wire \u_cpu.PC_F[31] ;
 wire \u_cpu.PC_F[3] ;
 wire \u_cpu.PC_F[4] ;
 wire \u_cpu.PC_F[5] ;
 wire \u_cpu.PC_F[6] ;
 wire \u_cpu.PC_F[7] ;
 wire \u_cpu.PC_F[8] ;
 wire \u_cpu.PC_F[9] ;
 wire \u_cpu.counter[0] ;
 wire \u_cpu.counter[10] ;
 wire \u_cpu.counter[11] ;
 wire \u_cpu.counter[12] ;
 wire \u_cpu.counter[13] ;
 wire \u_cpu.counter[14] ;
 wire \u_cpu.counter[15] ;
 wire \u_cpu.counter[16] ;
 wire \u_cpu.counter[17] ;
 wire \u_cpu.counter[18] ;
 wire \u_cpu.counter[19] ;
 wire \u_cpu.counter[1] ;
 wire \u_cpu.counter[20] ;
 wire \u_cpu.counter[21] ;
 wire \u_cpu.counter[22] ;
 wire \u_cpu.counter[23] ;
 wire \u_cpu.counter[24] ;
 wire \u_cpu.counter[25] ;
 wire \u_cpu.counter[2] ;
 wire \u_cpu.counter[3] ;
 wire \u_cpu.counter[4] ;
 wire \u_cpu.counter[5] ;
 wire \u_cpu.counter[6] ;
 wire \u_cpu.counter[7] ;
 wire \u_cpu.counter[8] ;
 wire \u_cpu.counter[9] ;

 sky130_fd_sc_hd__and3_2 _219_ (.A(\u_cpu.ALUResult_E[28] ),
    .B(\u_cpu.ALUResult_E[27] ),
    .C(\u_cpu.ALUResult_E[26] ),
    .X(_112_));
 sky130_fd_sc_hd__and2_2 _220_ (.A(\u_cpu.ALUResult_E[29] ),
    .B(_112_),
    .X(_113_));
 sky130_fd_sc_hd__and3_2 _221_ (.A(\u_cpu.ALUResult_E[24] ),
    .B(\u_cpu.ALUResult_E[23] ),
    .C(\u_cpu.ALUResult_E[22] ),
    .X(_114_));
 sky130_fd_sc_hd__and2_2 _222_ (.A(\u_cpu.ALUResult_E[25] ),
    .B(_114_),
    .X(_115_));
 sky130_fd_sc_hd__and4_2 _223_ (.A(\u_cpu.counter[0] ),
    .B(\u_cpu.counter[1] ),
    .C(\u_cpu.counter[3] ),
    .D(\u_cpu.counter[2] ),
    .X(_116_));
 sky130_fd_sc_hd__buf_1 _224_ (.A(_116_),
    .X(_117_));
 sky130_fd_sc_hd__and4_2 _225_ (.A(\u_cpu.counter[5] ),
    .B(\u_cpu.counter[4] ),
    .C(\u_cpu.counter[7] ),
    .D(\u_cpu.counter[6] ),
    .X(_118_));
 sky130_fd_sc_hd__and4_2 _226_ (.A(\u_cpu.counter[9] ),
    .B(\u_cpu.counter[8] ),
    .C(\u_cpu.counter[10] ),
    .D(\u_cpu.counter[11] ),
    .X(_119_));
 sky130_fd_sc_hd__and4_2 _227_ (.A(\u_cpu.counter[13] ),
    .B(\u_cpu.counter[12] ),
    .C(\u_cpu.counter[15] ),
    .D(\u_cpu.counter[14] ),
    .X(_120_));
 sky130_fd_sc_hd__and4_2 _228_ (.A(_117_),
    .B(_118_),
    .C(_119_),
    .D(_120_),
    .X(_121_));
 sky130_fd_sc_hd__buf_1 _229_ (.A(_121_),
    .X(_122_));
 sky130_fd_sc_hd__and4_2 _230_ (.A(\u_cpu.counter[17] ),
    .B(\u_cpu.counter[16] ),
    .C(\u_cpu.counter[19] ),
    .D(\u_cpu.counter[18] ),
    .X(_123_));
 sky130_fd_sc_hd__and4_2 _231_ (.A(\u_cpu.counter[21] ),
    .B(\u_cpu.counter[20] ),
    .C(\u_cpu.counter[23] ),
    .D(\u_cpu.counter[22] ),
    .X(_124_));
 sky130_fd_sc_hd__and2_2 _232_ (.A(\u_cpu.counter[24] ),
    .B(\u_cpu.counter[25] ),
    .X(_125_));
 sky130_fd_sc_hd__and4_2 _233_ (.A(_122_),
    .B(_123_),
    .C(_124_),
    .D(_125_),
    .X(_126_));
 sky130_fd_sc_hd__buf_1 _234_ (.A(_126_),
    .X(_127_));
 sky130_fd_sc_hd__and2_2 _235_ (.A(\u_cpu.ALUResult_E[19] ),
    .B(\u_cpu.ALUResult_E[18] ),
    .X(_128_));
 sky130_fd_sc_hd__and4_2 _236_ (.A(io_out[35]),
    .B(io_out[34]),
    .C(io_out[33]),
    .D(io_out[32]),
    .X(_129_));
 sky130_fd_sc_hd__and2_2 _237_ (.A(io_out[37]),
    .B(io_out[36]),
    .X(_130_));
 sky130_fd_sc_hd__and3_2 _238_ (.A(\u_cpu.ALUResult_E[17] ),
    .B(\u_cpu.ALUResult_E[16] ),
    .C(_130_),
    .X(_131_));
 sky130_fd_sc_hd__and2_2 _239_ (.A(io_out[29]),
    .B(io_out[28]),
    .X(_132_));
 sky130_fd_sc_hd__and4_2 _240_ (.A(io_out[27]),
    .B(io_out[26]),
    .C(io_out[25]),
    .D(io_out[24]),
    .X(_133_));
 sky130_fd_sc_hd__and4_2 _241_ (.A(io_out[31]),
    .B(io_out[30]),
    .C(_132_),
    .D(_133_),
    .X(_134_));
 sky130_fd_sc_hd__and4_2 _242_ (.A(_128_),
    .B(_129_),
    .C(_131_),
    .D(_134_),
    .X(_135_));
 sky130_fd_sc_hd__and4_2 _243_ (.A(\u_cpu.ALUResult_E[21] ),
    .B(\u_cpu.ALUResult_E[20] ),
    .C(_127_),
    .D(_135_),
    .X(_136_));
 sky130_fd_sc_hd__buf_1 _244_ (.A(_136_),
    .X(_137_));
 sky130_fd_sc_hd__and4_2 _245_ (.A(\u_cpu.ALUResult_E[30] ),
    .B(_113_),
    .C(_115_),
    .D(_137_),
    .X(_138_));
 sky130_fd_sc_hd__xor2_2 _246_ (.A(\u_cpu.ALUResult_E[31] ),
    .B(_138_),
    .X(_111_));
 sky130_fd_sc_hd__and3_2 _247_ (.A(_113_),
    .B(_115_),
    .C(_136_),
    .X(_139_));
 sky130_fd_sc_hd__xor2_2 _248_ (.A(\u_cpu.ALUResult_E[30] ),
    .B(_139_),
    .X(_110_));
 sky130_fd_sc_hd__a31o_2 _249_ (.A1(_112_),
    .A2(_115_),
    .A3(_136_),
    .B1(\u_cpu.ALUResult_E[29] ),
    .X(_140_));
 sky130_fd_sc_hd__and2b_2 _250_ (.A_N(_139_),
    .B(_140_),
    .X(_141_));
 sky130_fd_sc_hd__buf_1 _251_ (.A(_141_),
    .X(_109_));
 sky130_fd_sc_hd__inv_2 _252_ (.A(_112_),
    .Y(_142_));
 sky130_fd_sc_hd__nand2_2 _253_ (.A(_115_),
    .B(_137_),
    .Y(_143_));
 sky130_fd_sc_hd__a41o_2 _254_ (.A1(\u_cpu.ALUResult_E[27] ),
    .A2(\u_cpu.ALUResult_E[26] ),
    .A3(_115_),
    .A4(_137_),
    .B1(\u_cpu.ALUResult_E[28] ),
    .X(_144_));
 sky130_fd_sc_hd__o21a_2 _255_ (.A1(_142_),
    .A2(_143_),
    .B1(_144_),
    .X(_108_));
 sky130_fd_sc_hd__nand2_2 _256_ (.A(\u_cpu.ALUResult_E[27] ),
    .B(\u_cpu.ALUResult_E[26] ),
    .Y(_145_));
 sky130_fd_sc_hd__a31o_2 _257_ (.A1(\u_cpu.ALUResult_E[26] ),
    .A2(_115_),
    .A3(_137_),
    .B1(\u_cpu.ALUResult_E[27] ),
    .X(_146_));
 sky130_fd_sc_hd__o21a_2 _258_ (.A1(_145_),
    .A2(_143_),
    .B1(_146_),
    .X(_107_));
 sky130_fd_sc_hd__xnor2_2 _259_ (.A(\u_cpu.ALUResult_E[26] ),
    .B(_143_),
    .Y(_106_));
 sky130_fd_sc_hd__a21o_2 _260_ (.A1(_114_),
    .A2(_137_),
    .B1(\u_cpu.ALUResult_E[25] ),
    .X(_147_));
 sky130_fd_sc_hd__and2_2 _261_ (.A(_143_),
    .B(_147_),
    .X(_148_));
 sky130_fd_sc_hd__buf_1 _262_ (.A(_148_),
    .X(_105_));
 sky130_fd_sc_hd__and3_2 _263_ (.A(\u_cpu.ALUResult_E[23] ),
    .B(\u_cpu.ALUResult_E[22] ),
    .C(_137_),
    .X(_149_));
 sky130_fd_sc_hd__o2bb2a_2 _264_ (.A1_N(_114_),
    .A2_N(_137_),
    .B1(_149_),
    .B2(\u_cpu.ALUResult_E[24] ),
    .X(_104_));
 sky130_fd_sc_hd__a21oi_2 _265_ (.A1(\u_cpu.ALUResult_E[22] ),
    .A2(_137_),
    .B1(\u_cpu.ALUResult_E[23] ),
    .Y(_150_));
 sky130_fd_sc_hd__nor2_2 _266_ (.A(_149_),
    .B(_150_),
    .Y(_103_));
 sky130_fd_sc_hd__xor2_2 _267_ (.A(\u_cpu.ALUResult_E[22] ),
    .B(_137_),
    .X(_102_));
 sky130_fd_sc_hd__buf_1 _268_ (.A(_127_),
    .X(_151_));
 sky130_fd_sc_hd__and2_2 _269_ (.A(_151_),
    .B(_135_),
    .X(_152_));
 sky130_fd_sc_hd__a21oi_2 _270_ (.A1(\u_cpu.ALUResult_E[20] ),
    .A2(_152_),
    .B1(\u_cpu.ALUResult_E[21] ),
    .Y(_153_));
 sky130_fd_sc_hd__nor2_2 _271_ (.A(_137_),
    .B(_153_),
    .Y(_101_));
 sky130_fd_sc_hd__xor2_2 _272_ (.A(\u_cpu.ALUResult_E[20] ),
    .B(_152_),
    .X(_100_));
 sky130_fd_sc_hd__and3_2 _273_ (.A(_129_),
    .B(_131_),
    .C(_134_),
    .X(_154_));
 sky130_fd_sc_hd__a31o_2 _274_ (.A1(\u_cpu.ALUResult_E[18] ),
    .A2(_127_),
    .A3(_154_),
    .B1(\u_cpu.ALUResult_E[19] ),
    .X(_155_));
 sky130_fd_sc_hd__and2b_2 _275_ (.A_N(_152_),
    .B(_155_),
    .X(_156_));
 sky130_fd_sc_hd__buf_1 _276_ (.A(_156_),
    .X(_099_));
 sky130_fd_sc_hd__nand2_2 _277_ (.A(_151_),
    .B(_154_),
    .Y(_157_));
 sky130_fd_sc_hd__xnor2_2 _278_ (.A(\u_cpu.ALUResult_E[18] ),
    .B(_157_),
    .Y(_098_));
 sky130_fd_sc_hd__inv_2 _279_ (.A(\u_cpu.ALUResult_E[16] ),
    .Y(_158_));
 sky130_fd_sc_hd__nand4_2 _280_ (.A(_127_),
    .B(_129_),
    .C(_130_),
    .D(_134_),
    .Y(_159_));
 sky130_fd_sc_hd__nor2_2 _281_ (.A(_158_),
    .B(_159_),
    .Y(_160_));
 sky130_fd_sc_hd__o21a_2 _282_ (.A1(\u_cpu.ALUResult_E[17] ),
    .A2(_160_),
    .B1(_157_),
    .X(_097_));
 sky130_fd_sc_hd__nand2_2 _283_ (.A(_158_),
    .B(_159_),
    .Y(_161_));
 sky130_fd_sc_hd__and2b_2 _284_ (.A_N(_160_),
    .B(_161_),
    .X(_162_));
 sky130_fd_sc_hd__buf_1 _285_ (.A(_162_),
    .X(_096_));
 sky130_fd_sc_hd__and3_2 _286_ (.A(_127_),
    .B(_129_),
    .C(_134_),
    .X(_163_));
 sky130_fd_sc_hd__a21o_2 _287_ (.A1(io_out[36]),
    .A2(_163_),
    .B1(io_out[37]),
    .X(_164_));
 sky130_fd_sc_hd__and2_2 _288_ (.A(_159_),
    .B(_164_),
    .X(_165_));
 sky130_fd_sc_hd__buf_1 _289_ (.A(_165_),
    .X(_095_));
 sky130_fd_sc_hd__xor2_2 _290_ (.A(io_out[36]),
    .B(_163_),
    .X(_094_));
 sky130_fd_sc_hd__and4_2 _291_ (.A(io_out[33]),
    .B(io_out[32]),
    .C(_127_),
    .D(_134_),
    .X(_166_));
 sky130_fd_sc_hd__a21oi_2 _292_ (.A1(io_out[34]),
    .A2(_166_),
    .B1(io_out[35]),
    .Y(_167_));
 sky130_fd_sc_hd__nor2_2 _293_ (.A(_163_),
    .B(_167_),
    .Y(_093_));
 sky130_fd_sc_hd__xor2_2 _294_ (.A(io_out[34]),
    .B(_166_),
    .X(_092_));
 sky130_fd_sc_hd__a31o_2 _295_ (.A1(io_out[32]),
    .A2(_127_),
    .A3(_134_),
    .B1(io_out[33]),
    .X(_168_));
 sky130_fd_sc_hd__and2b_2 _296_ (.A_N(_166_),
    .B(_168_),
    .X(_169_));
 sky130_fd_sc_hd__buf_1 _297_ (.A(_169_),
    .X(_091_));
 sky130_fd_sc_hd__nand2_2 _298_ (.A(_151_),
    .B(_134_),
    .Y(_170_));
 sky130_fd_sc_hd__xnor2_2 _299_ (.A(io_out[32]),
    .B(_170_),
    .Y(_090_));
 sky130_fd_sc_hd__and2_2 _300_ (.A(_132_),
    .B(_133_),
    .X(_171_));
 sky130_fd_sc_hd__a31o_2 _301_ (.A1(io_out[30]),
    .A2(_127_),
    .A3(_171_),
    .B1(io_out[31]),
    .X(_172_));
 sky130_fd_sc_hd__and2_2 _302_ (.A(_170_),
    .B(_172_),
    .X(_173_));
 sky130_fd_sc_hd__buf_1 _303_ (.A(_173_),
    .X(_089_));
 sky130_fd_sc_hd__nand2_2 _304_ (.A(_151_),
    .B(_171_),
    .Y(_174_));
 sky130_fd_sc_hd__xnor2_2 _305_ (.A(io_out[30]),
    .B(_174_),
    .Y(_088_));
 sky130_fd_sc_hd__and3_2 _306_ (.A(io_out[28]),
    .B(_151_),
    .C(_133_),
    .X(_175_));
 sky130_fd_sc_hd__o21a_2 _307_ (.A1(io_out[29]),
    .A2(_175_),
    .B1(_174_),
    .X(_087_));
 sky130_fd_sc_hd__a21oi_2 _308_ (.A1(_151_),
    .A2(_133_),
    .B1(io_out[28]),
    .Y(_176_));
 sky130_fd_sc_hd__nor2_2 _309_ (.A(_175_),
    .B(_176_),
    .Y(_086_));
 sky130_fd_sc_hd__and3_2 _310_ (.A(io_out[25]),
    .B(io_out[24]),
    .C(_127_),
    .X(_177_));
 sky130_fd_sc_hd__and2_2 _311_ (.A(io_out[26]),
    .B(_177_),
    .X(_178_));
 sky130_fd_sc_hd__o2bb2a_2 _312_ (.A1_N(_151_),
    .A2_N(_133_),
    .B1(_178_),
    .B2(io_out[27]),
    .X(_085_));
 sky130_fd_sc_hd__xor2_2 _313_ (.A(io_out[26]),
    .B(_177_),
    .X(_084_));
 sky130_fd_sc_hd__a21oi_2 _314_ (.A1(io_out[24]),
    .A2(_151_),
    .B1(io_out[25]),
    .Y(_179_));
 sky130_fd_sc_hd__nor2_2 _315_ (.A(_177_),
    .B(_179_),
    .Y(_083_));
 sky130_fd_sc_hd__xor2_2 _316_ (.A(io_out[24]),
    .B(_151_),
    .X(_082_));
 sky130_fd_sc_hd__inv_2 _317_ (.A(\u_cpu.counter[0] ),
    .Y(_000_));
 sky130_fd_sc_hd__nand2_2 _318_ (.A(\u_cpu.counter[0] ),
    .B(\u_cpu.counter[1] ),
    .Y(_180_));
 sky130_fd_sc_hd__or2_2 _319_ (.A(\u_cpu.counter[0] ),
    .B(\u_cpu.counter[1] ),
    .X(_181_));
 sky130_fd_sc_hd__and2_2 _320_ (.A(_180_),
    .B(_181_),
    .X(_182_));
 sky130_fd_sc_hd__buf_1 _321_ (.A(_182_),
    .X(_011_));
 sky130_fd_sc_hd__xnor2_2 _322_ (.A(\u_cpu.counter[2] ),
    .B(_180_),
    .Y(_018_));
 sky130_fd_sc_hd__a31o_2 _323_ (.A1(\u_cpu.counter[0] ),
    .A2(\u_cpu.counter[1] ),
    .A3(\u_cpu.counter[2] ),
    .B1(\u_cpu.counter[3] ),
    .X(_183_));
 sky130_fd_sc_hd__and2b_2 _324_ (.A_N(_117_),
    .B(_183_),
    .X(_184_));
 sky130_fd_sc_hd__buf_1 _325_ (.A(_184_),
    .X(_019_));
 sky130_fd_sc_hd__xor2_2 _326_ (.A(\u_cpu.counter[4] ),
    .B(_117_),
    .X(_020_));
 sky130_fd_sc_hd__nand2_2 _327_ (.A(\u_cpu.counter[4] ),
    .B(_117_),
    .Y(_185_));
 sky130_fd_sc_hd__xnor2_2 _328_ (.A(\u_cpu.counter[5] ),
    .B(_185_),
    .Y(_021_));
 sky130_fd_sc_hd__and4_2 _329_ (.A(\u_cpu.counter[5] ),
    .B(\u_cpu.counter[4] ),
    .C(\u_cpu.counter[6] ),
    .D(_117_),
    .X(_186_));
 sky130_fd_sc_hd__a31o_2 _330_ (.A1(\u_cpu.counter[5] ),
    .A2(\u_cpu.counter[4] ),
    .A3(_117_),
    .B1(\u_cpu.counter[6] ),
    .X(_187_));
 sky130_fd_sc_hd__and2b_2 _331_ (.A_N(_186_),
    .B(_187_),
    .X(_188_));
 sky130_fd_sc_hd__buf_1 _332_ (.A(_188_),
    .X(_022_));
 sky130_fd_sc_hd__and2_2 _333_ (.A(_117_),
    .B(_118_),
    .X(_189_));
 sky130_fd_sc_hd__o21ba_2 _334_ (.A1(\u_cpu.counter[7] ),
    .A2(_186_),
    .B1_N(_189_),
    .X(_023_));
 sky130_fd_sc_hd__xor2_2 _335_ (.A(\u_cpu.counter[8] ),
    .B(_189_),
    .X(_024_));
 sky130_fd_sc_hd__and3_2 _336_ (.A(\u_cpu.counter[9] ),
    .B(\u_cpu.counter[8] ),
    .C(_189_),
    .X(_190_));
 sky130_fd_sc_hd__a31o_2 _337_ (.A1(\u_cpu.counter[8] ),
    .A2(_117_),
    .A3(_118_),
    .B1(\u_cpu.counter[9] ),
    .X(_191_));
 sky130_fd_sc_hd__and2b_2 _338_ (.A_N(_190_),
    .B(_191_),
    .X(_192_));
 sky130_fd_sc_hd__buf_1 _339_ (.A(_192_),
    .X(_025_));
 sky130_fd_sc_hd__xor2_2 _340_ (.A(\u_cpu.counter[10] ),
    .B(_190_),
    .X(_001_));
 sky130_fd_sc_hd__and3_2 _341_ (.A(_117_),
    .B(_118_),
    .C(_119_),
    .X(_193_));
 sky130_fd_sc_hd__a21o_2 _342_ (.A1(\u_cpu.counter[10] ),
    .A2(_190_),
    .B1(\u_cpu.counter[11] ),
    .X(_194_));
 sky130_fd_sc_hd__and2b_2 _343_ (.A_N(_193_),
    .B(_194_),
    .X(_195_));
 sky130_fd_sc_hd__buf_1 _344_ (.A(_195_),
    .X(_002_));
 sky130_fd_sc_hd__and2_2 _345_ (.A(\u_cpu.counter[12] ),
    .B(_193_),
    .X(_196_));
 sky130_fd_sc_hd__nor2_2 _346_ (.A(\u_cpu.counter[12] ),
    .B(_193_),
    .Y(_197_));
 sky130_fd_sc_hd__nor2_2 _347_ (.A(_196_),
    .B(_197_),
    .Y(_003_));
 sky130_fd_sc_hd__xor2_2 _348_ (.A(\u_cpu.counter[13] ),
    .B(_196_),
    .X(_004_));
 sky130_fd_sc_hd__a21oi_2 _349_ (.A1(\u_cpu.counter[13] ),
    .A2(_196_),
    .B1(\u_cpu.counter[14] ),
    .Y(_198_));
 sky130_fd_sc_hd__and3_2 _350_ (.A(\u_cpu.counter[13] ),
    .B(\u_cpu.counter[14] ),
    .C(_196_),
    .X(_199_));
 sky130_fd_sc_hd__nor2_2 _351_ (.A(_198_),
    .B(_199_),
    .Y(_005_));
 sky130_fd_sc_hd__o21ba_2 _352_ (.A1(\u_cpu.counter[15] ),
    .A2(_199_),
    .B1_N(_122_),
    .X(_006_));
 sky130_fd_sc_hd__xor2_2 _353_ (.A(\u_cpu.counter[16] ),
    .B(_122_),
    .X(_007_));
 sky130_fd_sc_hd__and3_2 _354_ (.A(\u_cpu.counter[17] ),
    .B(\u_cpu.counter[16] ),
    .C(_122_),
    .X(_200_));
 sky130_fd_sc_hd__a21oi_2 _355_ (.A1(\u_cpu.counter[16] ),
    .A2(_122_),
    .B1(\u_cpu.counter[17] ),
    .Y(_201_));
 sky130_fd_sc_hd__nor2_2 _356_ (.A(_200_),
    .B(_201_),
    .Y(_008_));
 sky130_fd_sc_hd__and2_2 _357_ (.A(\u_cpu.counter[18] ),
    .B(_200_),
    .X(_202_));
 sky130_fd_sc_hd__nor2_2 _358_ (.A(\u_cpu.counter[18] ),
    .B(_200_),
    .Y(_203_));
 sky130_fd_sc_hd__nor2_2 _359_ (.A(_202_),
    .B(_203_),
    .Y(_009_));
 sky130_fd_sc_hd__and2_2 _360_ (.A(_122_),
    .B(_123_),
    .X(_204_));
 sky130_fd_sc_hd__o21ba_2 _361_ (.A1(\u_cpu.counter[19] ),
    .A2(_202_),
    .B1_N(_204_),
    .X(_010_));
 sky130_fd_sc_hd__xor2_2 _362_ (.A(\u_cpu.counter[20] ),
    .B(_204_),
    .X(_012_));
 sky130_fd_sc_hd__and3_2 _363_ (.A(\u_cpu.counter[21] ),
    .B(\u_cpu.counter[20] ),
    .C(_204_),
    .X(_205_));
 sky130_fd_sc_hd__a31o_2 _364_ (.A1(\u_cpu.counter[20] ),
    .A2(_122_),
    .A3(_123_),
    .B1(\u_cpu.counter[21] ),
    .X(_206_));
 sky130_fd_sc_hd__and2b_2 _365_ (.A_N(_205_),
    .B(_206_),
    .X(_207_));
 sky130_fd_sc_hd__buf_1 _366_ (.A(_207_),
    .X(_013_));
 sky130_fd_sc_hd__and2_2 _367_ (.A(\u_cpu.counter[22] ),
    .B(_205_),
    .X(_208_));
 sky130_fd_sc_hd__nor2_2 _368_ (.A(\u_cpu.counter[22] ),
    .B(_205_),
    .Y(_209_));
 sky130_fd_sc_hd__nor2_2 _369_ (.A(_208_),
    .B(_209_),
    .Y(_014_));
 sky130_fd_sc_hd__and3_2 _370_ (.A(_122_),
    .B(_123_),
    .C(_124_),
    .X(_210_));
 sky130_fd_sc_hd__o21ba_2 _371_ (.A1(\u_cpu.counter[23] ),
    .A2(_208_),
    .B1_N(_210_),
    .X(_015_));
 sky130_fd_sc_hd__and2_2 _372_ (.A(\u_cpu.counter[24] ),
    .B(_210_),
    .X(_211_));
 sky130_fd_sc_hd__nor2_2 _373_ (.A(\u_cpu.counter[24] ),
    .B(_210_),
    .Y(_212_));
 sky130_fd_sc_hd__nor2_2 _374_ (.A(_211_),
    .B(_212_),
    .Y(_016_));
 sky130_fd_sc_hd__o21ba_2 _375_ (.A1(\u_cpu.counter[25] ),
    .A2(_211_),
    .B1_N(_151_),
    .X(_017_));
 sky130_fd_sc_hd__buf_1 _376_ (.A(wb_rst_i),
    .X(_213_));
 sky130_fd_sc_hd__buf_1 _377_ (.A(_213_),
    .X(_214_));
 sky130_fd_sc_hd__inv_2 _378_ (.A(_214_),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _379_ (.A(_214_),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _380_ (.A(_214_),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _381_ (.A(_214_),
    .Y(_029_));
 sky130_fd_sc_hd__inv_2 _382_ (.A(_214_),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _383_ (.A(_214_),
    .Y(_031_));
 sky130_fd_sc_hd__inv_2 _384_ (.A(_214_),
    .Y(_032_));
 sky130_fd_sc_hd__inv_2 _385_ (.A(_214_),
    .Y(_033_));
 sky130_fd_sc_hd__inv_2 _386_ (.A(_214_),
    .Y(_034_));
 sky130_fd_sc_hd__inv_2 _387_ (.A(_214_),
    .Y(_035_));
 sky130_fd_sc_hd__buf_1 _388_ (.A(_213_),
    .X(_215_));
 sky130_fd_sc_hd__inv_2 _389_ (.A(_215_),
    .Y(_036_));
 sky130_fd_sc_hd__inv_2 _390_ (.A(_215_),
    .Y(_037_));
 sky130_fd_sc_hd__inv_2 _391_ (.A(_215_),
    .Y(_038_));
 sky130_fd_sc_hd__inv_2 _392_ (.A(_215_),
    .Y(_039_));
 sky130_fd_sc_hd__inv_2 _393_ (.A(_215_),
    .Y(_040_));
 sky130_fd_sc_hd__inv_2 _394_ (.A(_215_),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _395_ (.A(_215_),
    .Y(_042_));
 sky130_fd_sc_hd__inv_2 _396_ (.A(_215_),
    .Y(_043_));
 sky130_fd_sc_hd__inv_2 _397_ (.A(_215_),
    .Y(_044_));
 sky130_fd_sc_hd__inv_2 _398_ (.A(_215_),
    .Y(_045_));
 sky130_fd_sc_hd__buf_1 _399_ (.A(_213_),
    .X(_216_));
 sky130_fd_sc_hd__inv_2 _400_ (.A(_216_),
    .Y(_046_));
 sky130_fd_sc_hd__inv_2 _401_ (.A(_216_),
    .Y(_047_));
 sky130_fd_sc_hd__inv_2 _402_ (.A(_216_),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _403_ (.A(_216_),
    .Y(_049_));
 sky130_fd_sc_hd__inv_2 _404_ (.A(_216_),
    .Y(_050_));
 sky130_fd_sc_hd__inv_2 _405_ (.A(_216_),
    .Y(_051_));
 sky130_fd_sc_hd__inv_2 _406_ (.A(_216_),
    .Y(_052_));
 sky130_fd_sc_hd__inv_2 _407_ (.A(_216_),
    .Y(_053_));
 sky130_fd_sc_hd__inv_2 _408_ (.A(_216_),
    .Y(_054_));
 sky130_fd_sc_hd__inv_2 _409_ (.A(_216_),
    .Y(_055_));
 sky130_fd_sc_hd__buf_1 _410_ (.A(_213_),
    .X(_217_));
 sky130_fd_sc_hd__inv_2 _411_ (.A(_217_),
    .Y(_056_));
 sky130_fd_sc_hd__inv_2 _412_ (.A(_217_),
    .Y(_057_));
 sky130_fd_sc_hd__inv_2 _413_ (.A(_217_),
    .Y(_058_));
 sky130_fd_sc_hd__inv_2 _414_ (.A(_217_),
    .Y(_059_));
 sky130_fd_sc_hd__inv_2 _415_ (.A(_217_),
    .Y(_060_));
 sky130_fd_sc_hd__inv_2 _416_ (.A(_217_),
    .Y(_061_));
 sky130_fd_sc_hd__inv_2 _417_ (.A(_217_),
    .Y(_062_));
 sky130_fd_sc_hd__inv_2 _418_ (.A(_217_),
    .Y(_063_));
 sky130_fd_sc_hd__inv_2 _419_ (.A(_217_),
    .Y(_064_));
 sky130_fd_sc_hd__inv_2 _420_ (.A(_217_),
    .Y(_065_));
 sky130_fd_sc_hd__buf_1 _421_ (.A(wb_rst_i),
    .X(_218_));
 sky130_fd_sc_hd__inv_2 _422_ (.A(_218_),
    .Y(_066_));
 sky130_fd_sc_hd__inv_2 _423_ (.A(_218_),
    .Y(_067_));
 sky130_fd_sc_hd__inv_2 _424_ (.A(_218_),
    .Y(_068_));
 sky130_fd_sc_hd__inv_2 _425_ (.A(_218_),
    .Y(_069_));
 sky130_fd_sc_hd__inv_2 _426_ (.A(_218_),
    .Y(_070_));
 sky130_fd_sc_hd__inv_2 _427_ (.A(_218_),
    .Y(_071_));
 sky130_fd_sc_hd__inv_2 _428_ (.A(_218_),
    .Y(_072_));
 sky130_fd_sc_hd__inv_2 _429_ (.A(_218_),
    .Y(_073_));
 sky130_fd_sc_hd__inv_2 _430_ (.A(_218_),
    .Y(_074_));
 sky130_fd_sc_hd__inv_2 _431_ (.A(_218_),
    .Y(_075_));
 sky130_fd_sc_hd__inv_2 _432_ (.A(_213_),
    .Y(_076_));
 sky130_fd_sc_hd__inv_2 _433_ (.A(_213_),
    .Y(_077_));
 sky130_fd_sc_hd__inv_2 _434_ (.A(_213_),
    .Y(_078_));
 sky130_fd_sc_hd__inv_2 _435_ (.A(_213_),
    .Y(_079_));
 sky130_fd_sc_hd__inv_2 _436_ (.A(_213_),
    .Y(_080_));
 sky130_fd_sc_hd__inv_2 _437_ (.A(_213_),
    .Y(_081_));
 sky130_fd_sc_hd__dfrtp_2 _438_ (.CLK(wb_clk_i),
    .D(_082_),
    .RESET_B(_026_),
    .Q(io_out[24]));
 sky130_fd_sc_hd__dfrtp_2 _439_ (.CLK(wb_clk_i),
    .D(_083_),
    .RESET_B(_027_),
    .Q(io_out[25]));
 sky130_fd_sc_hd__dfrtp_2 _440_ (.CLK(wb_clk_i),
    .D(_084_),
    .RESET_B(_028_),
    .Q(io_out[26]));
 sky130_fd_sc_hd__dfrtp_2 _441_ (.CLK(wb_clk_i),
    .D(_085_),
    .RESET_B(_029_),
    .Q(io_out[27]));
 sky130_fd_sc_hd__dfrtp_2 _442_ (.CLK(wb_clk_i),
    .D(_086_),
    .RESET_B(_030_),
    .Q(io_out[28]));
 sky130_fd_sc_hd__dfrtp_2 _443_ (.CLK(wb_clk_i),
    .D(_087_),
    .RESET_B(_031_),
    .Q(io_out[29]));
 sky130_fd_sc_hd__dfrtp_2 _444_ (.CLK(wb_clk_i),
    .D(_088_),
    .RESET_B(_032_),
    .Q(io_out[30]));
 sky130_fd_sc_hd__dfrtp_2 _445_ (.CLK(wb_clk_i),
    .D(_089_),
    .RESET_B(_033_),
    .Q(io_out[31]));
 sky130_fd_sc_hd__dfrtp_2 _446_ (.CLK(wb_clk_i),
    .D(_090_),
    .RESET_B(_034_),
    .Q(io_out[32]));
 sky130_fd_sc_hd__dfrtp_2 _447_ (.CLK(wb_clk_i),
    .D(_091_),
    .RESET_B(_035_),
    .Q(io_out[33]));
 sky130_fd_sc_hd__dfrtp_2 _448_ (.CLK(wb_clk_i),
    .D(_092_),
    .RESET_B(_036_),
    .Q(io_out[34]));
 sky130_fd_sc_hd__dfrtp_2 _449_ (.CLK(wb_clk_i),
    .D(_093_),
    .RESET_B(_037_),
    .Q(io_out[35]));
 sky130_fd_sc_hd__dfrtp_2 _450_ (.CLK(wb_clk_i),
    .D(_094_),
    .RESET_B(_038_),
    .Q(io_out[36]));
 sky130_fd_sc_hd__dfrtp_2 _451_ (.CLK(wb_clk_i),
    .D(_095_),
    .RESET_B(_039_),
    .Q(io_out[37]));
 sky130_fd_sc_hd__dfrtp_2 _452_ (.CLK(wb_clk_i),
    .D(_096_),
    .RESET_B(_040_),
    .Q(\u_cpu.ALUResult_E[16] ));
 sky130_fd_sc_hd__dfrtp_2 _453_ (.CLK(wb_clk_i),
    .D(_097_),
    .RESET_B(_041_),
    .Q(\u_cpu.ALUResult_E[17] ));
 sky130_fd_sc_hd__dfrtp_2 _454_ (.CLK(wb_clk_i),
    .D(_098_),
    .RESET_B(_042_),
    .Q(\u_cpu.ALUResult_E[18] ));
 sky130_fd_sc_hd__dfrtp_2 _455_ (.CLK(wb_clk_i),
    .D(_099_),
    .RESET_B(_043_),
    .Q(\u_cpu.ALUResult_E[19] ));
 sky130_fd_sc_hd__dfrtp_2 _456_ (.CLK(wb_clk_i),
    .D(_100_),
    .RESET_B(_044_),
    .Q(\u_cpu.ALUResult_E[20] ));
 sky130_fd_sc_hd__dfrtp_2 _457_ (.CLK(wb_clk_i),
    .D(_101_),
    .RESET_B(_045_),
    .Q(\u_cpu.ALUResult_E[21] ));
 sky130_fd_sc_hd__dfrtp_2 _458_ (.CLK(wb_clk_i),
    .D(_102_),
    .RESET_B(_046_),
    .Q(\u_cpu.ALUResult_E[22] ));
 sky130_fd_sc_hd__dfrtp_2 _459_ (.CLK(wb_clk_i),
    .D(_103_),
    .RESET_B(_047_),
    .Q(\u_cpu.ALUResult_E[23] ));
 sky130_fd_sc_hd__dfrtp_2 _460_ (.CLK(wb_clk_i),
    .D(_104_),
    .RESET_B(_048_),
    .Q(\u_cpu.ALUResult_E[24] ));
 sky130_fd_sc_hd__dfrtp_2 _461_ (.CLK(wb_clk_i),
    .D(_105_),
    .RESET_B(_049_),
    .Q(\u_cpu.ALUResult_E[25] ));
 sky130_fd_sc_hd__dfrtp_2 _462_ (.CLK(wb_clk_i),
    .D(_106_),
    .RESET_B(_050_),
    .Q(\u_cpu.ALUResult_E[26] ));
 sky130_fd_sc_hd__dfrtp_2 _463_ (.CLK(wb_clk_i),
    .D(_107_),
    .RESET_B(_051_),
    .Q(\u_cpu.ALUResult_E[27] ));
 sky130_fd_sc_hd__dfrtp_2 _464_ (.CLK(wb_clk_i),
    .D(_108_),
    .RESET_B(_052_),
    .Q(\u_cpu.ALUResult_E[28] ));
 sky130_fd_sc_hd__dfrtp_2 _465_ (.CLK(wb_clk_i),
    .D(_109_),
    .RESET_B(_053_),
    .Q(\u_cpu.ALUResult_E[29] ));
 sky130_fd_sc_hd__dfrtp_2 _466_ (.CLK(wb_clk_i),
    .D(_110_),
    .RESET_B(_054_),
    .Q(\u_cpu.ALUResult_E[30] ));
 sky130_fd_sc_hd__dfrtp_2 _467_ (.CLK(wb_clk_i),
    .D(_111_),
    .RESET_B(_055_),
    .Q(\u_cpu.ALUResult_E[31] ));
 sky130_fd_sc_hd__dfrtp_2 _468_ (.CLK(wb_clk_i),
    .D(_000_),
    .RESET_B(_056_),
    .Q(\u_cpu.counter[0] ));
 sky130_fd_sc_hd__dfrtp_2 _469_ (.CLK(wb_clk_i),
    .D(_011_),
    .RESET_B(_057_),
    .Q(\u_cpu.counter[1] ));
 sky130_fd_sc_hd__dfrtp_2 _470_ (.CLK(wb_clk_i),
    .D(_018_),
    .RESET_B(_058_),
    .Q(\u_cpu.counter[2] ));
 sky130_fd_sc_hd__dfrtp_2 _471_ (.CLK(wb_clk_i),
    .D(_019_),
    .RESET_B(_059_),
    .Q(\u_cpu.counter[3] ));
 sky130_fd_sc_hd__dfrtp_2 _472_ (.CLK(wb_clk_i),
    .D(_020_),
    .RESET_B(_060_),
    .Q(\u_cpu.counter[4] ));
 sky130_fd_sc_hd__dfrtp_2 _473_ (.CLK(wb_clk_i),
    .D(_021_),
    .RESET_B(_061_),
    .Q(\u_cpu.counter[5] ));
 sky130_fd_sc_hd__dfrtp_2 _474_ (.CLK(wb_clk_i),
    .D(_022_),
    .RESET_B(_062_),
    .Q(\u_cpu.counter[6] ));
 sky130_fd_sc_hd__dfrtp_2 _475_ (.CLK(wb_clk_i),
    .D(_023_),
    .RESET_B(_063_),
    .Q(\u_cpu.counter[7] ));
 sky130_fd_sc_hd__dfrtp_2 _476_ (.CLK(wb_clk_i),
    .D(_024_),
    .RESET_B(_064_),
    .Q(\u_cpu.counter[8] ));
 sky130_fd_sc_hd__dfrtp_2 _477_ (.CLK(wb_clk_i),
    .D(_025_),
    .RESET_B(_065_),
    .Q(\u_cpu.counter[9] ));
 sky130_fd_sc_hd__dfrtp_2 _478_ (.CLK(wb_clk_i),
    .D(_001_),
    .RESET_B(_066_),
    .Q(\u_cpu.counter[10] ));
 sky130_fd_sc_hd__dfrtp_2 _479_ (.CLK(wb_clk_i),
    .D(_002_),
    .RESET_B(_067_),
    .Q(\u_cpu.counter[11] ));
 sky130_fd_sc_hd__dfrtp_2 _480_ (.CLK(wb_clk_i),
    .D(_003_),
    .RESET_B(_068_),
    .Q(\u_cpu.counter[12] ));
 sky130_fd_sc_hd__dfrtp_2 _481_ (.CLK(wb_clk_i),
    .D(_004_),
    .RESET_B(_069_),
    .Q(\u_cpu.counter[13] ));
 sky130_fd_sc_hd__dfrtp_2 _482_ (.CLK(wb_clk_i),
    .D(_005_),
    .RESET_B(_070_),
    .Q(\u_cpu.counter[14] ));
 sky130_fd_sc_hd__dfrtp_2 _483_ (.CLK(wb_clk_i),
    .D(_006_),
    .RESET_B(_071_),
    .Q(\u_cpu.counter[15] ));
 sky130_fd_sc_hd__dfrtp_2 _484_ (.CLK(wb_clk_i),
    .D(_007_),
    .RESET_B(_072_),
    .Q(\u_cpu.counter[16] ));
 sky130_fd_sc_hd__dfrtp_2 _485_ (.CLK(wb_clk_i),
    .D(_008_),
    .RESET_B(_073_),
    .Q(\u_cpu.counter[17] ));
 sky130_fd_sc_hd__dfrtp_2 _486_ (.CLK(wb_clk_i),
    .D(_009_),
    .RESET_B(_074_),
    .Q(\u_cpu.counter[18] ));
 sky130_fd_sc_hd__dfrtp_2 _487_ (.CLK(wb_clk_i),
    .D(_010_),
    .RESET_B(_075_),
    .Q(\u_cpu.counter[19] ));
 sky130_fd_sc_hd__dfrtp_2 _488_ (.CLK(wb_clk_i),
    .D(_012_),
    .RESET_B(_076_),
    .Q(\u_cpu.counter[20] ));
 sky130_fd_sc_hd__dfrtp_2 _489_ (.CLK(wb_clk_i),
    .D(_013_),
    .RESET_B(_077_),
    .Q(\u_cpu.counter[21] ));
 sky130_fd_sc_hd__dfrtp_2 _490_ (.CLK(wb_clk_i),
    .D(_014_),
    .RESET_B(_078_),
    .Q(\u_cpu.counter[22] ));
 sky130_fd_sc_hd__dfrtp_2 _491_ (.CLK(wb_clk_i),
    .D(_015_),
    .RESET_B(_079_),
    .Q(\u_cpu.counter[23] ));
 sky130_fd_sc_hd__dfrtp_2 _492_ (.CLK(wb_clk_i),
    .D(_016_),
    .RESET_B(_080_),
    .Q(\u_cpu.counter[24] ));
 sky130_fd_sc_hd__dfrtp_2 _493_ (.CLK(wb_clk_i),
    .D(_017_),
    .RESET_B(_081_),
    .Q(\u_cpu.counter[25] ));
 sky130_fd_sc_hd__conb_1 _494_ (.LO(io_oeb[0]));
 sky130_fd_sc_hd__conb_1 _495_ (.LO(io_oeb[1]));
 sky130_fd_sc_hd__conb_1 _496_ (.LO(io_oeb[2]));
 sky130_fd_sc_hd__conb_1 _497_ (.LO(io_oeb[3]));
 sky130_fd_sc_hd__conb_1 _498_ (.LO(io_oeb[4]));
 sky130_fd_sc_hd__conb_1 _499_ (.LO(io_oeb[5]));
 sky130_fd_sc_hd__conb_1 _500_ (.LO(io_oeb[6]));
 sky130_fd_sc_hd__conb_1 _501_ (.LO(io_oeb[7]));
 sky130_fd_sc_hd__conb_1 _502_ (.LO(io_oeb[8]));
 sky130_fd_sc_hd__conb_1 _503_ (.LO(io_oeb[9]));
 sky130_fd_sc_hd__conb_1 _504_ (.LO(io_oeb[10]));
 sky130_fd_sc_hd__conb_1 _505_ (.LO(io_oeb[11]));
 sky130_fd_sc_hd__conb_1 _506_ (.LO(io_oeb[12]));
 sky130_fd_sc_hd__conb_1 _507_ (.LO(io_oeb[13]));
 sky130_fd_sc_hd__conb_1 _508_ (.LO(io_oeb[14]));
 sky130_fd_sc_hd__conb_1 _509_ (.LO(io_oeb[15]));
 sky130_fd_sc_hd__conb_1 _510_ (.LO(io_oeb[16]));
 sky130_fd_sc_hd__conb_1 _511_ (.LO(io_oeb[17]));
 sky130_fd_sc_hd__conb_1 _512_ (.LO(io_oeb[18]));
 sky130_fd_sc_hd__conb_1 _513_ (.LO(io_oeb[19]));
 sky130_fd_sc_hd__conb_1 _514_ (.LO(io_oeb[20]));
 sky130_fd_sc_hd__conb_1 _515_ (.LO(io_oeb[21]));
 sky130_fd_sc_hd__conb_1 _516_ (.LO(io_oeb[22]));
 sky130_fd_sc_hd__conb_1 _517_ (.LO(io_oeb[23]));
 sky130_fd_sc_hd__conb_1 _518_ (.LO(io_oeb[24]));
 sky130_fd_sc_hd__conb_1 _519_ (.LO(io_oeb[25]));
 sky130_fd_sc_hd__conb_1 _520_ (.LO(io_oeb[26]));
 sky130_fd_sc_hd__conb_1 _521_ (.LO(io_oeb[27]));
 sky130_fd_sc_hd__conb_1 _522_ (.LO(io_oeb[28]));
 sky130_fd_sc_hd__conb_1 _523_ (.LO(io_oeb[29]));
 sky130_fd_sc_hd__conb_1 _524_ (.LO(io_oeb[30]));
 sky130_fd_sc_hd__conb_1 _525_ (.LO(io_oeb[31]));
 sky130_fd_sc_hd__conb_1 _526_ (.LO(io_oeb[32]));
 sky130_fd_sc_hd__conb_1 _527_ (.LO(io_oeb[33]));
 sky130_fd_sc_hd__conb_1 _528_ (.LO(io_oeb[34]));
 sky130_fd_sc_hd__conb_1 _529_ (.LO(io_oeb[35]));
 sky130_fd_sc_hd__conb_1 _530_ (.LO(io_oeb[36]));
 sky130_fd_sc_hd__conb_1 _531_ (.LO(io_oeb[37]));
 sky130_fd_sc_hd__conb_1 _532_ (.LO(io_out[0]));
 sky130_fd_sc_hd__conb_1 _533_ (.LO(io_out[1]));
 sky130_fd_sc_hd__conb_1 _534_ (.LO(io_out[10]));
 sky130_fd_sc_hd__conb_1 _535_ (.LO(io_out[11]));
 sky130_fd_sc_hd__conb_1 _536_ (.LO(io_out[12]));
 sky130_fd_sc_hd__conb_1 _537_ (.LO(io_out[13]));
 sky130_fd_sc_hd__conb_1 _538_ (.LO(io_out[14]));
 sky130_fd_sc_hd__conb_1 _539_ (.LO(io_out[15]));
 sky130_fd_sc_hd__conb_1 _540_ (.LO(io_out[16]));
 sky130_fd_sc_hd__conb_1 _541_ (.LO(io_out[17]));
 sky130_fd_sc_hd__conb_1 _542_ (.LO(io_out[18]));
 sky130_fd_sc_hd__conb_1 _543_ (.LO(io_out[19]));
 sky130_fd_sc_hd__conb_1 _544_ (.LO(io_out[20]));
 sky130_fd_sc_hd__conb_1 _545_ (.LO(io_out[21]));
 sky130_fd_sc_hd__conb_1 _546_ (.LO(io_out[22]));
 sky130_fd_sc_hd__conb_1 _547_ (.LO(io_out[23]));
 sky130_fd_sc_hd__conb_1 _548_ (.LO(\u_cpu.ALUResult_E[0] ));
 sky130_fd_sc_hd__conb_1 _549_ (.LO(\u_cpu.ALUResult_E[1] ));
 sky130_fd_sc_hd__conb_1 _550_ (.LO(\u_cpu.Instr_D[0] ));
 sky130_fd_sc_hd__conb_1 _551_ (.LO(\u_cpu.Instr_D[1] ));
 sky130_fd_sc_hd__conb_1 _552_ (.LO(\u_cpu.Instr_D[2] ));
 sky130_fd_sc_hd__conb_1 _553_ (.LO(\u_cpu.Instr_D[3] ));
 sky130_fd_sc_hd__conb_1 _554_ (.LO(\u_cpu.Instr_D[4] ));
 sky130_fd_sc_hd__conb_1 _555_ (.LO(\u_cpu.Instr_D[5] ));
 sky130_fd_sc_hd__conb_1 _556_ (.LO(\u_cpu.Instr_D[6] ));
 sky130_fd_sc_hd__conb_1 _557_ (.LO(\u_cpu.Instr_D[7] ));
 sky130_fd_sc_hd__conb_1 _558_ (.LO(\u_cpu.Instr_D[8] ));
 sky130_fd_sc_hd__conb_1 _559_ (.LO(\u_cpu.Instr_D[9] ));
 sky130_fd_sc_hd__conb_1 _560_ (.LO(\u_cpu.Instr_D[10] ));
 sky130_fd_sc_hd__conb_1 _561_ (.LO(\u_cpu.Instr_D[11] ));
 sky130_fd_sc_hd__conb_1 _562_ (.LO(\u_cpu.Instr_D[12] ));
 sky130_fd_sc_hd__conb_1 _563_ (.LO(\u_cpu.Instr_D[13] ));
 sky130_fd_sc_hd__conb_1 _564_ (.LO(\u_cpu.Instr_D[14] ));
 sky130_fd_sc_hd__conb_1 _565_ (.LO(\u_cpu.Instr_D[15] ));
 sky130_fd_sc_hd__conb_1 _566_ (.LO(\u_cpu.Instr_D[16] ));
 sky130_fd_sc_hd__conb_1 _567_ (.LO(\u_cpu.Instr_D[17] ));
 sky130_fd_sc_hd__conb_1 _568_ (.LO(\u_cpu.Instr_D[18] ));
 sky130_fd_sc_hd__conb_1 _569_ (.LO(\u_cpu.Instr_D[19] ));
 sky130_fd_sc_hd__conb_1 _570_ (.LO(\u_cpu.Instr_D[20] ));
 sky130_fd_sc_hd__conb_1 _571_ (.LO(\u_cpu.Instr_D[21] ));
 sky130_fd_sc_hd__conb_1 _572_ (.LO(\u_cpu.Instr_D[22] ));
 sky130_fd_sc_hd__conb_1 _573_ (.LO(\u_cpu.Instr_D[23] ));
 sky130_fd_sc_hd__conb_1 _574_ (.LO(\u_cpu.Instr_D[24] ));
 sky130_fd_sc_hd__conb_1 _575_ (.LO(\u_cpu.Instr_D[25] ));
 sky130_fd_sc_hd__conb_1 _576_ (.LO(\u_cpu.Instr_D[26] ));
 sky130_fd_sc_hd__conb_1 _577_ (.LO(\u_cpu.Instr_D[27] ));
 sky130_fd_sc_hd__conb_1 _578_ (.LO(\u_cpu.Instr_D[28] ));
 sky130_fd_sc_hd__conb_1 _579_ (.LO(\u_cpu.Instr_D[29] ));
 sky130_fd_sc_hd__conb_1 _580_ (.LO(\u_cpu.Instr_D[30] ));
 sky130_fd_sc_hd__conb_1 _581_ (.LO(\u_cpu.Instr_D[31] ));
 sky130_fd_sc_hd__conb_1 _582_ (.LO(\u_cpu.Instr_F[0] ));
 sky130_fd_sc_hd__conb_1 _583_ (.LO(\u_cpu.Instr_F[1] ));
 sky130_fd_sc_hd__conb_1 _584_ (.LO(\u_cpu.Instr_F[2] ));
 sky130_fd_sc_hd__conb_1 _585_ (.LO(\u_cpu.Instr_F[3] ));
 sky130_fd_sc_hd__conb_1 _586_ (.LO(\u_cpu.Instr_F[4] ));
 sky130_fd_sc_hd__conb_1 _587_ (.LO(\u_cpu.Instr_F[5] ));
 sky130_fd_sc_hd__conb_1 _588_ (.LO(\u_cpu.Instr_F[6] ));
 sky130_fd_sc_hd__conb_1 _589_ (.LO(\u_cpu.Instr_F[7] ));
 sky130_fd_sc_hd__conb_1 _590_ (.LO(\u_cpu.Instr_F[8] ));
 sky130_fd_sc_hd__conb_1 _591_ (.LO(\u_cpu.Instr_F[9] ));
 sky130_fd_sc_hd__conb_1 _592_ (.LO(\u_cpu.Instr_F[10] ));
 sky130_fd_sc_hd__conb_1 _593_ (.LO(\u_cpu.Instr_F[11] ));
 sky130_fd_sc_hd__conb_1 _594_ (.LO(\u_cpu.Instr_F[12] ));
 sky130_fd_sc_hd__conb_1 _595_ (.LO(\u_cpu.Instr_F[13] ));
 sky130_fd_sc_hd__conb_1 _596_ (.LO(\u_cpu.Instr_F[14] ));
 sky130_fd_sc_hd__conb_1 _597_ (.LO(\u_cpu.Instr_F[15] ));
 sky130_fd_sc_hd__conb_1 _598_ (.LO(\u_cpu.Instr_F[16] ));
 sky130_fd_sc_hd__conb_1 _599_ (.LO(\u_cpu.Instr_F[17] ));
 sky130_fd_sc_hd__conb_1 _600_ (.LO(\u_cpu.Instr_F[18] ));
 sky130_fd_sc_hd__conb_1 _601_ (.LO(\u_cpu.Instr_F[19] ));
 sky130_fd_sc_hd__conb_1 _602_ (.LO(\u_cpu.Instr_F[20] ));
 sky130_fd_sc_hd__conb_1 _603_ (.LO(\u_cpu.Instr_F[21] ));
 sky130_fd_sc_hd__conb_1 _604_ (.LO(\u_cpu.Instr_F[22] ));
 sky130_fd_sc_hd__conb_1 _605_ (.LO(\u_cpu.Instr_F[23] ));
 sky130_fd_sc_hd__conb_1 _606_ (.LO(\u_cpu.Instr_F[24] ));
 sky130_fd_sc_hd__conb_1 _607_ (.LO(\u_cpu.Instr_F[25] ));
 sky130_fd_sc_hd__conb_1 _608_ (.LO(\u_cpu.Instr_F[26] ));
 sky130_fd_sc_hd__conb_1 _609_ (.LO(\u_cpu.Instr_F[27] ));
 sky130_fd_sc_hd__conb_1 _610_ (.LO(\u_cpu.Instr_F[28] ));
 sky130_fd_sc_hd__conb_1 _611_ (.LO(\u_cpu.Instr_F[29] ));
 sky130_fd_sc_hd__conb_1 _612_ (.LO(\u_cpu.Instr_F[30] ));
 sky130_fd_sc_hd__conb_1 _613_ (.LO(\u_cpu.Instr_F[31] ));
 sky130_fd_sc_hd__conb_1 _614_ (.LO(\u_cpu.PC_F[0] ));
 sky130_fd_sc_hd__conb_1 _615_ (.LO(\u_cpu.PC_F[1] ));
 sky130_fd_sc_hd__buf_2 _616_ (.A(io_out[26]),
    .X(\u_cpu.ALUResult_E[4] ));
 sky130_fd_sc_hd__buf_2 _617_ (.A(io_out[27]),
    .X(\u_cpu.ALUResult_E[5] ));
 sky130_fd_sc_hd__buf_2 _618_ (.A(io_out[28]),
    .X(\u_cpu.ALUResult_E[6] ));
 sky130_fd_sc_hd__buf_2 _619_ (.A(io_out[29]),
    .X(\u_cpu.ALUResult_E[7] ));
 sky130_fd_sc_hd__buf_2 _620_ (.A(io_out[30]),
    .X(\u_cpu.ALUResult_E[8] ));
 sky130_fd_sc_hd__buf_2 _621_ (.A(io_out[31]),
    .X(\u_cpu.ALUResult_E[9] ));
 sky130_fd_sc_hd__buf_2 _622_ (.A(io_out[32]),
    .X(\u_cpu.ALUResult_E[10] ));
 sky130_fd_sc_hd__buf_2 _623_ (.A(io_out[33]),
    .X(\u_cpu.ALUResult_E[11] ));
 sky130_fd_sc_hd__buf_2 _624_ (.A(io_out[34]),
    .X(\u_cpu.ALUResult_E[12] ));
 sky130_fd_sc_hd__buf_2 _625_ (.A(io_out[35]),
    .X(\u_cpu.ALUResult_E[13] ));
 sky130_fd_sc_hd__buf_2 _626_ (.A(io_out[36]),
    .X(\u_cpu.ALUResult_E[14] ));
 sky130_fd_sc_hd__buf_2 _627_ (.A(io_out[37]),
    .X(\u_cpu.ALUResult_E[15] ));
 sky130_fd_sc_hd__buf_2 _628_ (.A(io_out[24]),
    .X(\u_cpu.PC_F[2] ));
 sky130_fd_sc_hd__buf_2 _629_ (.A(io_out[25]),
    .X(\u_cpu.PC_F[3] ));
 sky130_fd_sc_hd__buf_2 _630_ (.A(io_out[26]),
    .X(\u_cpu.PC_F[4] ));
 sky130_fd_sc_hd__buf_2 _631_ (.A(io_out[27]),
    .X(\u_cpu.PC_F[5] ));
 sky130_fd_sc_hd__buf_2 _632_ (.A(io_out[28]),
    .X(\u_cpu.PC_F[6] ));
 sky130_fd_sc_hd__buf_2 _633_ (.A(io_out[29]),
    .X(\u_cpu.PC_F[7] ));
 sky130_fd_sc_hd__buf_2 _634_ (.A(io_out[30]),
    .X(\u_cpu.PC_F[8] ));
 sky130_fd_sc_hd__buf_2 _635_ (.A(io_out[31]),
    .X(\u_cpu.PC_F[9] ));
 sky130_fd_sc_hd__buf_2 _636_ (.A(io_out[32]),
    .X(\u_cpu.PC_F[10] ));
 sky130_fd_sc_hd__buf_2 _637_ (.A(io_out[33]),
    .X(\u_cpu.PC_F[11] ));
 sky130_fd_sc_hd__buf_2 _638_ (.A(io_out[34]),
    .X(\u_cpu.PC_F[12] ));
 sky130_fd_sc_hd__buf_2 _639_ (.A(io_out[35]),
    .X(\u_cpu.PC_F[13] ));
 sky130_fd_sc_hd__buf_2 _640_ (.A(io_out[36]),
    .X(\u_cpu.PC_F[14] ));
 sky130_fd_sc_hd__buf_2 _641_ (.A(io_out[37]),
    .X(\u_cpu.PC_F[15] ));
 sky130_fd_sc_hd__buf_2 _642_ (.A(\u_cpu.ALUResult_E[16] ),
    .X(\u_cpu.PC_F[16] ));
 sky130_fd_sc_hd__buf_2 _643_ (.A(\u_cpu.ALUResult_E[17] ),
    .X(\u_cpu.PC_F[17] ));
 sky130_fd_sc_hd__buf_2 _644_ (.A(\u_cpu.ALUResult_E[18] ),
    .X(\u_cpu.PC_F[18] ));
 sky130_fd_sc_hd__buf_2 _645_ (.A(\u_cpu.ALUResult_E[19] ),
    .X(\u_cpu.PC_F[19] ));
 sky130_fd_sc_hd__buf_2 _646_ (.A(\u_cpu.ALUResult_E[20] ),
    .X(\u_cpu.PC_F[20] ));
 sky130_fd_sc_hd__buf_2 _647_ (.A(\u_cpu.ALUResult_E[21] ),
    .X(\u_cpu.PC_F[21] ));
 sky130_fd_sc_hd__buf_2 _648_ (.A(\u_cpu.ALUResult_E[22] ),
    .X(\u_cpu.PC_F[22] ));
 sky130_fd_sc_hd__buf_2 _649_ (.A(\u_cpu.ALUResult_E[23] ),
    .X(\u_cpu.PC_F[23] ));
 sky130_fd_sc_hd__buf_2 _650_ (.A(\u_cpu.ALUResult_E[24] ),
    .X(\u_cpu.PC_F[24] ));
 sky130_fd_sc_hd__buf_2 _651_ (.A(\u_cpu.ALUResult_E[25] ),
    .X(\u_cpu.PC_F[25] ));
 sky130_fd_sc_hd__buf_2 _652_ (.A(\u_cpu.ALUResult_E[26] ),
    .X(\u_cpu.PC_F[26] ));
 sky130_fd_sc_hd__buf_2 _653_ (.A(\u_cpu.ALUResult_E[27] ),
    .X(\u_cpu.PC_F[27] ));
 sky130_fd_sc_hd__buf_2 _654_ (.A(\u_cpu.ALUResult_E[28] ),
    .X(\u_cpu.PC_F[28] ));
 sky130_fd_sc_hd__buf_2 _655_ (.A(\u_cpu.ALUResult_E[29] ),
    .X(\u_cpu.PC_F[29] ));
 sky130_fd_sc_hd__buf_2 _656_ (.A(\u_cpu.ALUResult_E[30] ),
    .X(\u_cpu.PC_F[30] ));
 sky130_fd_sc_hd__buf_2 _657_ (.A(\u_cpu.ALUResult_E[31] ),
    .X(\u_cpu.PC_F[31] ));
 sky130_fd_sc_hd__buf_2 _658_ (.A(io_out[24]),
    .X(\u_cpu.ALUResult_E[2] ));
 sky130_fd_sc_hd__buf_2 _659_ (.A(io_out[25]),
    .X(\u_cpu.ALUResult_E[3] ));
 sky130_fd_sc_hd__buf_2 _660_ (.A(io_out[24]),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_2 _661_ (.A(io_out[25]),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_2 _662_ (.A(io_out[26]),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_2 _663_ (.A(io_out[27]),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_2 _664_ (.A(io_out[28]),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_2 _665_ (.A(io_out[29]),
    .X(io_out[7]));
 sky130_fd_sc_hd__buf_2 _666_ (.A(io_out[30]),
    .X(io_out[8]));
 sky130_fd_sc_hd__buf_2 _667_ (.A(io_out[31]),
    .X(io_out[9]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__decap_3 PHY_572 ();
 sky130_fd_sc_hd__decap_3 PHY_573 ();
 sky130_fd_sc_hd__decap_3 PHY_574 ();
 sky130_fd_sc_hd__decap_3 PHY_575 ();
 sky130_fd_sc_hd__decap_3 PHY_576 ();
 sky130_fd_sc_hd__decap_3 PHY_577 ();
 sky130_fd_sc_hd__decap_3 PHY_578 ();
 sky130_fd_sc_hd__decap_3 PHY_579 ();
 sky130_fd_sc_hd__decap_3 PHY_580 ();
 sky130_fd_sc_hd__decap_3 PHY_581 ();
 sky130_fd_sc_hd__decap_3 PHY_582 ();
 sky130_fd_sc_hd__decap_3 PHY_583 ();
 sky130_fd_sc_hd__decap_3 PHY_584 ();
 sky130_fd_sc_hd__decap_3 PHY_585 ();
 sky130_fd_sc_hd__decap_3 PHY_586 ();
 sky130_fd_sc_hd__decap_3 PHY_587 ();
 sky130_fd_sc_hd__decap_3 PHY_588 ();
 sky130_fd_sc_hd__decap_3 PHY_589 ();
 sky130_fd_sc_hd__decap_3 PHY_590 ();
 sky130_fd_sc_hd__decap_3 PHY_591 ();
 sky130_fd_sc_hd__decap_3 PHY_592 ();
 sky130_fd_sc_hd__decap_3 PHY_593 ();
 sky130_fd_sc_hd__decap_3 PHY_594 ();
 sky130_fd_sc_hd__decap_3 PHY_595 ();
 sky130_fd_sc_hd__decap_3 PHY_596 ();
 sky130_fd_sc_hd__decap_3 PHY_597 ();
 sky130_fd_sc_hd__decap_3 PHY_598 ();
 sky130_fd_sc_hd__decap_3 PHY_599 ();
 sky130_fd_sc_hd__decap_3 PHY_600 ();
 sky130_fd_sc_hd__decap_3 PHY_601 ();
 sky130_fd_sc_hd__decap_3 PHY_602 ();
 sky130_fd_sc_hd__decap_3 PHY_603 ();
 sky130_fd_sc_hd__decap_3 PHY_604 ();
 sky130_fd_sc_hd__decap_3 PHY_605 ();
 sky130_fd_sc_hd__decap_3 PHY_606 ();
 sky130_fd_sc_hd__decap_3 PHY_607 ();
 sky130_fd_sc_hd__decap_3 PHY_608 ();
 sky130_fd_sc_hd__decap_3 PHY_609 ();
 sky130_fd_sc_hd__decap_3 PHY_610 ();
 sky130_fd_sc_hd__decap_3 PHY_611 ();
 sky130_fd_sc_hd__decap_3 PHY_612 ();
 sky130_fd_sc_hd__decap_3 PHY_613 ();
 sky130_fd_sc_hd__decap_3 PHY_614 ();
 sky130_fd_sc_hd__decap_3 PHY_615 ();
 sky130_fd_sc_hd__decap_3 PHY_616 ();
 sky130_fd_sc_hd__decap_3 PHY_617 ();
 sky130_fd_sc_hd__decap_3 PHY_618 ();
 sky130_fd_sc_hd__decap_3 PHY_619 ();
 sky130_fd_sc_hd__decap_3 PHY_620 ();
 sky130_fd_sc_hd__decap_3 PHY_621 ();
 sky130_fd_sc_hd__decap_3 PHY_622 ();
 sky130_fd_sc_hd__decap_3 PHY_623 ();
 sky130_fd_sc_hd__decap_3 PHY_624 ();
 sky130_fd_sc_hd__decap_3 PHY_625 ();
 sky130_fd_sc_hd__decap_3 PHY_626 ();
 sky130_fd_sc_hd__decap_3 PHY_627 ();
 sky130_fd_sc_hd__decap_3 PHY_628 ();
 sky130_fd_sc_hd__decap_3 PHY_629 ();
 sky130_fd_sc_hd__decap_3 PHY_630 ();
 sky130_fd_sc_hd__decap_3 PHY_631 ();
 sky130_fd_sc_hd__decap_3 PHY_632 ();
 sky130_fd_sc_hd__decap_3 PHY_633 ();
 sky130_fd_sc_hd__decap_3 PHY_634 ();
 sky130_fd_sc_hd__decap_3 PHY_635 ();
 sky130_fd_sc_hd__decap_3 PHY_636 ();
 sky130_fd_sc_hd__decap_3 PHY_637 ();
 sky130_fd_sc_hd__decap_3 PHY_638 ();
 sky130_fd_sc_hd__decap_3 PHY_639 ();
 sky130_fd_sc_hd__decap_3 PHY_640 ();
 sky130_fd_sc_hd__decap_3 PHY_641 ();
 sky130_fd_sc_hd__decap_3 PHY_642 ();
 sky130_fd_sc_hd__decap_3 PHY_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11659 ();
endmodule
