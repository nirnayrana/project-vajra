
.SUBCKT sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 y VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inor VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inor pmid VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 y VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inor VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inor pmid VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 y VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inor VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inor pmid VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 Y VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inor VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inor pmid VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 Y VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inor VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inor pmid VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 Y VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inor VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inor pmid VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA20 y A1 snd2A1 VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA21 snd2A1 A2 VGND VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21boi_0 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 net40 A1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 net40 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 net40 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 net40 A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 net40 A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 net40 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 net40 A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 net40 A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 net40 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 net40 A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 net40 A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 net40 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA20 y A1 snd2A1 VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA21 snd2A1 A2 VGND VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB20 pnd2B B1 pndA VPB pfet_01v8_hvt w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC20 y C1 pnd2B VPB pfet_01v8_hvt w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA20 y A1 snd2A1 VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA21 snd2A1 A2 VGND VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a222oi_1 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 Y C2 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 net62 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net62 C2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 y D1 pndC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 y D1 pndC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 y D1 pndC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111oi_0 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 Y D1 pndC VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 Y D1 pndC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 Y D1 pndC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 Y D1 pndC VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2_0 A B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=12 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=12 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_16 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__bufbuf_8 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 Abb Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 Abbb Abb VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X Abbb VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X Abbb VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Abbb Abb VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__bufbuf_16 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 Abb Ab VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 Abbb Abb VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X Abbb VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X Abbb VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 Abb Ab VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Abbb Abb VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__bufinv_8 A VGND VNB VPB VPWR Y
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 Abb Ab VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 Y Abb VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 Abb Ab VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 Y Abb VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
MMIN1 Ab A VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 Abb Ab VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 Y Abb VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 Abb Ab VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 Y Abb VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=8 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s15_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s15_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s18_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s18_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s25_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s50_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=8 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=12 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=24 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net36 A VGND VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 Y A net36 VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 Y A net31 VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net35 A VGND VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net31 A VGND VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Y A net35 VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
rI12 VGND LO sky130_fd_pr__res_generic_po
rI11 HI VPWR sky130_fd_pr__res_generic_po
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=0.59 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=0.59 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=1.05 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=1.05 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=1.97 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=1.97 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=2.89 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=2.89 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=4.73 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=4.73 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfbbn_1 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net141 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net162 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net125 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net125 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net110 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net82 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net162 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net93 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net93 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net82 RESET net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net82 S0 net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net81 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net218 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net162 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net82 S0 net221 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net218 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net165 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net210 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net210 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net82 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net221 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net165 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net162 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net82 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfbbn_2 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net141 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net162 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net125 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net125 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net110 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net82 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net162 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net93 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net93 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net82 RESET net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net82 S0 net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net81 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net218 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net162 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net82 S0 net221 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net218 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net165 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net210 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net210 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net82 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net221 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net165 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net162 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net82 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfbbp_1 CLK D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net141 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net162 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net118 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net118 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net110 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net82 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net162 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net93 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net93 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net82 RESET net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net82 S0 net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net81 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net218 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net162 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net82 S0 net221 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net218 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net165 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net210 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net210 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net82 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net221 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net165 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net162 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net82 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net99 s0 net125 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net125 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net118 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net110 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net110 M1 net118 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net98 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net99 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net98 net99 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI53 net142 net99 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 Q_N net142 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net190 net99 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net99 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net190 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net99 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net169 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net169 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net169 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net99 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI52 net142 net99 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI51 Q_N net142 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net99 s0 net125 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net125 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net118 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net110 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net110 M1 net118 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net98 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net99 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net98 net99 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI53 net142 net99 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 Q_N net142 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net181 net99 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net99 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net181 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net99 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net169 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net169 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net169 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net99 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI52 net142 net99 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI51 Q_N net142 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net83 net121 net109 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net109 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net102 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net94 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net94 M1 net102 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 net121 clkneg net82 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net83 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net82 net83 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos net121 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net166 net83 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net83 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 net121 clkpos net166 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net83 net121 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net145 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net145 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net145 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net83 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg net121 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net82 s0 net108 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net101 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net93 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net93 M1 net101 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net81 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net82 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net81 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net165 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net82 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net165 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net82 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net144 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net144 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net144 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net82 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net82 s0 net108 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net101 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net93 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net93 M1 net101 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net81 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net82 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net81 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net156 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net82 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net82 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net144 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net144 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net144 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net82 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net82 s0 net108 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net101 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net93 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net93 M1 net101 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net81 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net82 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net81 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net165 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net82 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net165 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net82 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net144 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net144 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net144 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net82 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfsbp_1 CLK D SET_B VGND VNB VPB VPWR Q Q_N
MI36 net129 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net112 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net80 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net129 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net97 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net89 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net89 S1 net97 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net80 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net112 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net141 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net141 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 Q_N S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net192 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net192 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net169 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net169 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net156 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net141 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net141 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 Q_N S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfsbp_2 CLK D SET_B VGND VNB VPB VPWR Q Q_N
MI36 net128 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net111 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net79 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net128 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net96 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net88 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net88 S1 net96 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net79 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net111 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net140 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net140 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 Q_N S0 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net191 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net191 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net168 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net168 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net155 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net140 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net140 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 Q_N S0 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
MI36 net120 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net103 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net71 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net120 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net88 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net80 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net80 S1 net88 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net71 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net103 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net128 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net128 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net179 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net179 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net156 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net143 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net143 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net128 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net128 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
MI36 net120 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net103 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net71 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net120 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net88 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net80 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net80 S1 net88 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net71 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net103 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net128 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net128 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net179 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net179 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net156 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net143 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net143 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net128 S0 VPWR VPB pfet_01v8_hvt m=1 w=1 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net128 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
MI36 net120 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net103 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net71 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net120 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net88 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net80 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net80 S1 net88 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net71 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net103 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net128 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net128 VGND VNB nfet_01v8 m=5 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net179 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net179 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net156 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net143 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net143 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net128 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net128 VPWR VPB pfet_01v8_hvt m=5 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxbp_1 CLK D VGND VNB VPB VPWR Q Q_N
MI657 M0 clkpos net96 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net96 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 net88 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net72 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net72 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 Q_N net88 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net128 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net147 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net88 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net147 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net128 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI666 Q_N net88 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxbp_2 CLK D VGND VNB VPB VPWR Q Q_N
MI657 M0 clkpos net96 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net96 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 net88 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net72 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net72 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 Q_N net88 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net128 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net147 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net88 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net147 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net128 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI666 Q_N net88 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
MI657 M0 clkpos net79 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net79 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net59 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net59 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net107 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net107 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
MI657 M0 clkpos net79 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net79 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net59 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net59 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net107 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net107 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
MI657 M0 clkpos net79 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net79 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net59 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net59 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net107 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net107 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
MI662 net75 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net75 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net63 CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net63 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net54 GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net63 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net110 VNB special_nfet_01v8 m=1 w=0.39 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 M0 clkpos net91 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net99 CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net63 m1 net99 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net91 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net63 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlclkp_2 CLK GATE VGND VNB VPB VPWR GCLK
MI662 net75 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net75 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net63 CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net63 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net54 GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net63 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net110 VNB special_nfet_01v8 m=1 w=0.39 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 M0 clkpos net91 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net99 CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net63 m1 net99 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net91 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net63 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlclkp_4 CLK GATE VGND VNB VPB VPWR GCLK
MI662 net75 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net75 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net63 CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net63 m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net54 GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net63 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net110 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 M0 clkpos net91 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net99 CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net63 m1 net99 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net91 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net63 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrbn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net125 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net61 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net125 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net61 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net57 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net57 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net125 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net125 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net116 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net116 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net108 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net96 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net96 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrbn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net125 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net61 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net125 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net61 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net57 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net57 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net125 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net125 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net116 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net116 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net108 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net96 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net96 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrbp_1 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net125 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net61 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net125 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net61 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net57 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net57 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net125 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net125 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net121 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net116 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net116 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net121 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net96 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net96 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrbp_2 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net125 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net61 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net125 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net61 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net57 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net57 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net125 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net125 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net116 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net116 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net108 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net96 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net96 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net54 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net50 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net50 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net93 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net101 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net101 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net93 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net81 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net81 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net54 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net50 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net50 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net93 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net101 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net101 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net93 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net81 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net81 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtn_4 D GATE_N RESET_B VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net55 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net55 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net51 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net94 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net102 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net102 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net94 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net82 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net82 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtp_1 D GATE RESET_B VGND VNB VPB VPWR Q
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net54 VPB special_pfet_01v8_hvt m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net54 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net50 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net50 VPB special_pfet_01v8_hvt m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net93 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net101 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net101 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net93 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net81 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net81 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtp_2 D GATE RESET_B VGND VNB VPB VPWR Q
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net54 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net50 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net50 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net93 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net101 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net101 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net93 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net81 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net81 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtp_4 D GATE RESET_B VGND VNB VPB VPWR Q
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net55 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net55 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net51 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net94 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net102 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net102 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net94 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net82 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net82 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxbn_1 D GATE_N VGND VNB VPB VPWR Q Q_N
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net112 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net56 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net112 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net56 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net52 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net52 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net112 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net112 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net107 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net107 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net87 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net87 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxbn_2 D GATE_N VGND VNB VPB VPWR Q Q_N
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net114 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net58 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net114 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net58 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net54 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net114 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net114 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net109 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net109 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net89 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net89 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net114 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net58 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net114 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net58 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net54 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net114 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net114 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net109 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net109 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net89 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net89 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net53 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net53 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net44 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net44 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net96 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net96 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net76 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net76 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net51 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net47 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net47 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net94 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net94 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net74 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net74 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxtn_4 D GATE_N VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net51 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net47 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net47 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net94 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net94 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net74 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net74 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net51 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net47 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net47 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net94 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net94 m1 VGND VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net74 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net74 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
MMIN1 Ab net34 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net34 net30 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net30 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net34 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net34 net30 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net30 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlygate4sd2_1 A VGND VNB VPB VPWR X
MMIN1 Ab net34 VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net34 net30 VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net30 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net34 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.18 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net34 net30 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.18 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net30 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
MMIN1 Ab net34 VGND VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net34 net30 VGND VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net30 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net34 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net34 net30 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net30 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
MMIN1 Ab net55 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 net59 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net55 net47 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 net51 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net47 X VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 X net51 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net55 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 net59 Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net55 net47 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net47 X VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 X net51 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 net51 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlymetal6s4s_1 A VGND VNB VPB VPWR X
MMIN1 Ab X VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 net59 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X net47 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 net51 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net47 net43 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net43 net51 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab X VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 net59 Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 X net47 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net47 net43 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net43 net51 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 net51 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlymetal6s6s_1 A VGND VNB VPB VPWR X
MMIN1 Ab net56 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net56 net48 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 net52 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net48 net44 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net44 net52 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net56 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net56 net48 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net48 net44 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net44 net52 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 net52 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
MMN0 Z net35 sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net39 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net39 TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net35 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB net35 Z VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net39 TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net35 A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
MMN0 Z net35 sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net39 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net39 TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net35 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=2 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB net35 Z VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net39 TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net35 A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ebufn_4 A TE_B VGND VNB VPB VPWR Z
MMN0 Z net35 sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net39 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net39 TE_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net35 A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=4 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB net35 Z VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net39 TE_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net35 A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
MMN0 Z net35 sndA VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net39 VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net39 TE_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net35 A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=8 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB net35 Z VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net39 TE_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net35 A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__edfxbp_1 CLK D DE VGND VNB VPB VPWR Q Q_N
MI14 net124 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net124 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 net68 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net109 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net92 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net92 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net109 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net85 DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 db S1 net85 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 db D net68 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 Q_N S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net193 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net193 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net148 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net168 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net168 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net161 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net161 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 db D net148 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 db S1 net141 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 net141 deneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 Q_N S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__edfxtp_1 CLK D DE VGND VNB VPB VPWR Q
MI14 net115 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net115 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 net59 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net79 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net83 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net83 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net79 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net76 DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 db S1 net76 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 db D net59 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net175 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net175 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net172 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net160 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net160 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net148 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net148 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 db D net172 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 db S1 net128 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 net128 deneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_0 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net25 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net25 TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net25 TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_1 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net25 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net25 TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net25 TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_2 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TE TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=2 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TE TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_4 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TE TE_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=4 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TE TE_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_8 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TE TE_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=8 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TE TE_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvp_1 A TE VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TEB TE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TEB sndTEB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TEB TE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvp_2 A TE VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TEB TE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TEB sndTEB VPB pfet_01v8_hvt m=2 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TEB TE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvp_4 A TE VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TEB TE VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TEB sndTEB VPB pfet_01v8_hvt m=4 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TEB TE VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TEB TE VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TEB sndTEB VPB pfet_01v8_hvt m=8 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TEB TE VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM
MMNs1s nint1 majb sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 COUT majb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj10 majb B sndNAp1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj11 sndNAp1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj30 majb CIN sndNCINn3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj31 sndNCINn3 B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj20 VGND A sndNCINn3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s0 VGND A sndNAn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s1 sndNAn4 B sndNBn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s2 sndNBn4 CIN sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s0 nint1 B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s1 nint1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s2 nint1 CIN VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj10 VPWR A sndPAp1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj11 sndPAp1 B majb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj20 VPWR A sndPCINp3 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj21 sndPCINp3 CIN majb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj31 sndPCINp3 B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s0 VPWR A sndPAp4 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s1 sndPAp4 B sndPBp4 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s2 sndPBp4 CIN sumb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s0 pint1 B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s1 pint1 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s2 pint1 CIN VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1s pint1 majb sumb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fa_2 A B CIN VGND VNB VPB VPWR COUT SUM
MMNs1s nint1 majb sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 COUT majb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj10 majb B sndNAp1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj11 sndNAp1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj30 majb CIN nmajmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj21 nmajmid A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj20 VGND B nmajmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s0 VGND A sndNAn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s1 sndNAn4 B sndNBn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s2 sndNBn4 CIN sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s0 nint1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s1 nint1 B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s2 nint1 CIN VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj10 VPWR A sndPAp1 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj11 sndPAp1 B majb VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj20 VPWR B pmajmid VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj30 pmajmid CIN majb VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj21 pmajmid A VPWR VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s0 VPWR A sndPAp4 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s1 sndPAp4 B sndPBp4 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s2 sndPBp4 CIN sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s0 pint1 A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s1 pint1 B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s2 pint1 CIN VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1s pint1 majb sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fa_4 A B CIN VGND VNB VPB VPWR COUT SUM
MMNs1s nint1 majb sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 COUT majb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj10 majb B sndNAp1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj11 sndNAp1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj30 majb CIN nmajmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj21 nmajmid A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj20 VGND B nmajmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s0 VGND A sndNAn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s1 sndNAn4 B sndNBn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s2 sndNBn4 CIN sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s0 nint1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s1 nint1 B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s2 nint1 CIN VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj10 VPWR A sndPAp1 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj11 sndPAp1 B majb VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj20 VPWR B pmajmid VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj30 pmajmid CIN majb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj21 pmajmid A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s0 VPWR A sndPAp4 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s1 sndPAp4 B sndPBp4 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s2 sndPBp4 CIN sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s0 pint1 A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s1 pint1 B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s2 pint1 CIN VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1s pint1 majb sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fah_1 A B CI VGND VNB VPB VPWR COUT SUM
MMIN2 COUT net195 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM net123 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 CIb mid2 net195 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Bb mid1 net195 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 CIbb mid2 net123 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 CIb mid1 net123 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 CIbb CIb VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 CIb CI VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 Ab2 A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 Abb2 Ab2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI14 Ab1 A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 Abb2 B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 Ab1 Bb mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Abb2 Bb mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Ab1 B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT net195 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM net123 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 CIb mid1 net195 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 Bb mid2 net195 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 CIbb mid1 net123 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 CIb mid2 net123 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 CIbb CIb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 CIb CI VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 Ab2 A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 Abb2 Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 Ab1 A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 Abb2 Bb mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 Ab1 B mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 Abb2 B mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 Ab1 Bb mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fahcin_1 A B CIN VGND VNB VPB VPWR COUT SUM
MMIP3 SUM net144 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 Bbb Bb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 Ab Bb mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 Abb B mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 Abb Bb mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 Ab B mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 CINb1 CIN VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 CINbb2 CINb2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 CINb2 CIN VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 CINbb2 mid2 net144 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 CINb2 mid1 net144 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 Bbb mid2 COUT VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 CINb1 mid1 COUT VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM net144 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 CINb1 mid2 COUT VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Ab B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Abb Bb mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 Ab Bb mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 Abb B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI14 CINb1 CIN VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 CINbb2 CINb2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 CINb2 CIN VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 CINbb2 mid1 net144 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 CINb2 mid2 net144 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 Bbb mid1 COUT VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Bbb Bb VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fahcon_1 A B CI VGND VNB VPB VPWR COUT_N SUM
MMIP3 SUM net146 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 Bb2 B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 Ab Bb1 mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 Abb B mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 Abb Bb1 mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 Ab B mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 CIb1 CI VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 CIbb2 CIb2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 CIb2 CI VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb1 B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 CIb2 mid2 net146 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 CIbb2 mid1 net146 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 Bb2 mid2 COUT_N VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 CIb1 mid1 COUT_N VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM net146 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 CIb1 mid2 COUT_N VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Ab B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Abb Bb1 mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 Ab Bb1 mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 Abb B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI14 CIb1 CI VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 CIbb2 CIb2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 CIb2 CI VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb1 B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 CIb2 mid1 net146 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 CIbb2 mid2 net146 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 Bb2 mid1 COUT_N VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Bb2 B VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__fill_4 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__fill_8 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__ha_1 A B VGND VNB VPB VPWR COUT SUM
MMIN2 COUT majb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A sndNA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B majb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs1 sumb majb nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs20 VGND A nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs21 VGND B nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 majb A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 majb B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1 VPWR majb sumb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs20 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs21 sndPA B sumb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ha_2 A B VGND VNB VPB VPWR COUT SUM
MMIN2 COUT majb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A sndNA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B majb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs1 sumb majb nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs20 VGND A nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs21 VGND B nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 majb A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 majb B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1 VPWR majb sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs20 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs21 sndPA B sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ha_4 A B VGND VNB VPB VPWR COUT SUM
MMIN2 COUT majb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A sndNA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B majb VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs1 sumb majb nint1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs20 VGND A nint1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs21 VGND B nint1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 majb A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 majb B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1 VPWR majb sumb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs20 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs21 sndPA B sumb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Y A VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=12 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=12 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_bleeder_1 SHORT VGND VNB VPB VPWR
MI2 net29 SHORT net25 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net25 SHORT net24 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 VPWR SHORT net29 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 net24 SHORT net16 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net16 SHORT VGND VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_1 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_2 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_4 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_8 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=8 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_16 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_1 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=2 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_2 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_4 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_8 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=8 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=12 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_16 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=24 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_3 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=0.59 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=0.59 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_4 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=1.05 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=1.05 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_6 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=1.97 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=1.97 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_8 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=2.89 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=2.89 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_12 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=4.73 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=4.73 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputiso0n_1 A SLEEP_B VGND VNB VPB VPWR X
MI14 X net36 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 net36 A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 sndA SLEEP_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 net36 SLEEP_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 X net36 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 net36 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputiso0p_1 A SLEEP VGND VNB VPB VPWR X
MI8 net36 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net36 sleepb VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 X net36 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 sleepb SLEEP VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net36 sleepb sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 X net36 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 sleepb SLEEP VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 sndA A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputiso1n_1 A SLEEP_B VGND VNB VPB VPWR X
MI23 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 VPWR net44 X VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 net56 SLEEP_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 sndPA net56 net44 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 net56 SLEEP_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net44 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X net44 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net44 net56 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputiso1p_1 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 sndPA A net36 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 VPWR net36 X VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net36 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net36 SLEEP VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI14 X net36 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputisolatch_1 D SLEEP_B VGND VNB VPB VPWR Q
MI677 Q s0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 sleepneg sleeppos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI674 net39 s0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 s0 sleepneg net49 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net49 D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 sleeppos net38 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net38 net39 VGND VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 sleeppos SLEEP_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 sleeppos SLEEP_B VPWR VPB pfet_01v8_hvt m=1 w=0.55 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 sleepneg sleeppos VPWR VPB pfet_01v8_hvt m=1 w=0.55 l=0.15
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
MI662 net86 net39 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 sleepneg net86 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net39 s0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q s0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 s0 sleeppos net69 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net69 D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_1 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA Ab X VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_2 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA Ab X VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_4 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA Ab X VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_8 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR Ab sndPA VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA SLEEP X VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_16 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR Ab sndPA VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA SLEEP X VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrckapwr_16 A SLEEP KAPWR VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA net58 net66 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net58 A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab net66 KAPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 X Ab KAPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 net66 SLEEP VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 net66 net58 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net58 A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 Ab net66 VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 X Ab VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1 A VGND VPB VPWRIN VPWR X
M1000 X a_1028_32# VPWR VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=2.1725e+11p pd=2.13e+06u as=4.7795e+11p ps=4.37e+06u
M1001 VPWR a_620_911# a_714_58# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
M1002 a_1028_32# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1003 X a_1028_32# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.8525e+11p pd=1.87e+06u as=1.4178e+12p ps=1.319e+07u
M1004 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=0p ps=0u
M1005 a_714_58# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1006 a_714_58# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1007 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1008 a_1028_32# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1009 a_505_297# A VPWRIN VPWRIN pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1010 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1011 VGND A a_714_58# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1012 VGND A a_714_58# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1013 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1014 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_714_58# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2 A VGND VPB VPWRIN VPWR X
M1000 VPWR a_620_911# a_714_47# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=8.352e+11p pd=7.41e+06u as=2.1725e+11p ps=2.13e+06u
M1001 a_1032_911# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.62905e+12p ps=1.514e+07u
M1003 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1004 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1005 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=2.405e+11p pd=2.04e+06u as=0p ps=0u
M1006 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=3.7e+11p ps=2.74e+06u
M1007 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1008 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1009 a_1032_911# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1010 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1011 a_505_297# A VPWRIN VPWRIN pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1012 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1013 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1014 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1015 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1016 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_714_47# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4 A VGND VPB VPWRIN VPWR X
M1000 VPWR a_620_911# a_714_47# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=1.1152e+12p pd=9.97e+06u as=2.1725e+11p ps=2.13e+06u
M1001 a_1032_911# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u
+ ad=6.5e+11p pd=5.3e+06u as=0p ps=0u
M1003 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.81105e+12p ps=1.7e+07u
M1004 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1005 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1006 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=4.225e+11p pd=3.9e+06u as=0p ps=0u
M1007 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1008 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1009 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1010 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1011 a_1032_911# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1012 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1013 a_505_297# A VPWRIN VPWRIN pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1014 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1015 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1016 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1017 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1018 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1019 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1020 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_714_47# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4 A LOWLVPWR VGND VNB VPB VPWR X
MI2 net72 cross1 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 cross1 net72 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 Ab A LOWLVPWR LOWLVPWR pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 X net60 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 net60 cross1 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 cross1 Ab VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 net72 A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 X net60 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 net60 cross1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1 A LOWLVPWR VGND VPB VPWR X
M1000 X a_1028_32# VPWR VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=2.1725e+11p pd=2.13e+06u as=4.7795e+11p ps=4.37e+06u
M1001 VPWR a_620_911# a_714_58# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
M1002 a_1028_32# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1003 X a_1028_32# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.8525e+11p pd=1.87e+06u as=1.4178e+12p ps=1.319e+07u
M1004 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=0p ps=0u
M1005 a_714_58# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1006 a_714_58# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1007 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1008 a_1028_32# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1009 a_505_297# A LOWLVPWR LOWLVPWR pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1010 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1011 VGND A a_714_58# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1012 VGND A a_714_58# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1013 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1014 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_714_58# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2 A LOWLVPWR VGND VPB VPWR X
M1000 VPWR a_620_911# a_714_47# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=8.352e+11p pd=7.41e+06u as=2.1725e+11p ps=2.13e+06u
M1001 a_1032_911# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.62905e+12p ps=1.514e+07u
M1003 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1004 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1005 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=2.405e+11p pd=2.04e+06u as=0p ps=0u
M1006 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=3.7e+11p ps=2.74e+06u
M1007 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1008 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1009 a_1032_911# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1010 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1011 a_505_297# A LOWLVPWR LOWLVPWR pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1012 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1013 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1014 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1015 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1016 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_714_47# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4 A LOWLVPWR VGND VPB VPWR X
M1000 VPWR a_620_911# a_714_47# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=1.1152e+12p pd=9.97e+06u as=2.1725e+11p ps=2.13e+06u
M1001 a_1032_911# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u
+ ad=6.5e+11p pd=5.3e+06u as=0p ps=0u
M1003 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.81105e+12p ps=1.7e+07u
M1004 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1005 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1006 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=4.225e+11p pd=3.9e+06u as=0p ps=0u
M1007 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1008 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1009 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1010 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1011 a_1032_911# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1012 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1013 a_505_297# A LOWLVPWR LOWLVPWR pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1014 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1015 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1016 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1017 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1018 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1019 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1020 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_714_47# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__macro_sparecell VGND VNB VPB VPWR LO
XI1 VGND VNB VPB VPWR net59 LO / sky130_fd_sc_hd__conb_1
XI2 LO LO VGND VNB VPB VPWR nd2right / sky130_fd_sc_hd__nand2_2
XI3 LO LO VGND VNB VPB VPWR nd2left / sky130_fd_sc_hd__nand2_2
XI4 nd2right nd2right VGND VNB VPB VPWR nor2right / sky130_fd_sc_hd__nor2_2
XI5 nd2left nd2left VGND VNB VPB VPWR nor2left / sky130_fd_sc_hd__nor2_2
XI6 nor2right VGND VNB VPB VPWR invright / sky130_fd_sc_hd__inv_2
XI7 nor2left VGND VNB VPB VPWR invleft / sky130_fd_sc_hd__inv_2
.ENDS




.SUBCKT sky130_fd_sc_hd__maj3_1 A B C VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN10 y B sndNBa VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN11 sndNBa A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN20 y B sndNBc VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN21 sndNBc C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN30 y C sndNCa VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN31 sndNCa A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP10 VPWR A sndPAb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP11 sndPAb B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP20 VPWR C sndPCb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP21 sndPCb B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP30 VPWR A sndPAc VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP31 sndPAc C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__maj3_2 A B C VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN10 y B sndNBa VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN11 sndNBa A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN20 y B sndNBc VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN21 sndNBc C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN30 y C sndNCa VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN31 sndNCa A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP10 VPWR A sndPAb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP11 sndPAb B y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP20 VPWR C sndPCb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP21 sndPCb B y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP30 VPWR A sndPAc VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP31 sndPAc C y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__maj3_4 A B C VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN10 y B sndNBa VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN11 sndNBa A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN20 y B sndNBc VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN21 sndNBc C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN30 y C sndNCa VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN31 sndNCa A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP10 VPWR A sndPAb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP11 sndPAb B y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP20 VPWR C sndPCb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP21 sndPCb B y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP30 VPWR A sndPAc VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP31 sndPAc C y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
MMNA00 xb A0 smdNA0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 xb A1 sndNA1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X xb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 xb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 xb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X xb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
MMNA00 xb A0 smdNA0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 xb A1 sndNA1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X xb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 xb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 xb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X xb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
MMNA00 xb A0 smdNA0 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 xb A1 sndNA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X xb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 xb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 xb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X xb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
MMNA00 xb A0 smdNA0 VNB nfet_01v8 m=2 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=2 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 xb A1 sndNA1 VNB nfet_01v8 m=2 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=2 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X xb VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 xb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 xb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X xb VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2i_1 A0 A1 S VGND VNB VPB VPWR Y
MMNA00 Y A0 smdNA0 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 Y A1 sndNA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2i_2 A0 A1 S VGND VNB VPB VPWR Y
MMNA00 Y A0 smdNA0 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 Y A1 sndNA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2i_4 A0 A1 S VGND VNB VPB VPWR Y
MMNA00 Y A0 smdNA0 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 Y A1 sndNA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
MMNA00 sndNS0ba0 S0b xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA01 VGND A0 sndNS0ba0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA10 sndNS0a1 S0 xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA11 VGND A1 sndNS0a1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA20 sndNS0ba2 S0b xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA21 VGND A2 sndNS0ba2 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA30 sndNS0a3 S0 xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA31 VGND A3 sndNS0a3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs1o xb S1b xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs2o xb S1 xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN1 VGND S1 S1b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN2 VGND S0 S0b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN4 VGND xb X VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA00 sndPA0a0 A0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA01 xlowb S0 sndPA0a0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA10 sndPA1a1 A1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA11 xlowb S0b sndPA1a1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA20 sndPA2a2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA21 xhib S0 sndPA2a2 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA30 sndPA3a3 A3 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA31 xhib S0b sndPA3a3 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs1o xb S1 xlowb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs2o xb S1b xhib VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP1 VPWR S1 S1b VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP2 VPWR S0 S0b VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP4 VPWR xb X VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
MMNA00 sndNS0ba0 S0b xlowb VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA01 VGND A0 sndNS0ba0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA10 sndNS0a1 S0 xlowb VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA11 VGND A1 sndNS0a1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA20 sndNS0ba2 S0b xhib VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA21 VGND A2 sndNS0ba2 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA30 sndNS0a3 S0 xhib VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA31 VGND A3 sndNS0a3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs1o xb S1b xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs2o xb S1 xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN1 VGND S1 S1b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN2 VGND S0 S0b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN4 VGND xb X VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA00 sndPA0a0 A0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA01 xlowb S0 sndPA0a0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA10 sndPA1a1 A1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA11 xlowb S0b sndPA1a1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA20 sndPA2a2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA21 xhib S0 sndPA2a2 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA30 sndPA3a3 A3 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA31 xhib S0b sndPA3a3 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs1o xb S1 xlowb VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs2o xb S1b xhib VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP1 VPWR S1 S1b VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP2 VPWR S0 S0b VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP4 VPWR xb X VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__mux4_4 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
MMNA00 sndNS0ba0 S0b xlowb VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA01 VGND A0 sndNS0ba0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA10 sndNS0a1 S0 xlowb VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA11 VGND A1 sndNS0a1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA20 sndNS0ba2 S0b xhib VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA21 VGND A2 sndNS0ba2 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA30 sndNS0a3 S0 xhib VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA31 VGND A3 sndNS0a3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs1o xb S1b xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs2o xb S1 xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN1 VGND S1 S1b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN2 VGND S0 S0b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN4 VGND xb X VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA00 sndPA0a0 A0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA01 xlowb S0 sndPA0a0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA10 sndPA1a1 A1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA11 xlowb S0b sndPA1a1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA20 sndPA2a2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA21 xhib S0 sndPA2a2 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA30 sndPA3a3 A3 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA31 xhib S0b sndPA3a3 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs1o xb S1 xlowb VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs2o xb S1b xhib VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP1 VPWR S1 S1b VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP2 VPWR S0 S0b VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP4 VPWR xb X VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP3 sndPC D Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN3 Y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP3 sndPC D Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN3 Y D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP3 sndPC D Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN3 Y D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4bb_1 A B C_N D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4bb_2 A B C_N D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4bb_4 A B C_N D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inand nmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inand VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inand nmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inand VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inand nmid VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inand VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA20 VPWR A1 snd2A1 VPB pfet_01v8_hvt w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA21 snd2A1 A2 y VPB pfet_01v8_hvt w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ai_0 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=0.7 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311ai_0 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 pndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 pndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 pndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 pndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 pndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 pndC VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2_0 A B VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__probe_p_8 A VGND VNB VPB VPWR X
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 net29 Ab VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 net29 Ab VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
rI112 net29 X sky130_fd_pr__res_generic_m5
.ENDS




.SUBCKT sky130_fd_sc_hd__probec_p_8 A VGND VNB VPB VPWR X
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 net33 Ab VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 net33 Ab VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
rI112 net33 X short
rI120 VGND met5vgnd short
rI119 VPWR met5vpwr short
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfbbn_1 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI98 net105 D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 net105 SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net176 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net213 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net153 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net153 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net145 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net145 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net117 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net213 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net105 clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net125 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net125 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net117 RESET net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net117 S0 net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net116 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 net105 D p0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 net105 sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net265 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net213 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net117 S0 net268 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net265 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net216 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net257 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net257 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net117 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net268 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net241 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net105 clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net241 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net216 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net213 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net117 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfbbn_2 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI98 net105 D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 net105 SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net176 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net213 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net160 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net160 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net145 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net145 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net117 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net213 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net105 clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net128 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net128 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net117 RESET net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net117 S0 net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net116 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 net105 D p0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 net105 sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net265 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net213 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net117 S0 net268 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net265 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net216 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net257 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net257 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net117 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net268 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net241 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net105 clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net241 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net216 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net213 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net117 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfbbp_1 CLK D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI98 net105 D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 net105 SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net176 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net213 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net160 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net160 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net145 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net145 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net117 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net213 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net105 clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net125 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net125 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net117 RESET net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net117 S0 net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net116 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 net105 D p0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 net105 sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net265 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net213 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net117 S0 net268 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net265 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net216 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net257 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net257 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net117 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net268 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net241 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net105 clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net241 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net216 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net213 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net117 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrbp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net92 S0 net134 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net134 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net127 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net115 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net115 M1 net127 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net103 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net92 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net103 net92 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI672 net171 net92 VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 Q_N net171 VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net215 net92 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net92 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net215 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net92 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net194 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net92 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI673 net171 net92 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI671 Q_N net171 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrbp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net92 S0 net134 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net134 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net127 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net115 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net115 M1 net127 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net110 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net92 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 net92 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI672 net171 net92 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 Q_N net171 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net215 net92 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net92 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net215 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net92 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net194 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net92 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI673 net171 net92 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI671 Q_N net171 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrtn_1 CLK_N D RESET_B SCD SCE VGND VNB VPB VPWR Q
MI642 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net87 net153 net117 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net117 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net110 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net98 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net98 M1 net110 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 net153 clkneg net93 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net87 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net93 net87 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos net153 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net190 net87 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net87 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 net153 clkpos net190 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net87 net153 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net169 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net169 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net169 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net87 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg net153 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net84 S0 net114 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net114 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net107 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net95 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net95 M1 net107 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net83 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net84 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net83 net84 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net187 net84 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net84 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net187 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net84 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net166 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net166 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net166 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net84 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net84 S0 net114 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net114 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net107 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net95 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net95 M1 net107 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net90 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net84 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net90 net84 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net187 net84 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net84 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net187 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net84 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net166 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net166 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net166 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net84 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrtp_4 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net84 S0 net114 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net114 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net107 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net95 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net95 M1 net107 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net90 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net84 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net90 net84 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net187 net84 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net84 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net187 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net84 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net166 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net166 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net166 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net84 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfsbp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net159 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net159 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net138 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net138 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net199 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net199 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net98 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net98 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI27 net243 S1 net215 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net230 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net227 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net199 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net215 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net206 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net199 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net227 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net206 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net230 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net243 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfsbp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net195 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net195 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net130 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net130 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net107 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net107 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N S0 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI34 S0 clkpos net219 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net239 S1 net187 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net230 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net199 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net230 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net219 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net239 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net199 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net195 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net187 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net195 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N S0 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfstp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net165 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net165 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net109 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net109 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net96 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net96 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net84 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net84 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net189 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net209 S1 net157 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net200 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net169 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net189 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net209 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net169 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net165 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net157 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net165 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfstp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net165 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net165 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net109 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net109 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net96 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net96 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net84 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net84 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net212 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net209 S1 net157 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net200 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net196 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net212 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net209 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net196 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net165 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net157 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net165 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfstp_4 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net165 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net165 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net104 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net104 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net96 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net96 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net84 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net84 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net189 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net209 S1 net157 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net200 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net169 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net189 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net209 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net169 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net165 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net157 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net165 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxbp_1 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI657 M0 clkpos net129 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net129 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net120 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net120 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net153 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net153 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net177 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net160 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q_N net153 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net177 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net160 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 net153 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxbp_2 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI657 M0 clkpos net129 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net129 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net120 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net120 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net153 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net153 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net196 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net189 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q_N net153 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net196 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net189 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 net153 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxtp_1 CLK D SCD SCE VGND VNB VPB VPWR Q
MI652 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net78 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net78 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net54 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net54 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net155 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxtp_2 CLK D SCD SCE VGND VNB VPB VPWR Q
MI652 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net78 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net78 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net54 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net54 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 net163 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net138 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net138 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net163 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxtp_4 CLK D SCD SCE VGND VNB VPB VPWR Q
MI652 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net78 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net78 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net54 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net54 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 net163 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net155 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net163 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdlclkp_1 CLK GATE SCE VGND VNB VPB VPWR GCLK
MI662 net88 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net88 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net76 CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net76 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 net63 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 net116 GATE net63 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net76 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net116 clkneg M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net116 clkpos M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net123 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net123 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 net116 SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net112 CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net76 m1 net112 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 net116 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net76 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdlclkp_2 CLK GATE SCE VGND VNB VPB VPWR GCLK
MI662 net88 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net88 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net76 CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net76 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 net63 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 net116 GATE net63 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net76 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net116 clkneg M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net116 clkpos M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net123 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net123 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 net116 SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net112 CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net76 m1 net112 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 net116 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net76 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdlclkp_4 CLK GATE SCE VGND VNB VPB VPWR GCLK
MI662 net88 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net88 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net76 CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net76 m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 net63 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 net116 GATE net63 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net76 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net116 clkneg M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net116 clkpos M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net123 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net123 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 net116 SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net112 CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net76 m1 net112 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 net116 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net76 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxbp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
MI14 net155 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net123 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net127 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net127 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net123 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net116 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net107 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net107 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net104 D net116 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net104 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net104 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI52 Q_N q1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net235 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net235 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net224 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net224 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net104 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net104 D net203 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net200 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net192 q1 net104 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net192 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net203 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net176 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net176 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI53 Q_N q1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxbp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
MI14 net155 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net144 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net127 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net127 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net144 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net116 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net107 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net107 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net104 D net116 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net104 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net104 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI52 Q_N q1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net240 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net240 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net224 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net224 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net104 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net104 D net180 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net200 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net192 q1 net104 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net192 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net180 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net176 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net176 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI53 Q_N q1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxtp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q
MI14 net146 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net146 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net114 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net118 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net118 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net114 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net94 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net103 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net103 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net95 D net94 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net95 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net95 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net222 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net222 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net211 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net211 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net95 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net95 D net167 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net187 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net187 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net179 q1 net95 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net179 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net167 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net158 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net158 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxtp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q
MI14 net146 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net146 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net114 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net118 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net118 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net114 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net94 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net98 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net98 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net95 D net94 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net95 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net95 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net222 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net222 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net211 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net211 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net95 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net95 D net167 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net187 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net187 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net174 q1 net95 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net174 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net167 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net158 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net158 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxtp_4 CLK D DE SCD SCE VGND VNB VPB VPWR Q
MI14 net146 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net146 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net135 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net118 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net118 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net135 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net107 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net98 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net98 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net95 D net107 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net95 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net95 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net227 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net227 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net206 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net206 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net95 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net95 D net190 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net187 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net187 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net174 q1 net95 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net174 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net190 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net163 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net163 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__tap_1 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__tap_2 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__tapvgnd2_1 VGND VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__tapvgnd_1 VGND VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
MMNnand0 VGND A sndNA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B inand VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPA B Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
MMNnand0 VGND A sndNA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B inand VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPA B Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
MMNnand0 VGND A sndNA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B inand VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPA B Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor3_1 A B C VGND VNB VPB VPWR X
MMIN3 X net57 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 Cb net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 C net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X net57 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 C net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 mid2 Cb net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor3_2 A B C VGND VNB VPB VPWR X
MMIN3 X net57 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 Cb net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 C net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X net57 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 C net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 mid2 Cb net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor3_4 A B C VGND VNB VPB VPWR X
MMIN3 X net57 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 Cb net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 C net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X net57 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 C net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 mid2 Cb net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
MMNnor0 inor A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND A sndNA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNA B X VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 X inor VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA B inor VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 X inor pmid VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
MMNnor0 inor A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND A sndNA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNA B X VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 X inor VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA B inor VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 X inor pmid VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
MMNnor0 inor A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND A sndNA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNA B X VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 X inor VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA B inor VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 X inor pmid VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor3_1 A B C VGND VNB VPB VPWR X
MMIP3 X net117 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 Cb net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 mid2 C net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X net117 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 C net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 Cb net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor3_2 A B C VGND VNB VPB VPWR X
MMIP3 X net117 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 Cb net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 mid2 C net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X net117 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 C net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 Cb net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor3_4 A B C VGND VNB VPB VPWR X
MMIP3 X net117 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 Cb net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 mid2 C net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X net117 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 C net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 Cb net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS














































.subckt riscv_pipeline_top M_AXI_ARADDR[10] M_AXI_ARADDR[11] M_AXI_ARADDR[12] M_AXI_ARADDR[22]
+ M_AXI_ARADDR[23] M_AXI_ARADDR[24] M_AXI_ARADDR[25] M_AXI_ARADDR[28] M_AXI_ARADDR[29]
+ M_AXI_ARADDR[3] M_AXI_ARADDR[4] M_AXI_ARADDR[5] M_AXI_ARADDR[9] M_AXI_ARREADY M_AXI_ARVALID
+ M_AXI_AWADDR[1] M_AXI_AWADDR[20] M_AXI_AWADDR[21] M_AXI_AWADDR[22] M_AXI_AWADDR[23]
+ M_AXI_AWADDR[24] M_AXI_AWADDR[25] M_AXI_AWADDR[26] M_AXI_AWADDR[27] M_AXI_AWADDR[28]
+ M_AXI_AWADDR[29] M_AXI_AWADDR[2] M_AXI_AWADDR[7] M_AXI_AWADDR[8] M_AXI_AWADDR[9]
+ M_AXI_AWREADY M_AXI_BREADY M_AXI_BRESP[0] M_AXI_BRESP[1] M_AXI_BVALID M_AXI_RDATA[0]
+ M_AXI_RDATA[10] M_AXI_RDATA[11] M_AXI_RDATA[12] M_AXI_RDATA[13] M_AXI_RDATA[14]
+ M_AXI_RDATA[15] M_AXI_RDATA[16] M_AXI_RDATA[17] M_AXI_RDATA[18] M_AXI_RDATA[19]
+ M_AXI_RDATA[1] M_AXI_RDATA[20] M_AXI_RDATA[21] M_AXI_RDATA[22] M_AXI_RDATA[23] M_AXI_RDATA[24]
+ M_AXI_RDATA[25] M_AXI_RDATA[26] M_AXI_RDATA[27] M_AXI_RDATA[28] M_AXI_RDATA[29]
+ M_AXI_RDATA[2] M_AXI_RDATA[30] M_AXI_RDATA[31] M_AXI_RDATA[3] M_AXI_RDATA[4] M_AXI_RDATA[5]
+ M_AXI_RDATA[6] M_AXI_RDATA[7] M_AXI_RDATA[8] M_AXI_RDATA[9] M_AXI_RREADY M_AXI_RRESP[0]
+ M_AXI_RRESP[1] M_AXI_RVALID M_AXI_WDATA[0] M_AXI_WDATA[15] M_AXI_WDATA[16] M_AXI_WDATA[17]
+ M_AXI_WDATA[18] M_AXI_WDATA[19] M_AXI_WDATA[1] M_AXI_WDATA[22] M_AXI_WDATA[23] M_AXI_WDATA[24]
+ M_AXI_WDATA[25] M_AXI_WDATA[26] M_AXI_WDATA[27] M_AXI_WDATA[2] M_AXI_WDATA[30] M_AXI_WDATA[31]
+ M_AXI_WDATA[3] M_AXI_WDATA[4] M_AXI_WDATA[5] M_AXI_WREADY M_AXI_WSTRB[0] M_AXI_WSTRB[1]
+ M_AXI_WSTRB[2] M_AXI_WSTRB[3] M_AXI_WVALID VGND VPWR clk led[0] led[1] led[2] led[3]
+ led[5] led[6] led[7] led[8] led[9] rst_n M_AXI_WDATA[21] M_AXI_WDATA[20] M_AXI_ARADDR[15]
+ M_AXI_ARADDR[14] M_AXI_ARADDR[13] M_AXI_ARADDR[2] M_AXI_ARADDR[1] M_AXI_AWADDR[12]
+ M_AXI_AWADDR[11] M_AXI_AWADDR[0] M_AXI_ARADDR[0] M_AXI_AWVALID M_AXI_AWADDR[10]
+ M_AXI_ARADDR[21] M_AXI_ARADDR[20] M_AXI_ARADDR[31] M_AXI_WDATA[9] M_AXI_AWADDR[31]
+ M_AXI_ARADDR[8] M_AXI_WDATA[8] M_AXI_AWADDR[19] M_AXI_ARADDR[30] M_AXI_ARADDR[19]
+ M_AXI_AWADDR[30] M_AXI_ARADDR[7] M_AXI_ARADDR[18] M_AXI_WDATA[7] M_AXI_AWADDR[18]
+ M_AXI_WDATA[6] M_AXI_AWADDR[6] M_AXI_ARADDR[6] M_AXI_AWADDR[17] M_AXI_ARADDR[17]
+ M_AXI_AWADDR[5] M_AXI_AWADDR[16] M_AXI_ARADDR[27] M_AXI_ARADDR[16] M_AXI_AWADDR[4]
+ M_AXI_ARADDR[26] M_AXI_AWADDR[15] M_AXI_AWADDR[3] M_AXI_WDATA[14] M_AXI_AWADDR[14]
+ M_AXI_AWADDR[13] M_AXI_WDATA[13] M_AXI_WDATA[12] M_AXI_WDATA[11] M_AXI_WDATA[10]
+ M_AXI_WDATA[29] M_AXI_WDATA[28] led[4]
XFILLER_0_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_61 VGND VGND VPWR VPWR riscv_pipeline_top_61/HI M_AXI_AWADDR[14]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_139_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_72 VGND VGND VPWR VPWR riscv_pipeline_top_72/HI M_AXI_AWADDR[25]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_50 VGND VGND VPWR VPWR riscv_pipeline_top_50/HI M_AXI_AWADDR[3]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_83 VGND VGND VPWR VPWR riscv_pipeline_top_83/HI M_AXI_WDATA[3]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_94 VGND VGND VPWR VPWR riscv_pipeline_top_94/HI M_AXI_WDATA[14]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_155_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_200_ clknet_1_1__leaf_clk _011_ net11 VGND VGND VPWR VPWR counter\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_131_ _044_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_109 VGND VGND VPWR VPWR riscv_pipeline_top_109/HI M_AXI_WDATA[29]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_173_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_114_ _091_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput7 net7 VGND VGND VPWR VPWR M_AXI_BREADY sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_73 VGND VGND VPWR VPWR riscv_pipeline_top_73/HI M_AXI_AWADDR[26]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_102_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xriscv_pipeline_top_40 VGND VGND VPWR VPWR riscv_pipeline_top_40/HI M_AXI_ARADDR[26]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_62 VGND VGND VPWR VPWR riscv_pipeline_top_62/HI M_AXI_AWADDR[15]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_51 VGND VGND VPWR VPWR riscv_pipeline_top_51/HI M_AXI_AWADDR[4]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_31_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_84 VGND VGND VPWR VPWR riscv_pipeline_top_84/HI M_AXI_WDATA[4]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_95 VGND VGND VPWR VPWR riscv_pipeline_top_95/HI M_AXI_WDATA[15]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_155_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_130_ _042_ _043_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__and2b_1
XFILLER_0_93_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_113_ _089_ _090_ VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__and2b_1
XFILLER_0_62_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput8 net8 VGND VGND VPWR VPWR M_AXI_RREADY sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_30 VGND VGND VPWR VPWR riscv_pipeline_top_30/HI M_AXI_ARADDR[16]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_20_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xriscv_pipeline_top_41 VGND VGND VPWR VPWR riscv_pipeline_top_41/HI M_AXI_ARADDR[27]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_52 VGND VGND VPWR VPWR riscv_pipeline_top_52/HI M_AXI_AWADDR[5]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_63 VGND VGND VPWR VPWR riscv_pipeline_top_63/HI M_AXI_AWADDR[16]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_31_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_74 VGND VGND VPWR VPWR riscv_pipeline_top_74/HI M_AXI_AWADDR[27]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_85 VGND VGND VPWR VPWR riscv_pipeline_top_85/HI M_AXI_WDATA[5]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_102_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_96 VGND VGND VPWR VPWR riscv_pipeline_top_96/HI M_AXI_WDATA[16]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_917 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_189_ clknet_1_0__leaf_clk _025_ net10 VGND VGND VPWR VPWR counter\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_112_ counter\[1\] counter\[0\] counter\[2\] counter\[3\] VGND VGND VPWR VPWR _090_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_123_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold10 counter\[15\] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput9 net9 VGND VGND VPWR VPWR M_AXI_WVALID sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xriscv_pipeline_top_20 VGND VGND VPWR VPWR riscv_pipeline_top_20/HI M_AXI_ARADDR[6]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_31_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_31 VGND VGND VPWR VPWR riscv_pipeline_top_31/HI M_AXI_ARADDR[17]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_42 VGND VGND VPWR VPWR riscv_pipeline_top_42/HI M_AXI_ARADDR[28]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_130_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_53 VGND VGND VPWR VPWR riscv_pipeline_top_53/HI M_AXI_AWADDR[6]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_64 VGND VGND VPWR VPWR riscv_pipeline_top_64/HI M_AXI_AWADDR[17]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_43_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xriscv_pipeline_top_86 VGND VGND VPWR VPWR riscv_pipeline_top_86/HI M_AXI_WDATA[6]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_75 VGND VGND VPWR VPWR riscv_pipeline_top_75/HI M_AXI_AWADDR[28]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_20_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xriscv_pipeline_top_97 VGND VGND VPWR VPWR riscv_pipeline_top_97/HI M_AXI_WDATA[17]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_101_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_188_ clknet_1_1__leaf_clk _024_ net11 VGND VGND VPWR VPWR counter\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_111_ _088_ VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__buf_2
XFILLER_0_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold11 counter\[2\] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xriscv_pipeline_top_21 VGND VGND VPWR VPWR riscv_pipeline_top_21/HI M_AXI_ARADDR[7]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_20_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_54 VGND VGND VPWR VPWR riscv_pipeline_top_54/HI M_AXI_AWADDR[7]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_43 VGND VGND VPWR VPWR riscv_pipeline_top_43/HI M_AXI_ARADDR[29]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_32 VGND VGND VPWR VPWR riscv_pipeline_top_32/HI M_AXI_ARADDR[18]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xriscv_pipeline_top_65 VGND VGND VPWR VPWR riscv_pipeline_top_65/HI M_AXI_AWADDR[18]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_130_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xriscv_pipeline_top_76 VGND VGND VPWR VPWR riscv_pipeline_top_76/HI M_AXI_AWADDR[29]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_87 VGND VGND VPWR VPWR riscv_pipeline_top_87/HI M_AXI_WDATA[7]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_98 VGND VGND VPWR VPWR riscv_pipeline_top_98/HI M_AXI_WDATA[18]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_187_ clknet_1_1__leaf_clk _017_ net11 VGND VGND VPWR VPWR counter\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_110_ counter\[1\] counter\[0\] counter\[2\] counter\[3\] VGND VGND VPWR VPWR _088_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold12 counter\[8\] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_959 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_33 VGND VGND VPWR VPWR riscv_pipeline_top_33/HI M_AXI_ARADDR[19]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_55 VGND VGND VPWR VPWR riscv_pipeline_top_55/HI M_AXI_AWADDR[8]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_130_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_44 VGND VGND VPWR VPWR riscv_pipeline_top_44/HI M_AXI_ARADDR[30]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_20_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_22 VGND VGND VPWR VPWR riscv_pipeline_top_22/HI M_AXI_ARADDR[8]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_77 VGND VGND VPWR VPWR riscv_pipeline_top_77/HI M_AXI_AWADDR[30]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_66 VGND VGND VPWR VPWR riscv_pipeline_top_66/HI M_AXI_AWADDR[19]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_88 VGND VGND VPWR VPWR riscv_pipeline_top_88/HI M_AXI_WDATA[8]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_99 VGND VGND VPWR VPWR riscv_pipeline_top_99/HI M_AXI_WDATA[19]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_99_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_970 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_186_ clknet_1_1__leaf_clk _006_ net10 VGND VGND VPWR VPWR counter\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_169_ _067_ _068_ VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__and2b_1
XFILLER_0_97_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold13 counter\[13\] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xriscv_pipeline_top_23 VGND VGND VPWR VPWR riscv_pipeline_top_23/HI M_AXI_ARADDR[9]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_34 VGND VGND VPWR VPWR riscv_pipeline_top_34/HI M_AXI_ARADDR[20]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_45 VGND VGND VPWR VPWR riscv_pipeline_top_45/HI M_AXI_ARADDR[31]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_20_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_78 VGND VGND VPWR VPWR riscv_pipeline_top_78/HI M_AXI_AWADDR[31]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_56 VGND VGND VPWR VPWR riscv_pipeline_top_56/HI M_AXI_AWADDR[9]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_67 VGND VGND VPWR VPWR riscv_pipeline_top_67/HI M_AXI_AWADDR[20]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_89 VGND VGND VPWR VPWR riscv_pipeline_top_89/HI M_AXI_WDATA[9]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_99_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_982 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_185_ net2 AXI_BRIDGE.state\[3\] _077_ _078_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__a31o_1
XFILLER_0_52_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_168_ counter\[22\] _054_ _059_ _062_ counter\[23\] VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__a41o_1
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_099_ AXI_BRIDGE.state\[1\] net1 _081_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold14 counter\[4\] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xriscv_pipeline_top_24 VGND VGND VPWR VPWR riscv_pipeline_top_24/HI M_AXI_ARADDR[10]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_35 VGND VGND VPWR VPWR riscv_pipeline_top_35/HI M_AXI_ARADDR[21]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_46 VGND VGND VPWR VPWR riscv_pipeline_top_46/HI M_AXI_ARVALID
+ sky130_fd_sc_hd__conb_1
XFILLER_0_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xriscv_pipeline_top_57 VGND VGND VPWR VPWR riscv_pipeline_top_57/HI M_AXI_AWADDR[10]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_68 VGND VGND VPWR VPWR riscv_pipeline_top_68/HI M_AXI_AWADDR[21]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_79 VGND VGND VPWR VPWR riscv_pipeline_top_79/HI M_AXI_AWVALID
+ sky130_fd_sc_hd__conb_1
XFILLER_0_98_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_184_ _079_ _001_ _075_ net9 VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__o31a_1
XFILLER_0_91_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_167_ _053_ _059_ _066_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_098_ net4 AXI_BRIDGE.state\[4\] VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold15 counter\[12\] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_219_ AXI_BRIDGE.clk _033_ net12 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_107_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xriscv_pipeline_top_14 VGND VGND VPWR VPWR riscv_pipeline_top_14/HI M_AXI_ARADDR[0]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_36 VGND VGND VPWR VPWR riscv_pipeline_top_36/HI M_AXI_ARADDR[22]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_25 VGND VGND VPWR VPWR riscv_pipeline_top_25/HI M_AXI_ARADDR[11]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_43_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xriscv_pipeline_top_69 VGND VGND VPWR VPWR riscv_pipeline_top_69/HI M_AXI_AWADDR[22]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_47 VGND VGND VPWR VPWR riscv_pipeline_top_47/HI M_AXI_AWADDR[0]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_58 VGND VGND VPWR VPWR riscv_pipeline_top_58/HI M_AXI_AWADDR[11]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_183_ _079_ VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_166_ counter\[22\] counter\[23\] _062_ VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_097_ _080_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold16 counter\[16\] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_218_ AXI_BRIDGE.clk _032_ net13 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_53_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_149_ counter\[16\] counter\[17\] _054_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__nand3_1
XFILLER_0_13_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_37 VGND VGND VPWR VPWR riscv_pipeline_top_37/HI M_AXI_ARADDR[23]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_26 VGND VGND VPWR VPWR riscv_pipeline_top_26/HI M_AXI_ARADDR[12]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_102_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xriscv_pipeline_top_15 VGND VGND VPWR VPWR riscv_pipeline_top_15/HI M_AXI_ARADDR[1]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_4_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_48 VGND VGND VPWR VPWR riscv_pipeline_top_48/HI M_AXI_AWADDR[1]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_59 VGND VGND VPWR VPWR riscv_pipeline_top_59/HI M_AXI_AWADDR[12]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_153_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_182_ AXI_BRIDGE.state\[2\] net5 _074_ _076_ net7 VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__a32o_1
XFILLER_0_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_165_ net129 _063_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__xor2_1
XFILLER_0_80_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_096_ net1 AXI_BRIDGE.state\[1\] VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__and2b_1
XFILLER_0_21_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold17 AXI_BRIDGE.clk VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_217_ AXI_BRIDGE.clk _005_ net12 VGND VGND VPWR VPWR AXI_BRIDGE.state\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_148_ net141 _054_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__xor2_1
XFILLER_0_52_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_16 VGND VGND VPWR VPWR riscv_pipeline_top_16/HI M_AXI_ARADDR[2]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_142_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_27 VGND VGND VPWR VPWR riscv_pipeline_top_27/HI M_AXI_ARADDR[13]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_32_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_38 VGND VGND VPWR VPWR riscv_pipeline_top_38/HI M_AXI_ARADDR[24]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_102_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xriscv_pipeline_top_49 VGND VGND VPWR VPWR riscv_pipeline_top_49/HI M_AXI_AWADDR[2]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_181_ _082_ _075_ _083_ _079_ VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__a211o_1
XFILLER_0_80_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_164_ _065_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_095_ net2 AXI_BRIDGE.state\[3\] _079_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_216_ AXI_BRIDGE.clk _004_ net13 VGND VGND VPWR VPWR AXI_BRIDGE.state\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_147_ net135 _051_ _054_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_52_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_17 VGND VGND VPWR VPWR riscv_pipeline_top_17/HI M_AXI_ARADDR[3]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_13_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xriscv_pipeline_top_39 VGND VGND VPWR VPWR riscv_pipeline_top_39/HI M_AXI_ARADDR[25]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_28 VGND VGND VPWR VPWR riscv_pipeline_top_28/HI M_AXI_ARADDR[14]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_141_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout10 net6 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_180_ AXI_BRIDGE.state\[0\] AXI_BRIDGE.state\[2\] VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_163_ _063_ _064_ VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__and2b_1
XFILLER_0_80_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_094_ net5 AXI_BRIDGE.state\[2\] VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__and2b_1
XFILLER_0_33_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_215_ AXI_BRIDGE.clk _001_ net12 VGND VGND VPWR VPWR AXI_BRIDGE.state\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_146_ _053_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__buf_2
XFILLER_0_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_129_ counter\[8\] _089_ _038_ counter\[9\] VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xriscv_pipeline_top_18 VGND VGND VPWR VPWR riscv_pipeline_top_18/HI M_AXI_ARADDR[4]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_82_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_29 VGND VGND VPWR VPWR riscv_pipeline_top_29/HI M_AXI_ARADDR[15]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_149_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout11 net6 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_162_ counter\[20\] _054_ _059_ counter\[21\] VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_093_ net3 AXI_BRIDGE.state\[5\] net4 AXI_BRIDGE.state\[4\] AXI_BRIDGE.state\[0\]
+ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__a221o_1
XFILLER_0_150_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 M_AXI_ARREADY VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_2
XFILLER_0_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_214_ AXI_BRIDGE.clk _003_ net12 VGND VGND VPWR VPWR AXI_BRIDGE.state\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_145_ _089_ _038_ _046_ _052_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__and4_1
XFILLER_0_34_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_128_ counter\[8\] counter\[9\] _041_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_19 VGND VGND VPWR VPWR riscv_pipeline_top_19/HI M_AXI_ARADDR[5]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_149_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout12 net6 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_4
XFILLER_0_92_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_161_ _054_ _059_ _062_ VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput2 M_AXI_AWREADY VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_39_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_213_ AXI_BRIDGE.clk _000_ net13 VGND VGND VPWR VPWR AXI_BRIDGE.state\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_144_ counter\[12\] counter\[13\] counter\[14\] counter\[15\] VGND VGND VPWR VPWR
+ _052_ sky130_fd_sc_hd__and4_1
XFILLER_0_80_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_127_ _089_ _038_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout13 net6 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_2
XFILLER_0_77_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_160_ counter\[20\] counter\[21\] VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput3 M_AXI_BVALID VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_2
XFILLER_0_93_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_212_ AXI_BRIDGE.clk _002_ net12 VGND VGND VPWR VPWR AXI_BRIDGE.state\[0\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_108_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_143_ counter\[12\] counter\[13\] counter\[14\] _047_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__and4_1
XFILLER_0_80_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_126_ net137 _039_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_109_ net136 _085_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_871 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput4 M_AXI_RVALID VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_211_ clknet_1_0__leaf_clk _023_ net13 VGND VGND VPWR VPWR AXI_BRIDGE.clk sky130_fd_sc_hd__dfrtp_4
XFILLER_0_93_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_142_ net133 _050_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__xor2_1
XFILLER_0_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_125_ _040_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_108_ _087_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput5 M_AXI_WREADY VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_210_ clknet_1_0__leaf_clk _022_ net12 VGND VGND VPWR VPWR counter\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_141_ net138 _048_ _050_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_53_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_124_ _037_ _039_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_107_ _085_ _086_ VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput6 rst_n VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_160_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_140_ counter\[12\] counter\[13\] _047_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__and3_1
XFILLER_0_163_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_123_ _089_ _038_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_874 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_106_ counter\[1\] counter\[0\] VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_199_ clknet_1_1__leaf_clk _010_ net11 VGND VGND VPWR VPWR counter\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_122_ counter\[4\] counter\[5\] counter\[6\] counter\[7\] VGND VGND VPWR VPWR _038_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_68_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_105_ counter\[1\] counter\[0\] VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_198_ clknet_1_0__leaf_clk _009_ net11 VGND VGND VPWR VPWR counter\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_121_ counter\[4\] counter\[5\] counter\[6\] _089_ counter\[7\] VGND VGND VPWR VPWR
+ _037_ sky130_fd_sc_hd__a41o_1
XFILLER_0_68_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_104_ _084_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_197_ clknet_1_0__leaf_clk _008_ net10 VGND VGND VPWR VPWR counter\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_120_ net131 _092_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_103_ net2 AXI_BRIDGE.state\[3\] VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__and2b_1
XFILLER_0_62_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1 counter\[24\] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_196_ clknet_1_1__leaf_clk _007_ net10 VGND VGND VPWR VPWR counter\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_179_ _083_ VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_102_ AXI_BRIDGE.state\[2\] net5 _083_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2 counter\[0\] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_195_ clknet_1_0__leaf_clk _031_ net10 VGND VGND VPWR VPWR counter\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_985 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_178_ AXI_BRIDGE.state\[1\] net1 _071_ _073_ net8 VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__a32o_1
XFILLER_0_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_101_ net3 _082_ VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3 counter\[10\] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_194_ clknet_1_0__leaf_clk _030_ net10 VGND VGND VPWR VPWR counter\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_177_ _000_ _081_ _072_ VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__or3b_1
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_100_ AXI_BRIDGE.state\[5\] VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold4 counter\[22\] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_193_ clknet_1_0__leaf_clk _029_ net10 VGND VGND VPWR VPWR counter\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_942 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_176_ AXI_BRIDGE.state\[0\] AXI_BRIDGE.state\[4\] AXI_BRIDGE.state\[1\] VGND VGND
+ VPWR VPWR _072_ sky130_fd_sc_hd__or3_1
XFILLER_0_123_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_159_ net130 _060_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold5 counter\[20\] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_120 VGND VGND VPWR VPWR riscv_pipeline_top_120/HI led[5] sky130_fd_sc_hd__conb_1
XFILLER_0_158_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_192_ clknet_1_0__leaf_clk _028_ net10 VGND VGND VPWR VPWR counter\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_954 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_175_ _081_ VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_158_ _061_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold6 counter\[6\] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xriscv_pipeline_top_121 VGND VGND VPWR VPWR riscv_pipeline_top_121/HI led[6] sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_110 VGND VGND VPWR VPWR riscv_pipeline_top_110/HI M_AXI_WDATA[30]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_174_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_191_ clknet_1_0__leaf_clk _027_ net10 VGND VGND VPWR VPWR counter\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_899 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_966 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_174_ net127 VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_157_ _058_ _060_ VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold7 counter\[11\] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_209_ clknet_1_0__leaf_clk _021_ net12 VGND VGND VPWR VPWR counter\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_100 VGND VGND VPWR VPWR riscv_pipeline_top_100/HI M_AXI_WDATA[20]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_111 VGND VGND VPWR VPWR riscv_pipeline_top_111/HI M_AXI_WDATA[31]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_122 VGND VGND VPWR VPWR riscv_pipeline_top_122/HI led[7] sky130_fd_sc_hd__conb_1
XFILLER_0_58_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_190_ clknet_1_0__leaf_clk _026_ net10 VGND VGND VPWR VPWR counter\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_864 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_173_ net142 _070_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__xor2_1
XFILLER_0_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_818 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_156_ _054_ _059_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_973 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold8 counter\[14\] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_208_ clknet_1_1__leaf_clk _020_ net13 VGND VGND VPWR VPWR counter\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_139_ _048_ _049_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_101 VGND VGND VPWR VPWR riscv_pipeline_top_101/HI M_AXI_WDATA[21]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_112 VGND VGND VPWR VPWR riscv_pipeline_top_112/HI M_AXI_WSTRB[1]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_123 VGND VGND VPWR VPWR riscv_pipeline_top_123/HI led[8] sky130_fd_sc_hd__conb_1
XFILLER_0_89_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_172_ counter\[24\] _054_ _059_ _066_ VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__and4_1
XFILLER_0_80_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_155_ counter\[16\] counter\[17\] counter\[18\] counter\[19\] VGND VGND VPWR VPWR
+ _059_ sky130_fd_sc_hd__and4_2
XFILLER_0_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_985 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold9 counter\[18\] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_207_ clknet_1_1__leaf_clk _019_ net13 VGND VGND VPWR VPWR counter\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_138_ net140 _047_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_113 VGND VGND VPWR VPWR riscv_pipeline_top_113/HI M_AXI_WSTRB[2]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_124 VGND VGND VPWR VPWR riscv_pipeline_top_124/HI led[9] sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_102 VGND VGND VPWR VPWR riscv_pipeline_top_102/HI M_AXI_WDATA[22]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_89_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_861 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_171_ net126 _067_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__xor2_1
XFILLER_0_65_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_973 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_154_ counter\[16\] counter\[17\] counter\[18\] _054_ counter\[19\] VGND VGND VPWR
+ VPWR _058_ sky130_fd_sc_hd__a41o_1
XFILLER_0_150_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_206_ clknet_1_1__leaf_clk _018_ net13 VGND VGND VPWR VPWR counter\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_137_ counter\[12\] _047_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xriscv_pipeline_top_103 VGND VGND VPWR VPWR riscv_pipeline_top_103/HI M_AXI_WDATA[23]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_114 VGND VGND VPWR VPWR riscv_pipeline_top_114/HI M_AXI_WSTRB[3]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_125 VGND VGND VPWR VPWR M_AXI_WSTRB[0] riscv_pipeline_top_125/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_89_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_868 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_927 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_170_ _069_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_985 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_153_ net134 _055_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_205_ clknet_1_1__leaf_clk _016_ net12 VGND VGND VPWR VPWR counter\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_136_ net132 _045_ _047_ VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_104 VGND VGND VPWR VPWR riscv_pipeline_top_104/HI M_AXI_WDATA[24]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_115 VGND VGND VPWR VPWR riscv_pipeline_top_115/HI led[0] sky130_fd_sc_hd__conb_1
XFILLER_0_89_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_119_ _036_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_90 VGND VGND VPWR VPWR riscv_pipeline_top_90/HI M_AXI_WDATA[10]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_152_ _057_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_204_ clknet_1_1__leaf_clk _015_ net12 VGND VGND VPWR VPWR counter\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_135_ _089_ _038_ _046_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_105 VGND VGND VPWR VPWR riscv_pipeline_top_105/HI M_AXI_WDATA[25]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_116 VGND VGND VPWR VPWR riscv_pipeline_top_116/HI led[1] sky130_fd_sc_hd__conb_1
XFILLER_0_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_118_ _092_ _035_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_878 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_1 clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_80 VGND VGND VPWR VPWR riscv_pipeline_top_80/HI M_AXI_WDATA[0]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_91 VGND VGND VPWR VPWR riscv_pipeline_top_91/HI M_AXI_WDATA[11]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_20_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_220_ AXI_BRIDGE.clk _034_ net12 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_151_ _055_ _056_ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_203_ clknet_1_1__leaf_clk _014_ net11 VGND VGND VPWR VPWR counter\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_134_ counter\[8\] counter\[9\] counter\[10\] counter\[11\] VGND VGND VPWR VPWR _046_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_80_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xriscv_pipeline_top_106 VGND VGND VPWR VPWR riscv_pipeline_top_106/HI M_AXI_WDATA[26]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_101_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_117 VGND VGND VPWR VPWR riscv_pipeline_top_117/HI led[2] sky130_fd_sc_hd__conb_1
XFILLER_0_173_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_117_ counter\[4\] _089_ counter\[5\] VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_960 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xriscv_pipeline_top_70 VGND VGND VPWR VPWR riscv_pipeline_top_70/HI M_AXI_AWADDR[23]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_81 VGND VGND VPWR VPWR riscv_pipeline_top_81/HI M_AXI_WDATA[1]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_92 VGND VGND VPWR VPWR riscv_pipeline_top_92/HI M_AXI_WDATA[12]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_150_ counter\[16\] _054_ counter\[17\] VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__a21o_1
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_202_ clknet_1_1__leaf_clk _013_ net11 VGND VGND VPWR VPWR counter\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_133_ counter\[8\] counter\[9\] counter\[10\] _041_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__and4_1
XFILLER_0_80_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_107 VGND VGND VPWR VPWR riscv_pipeline_top_107/HI M_AXI_WDATA[27]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_118 VGND VGND VPWR VPWR riscv_pipeline_top_118/HI led[3] sky130_fd_sc_hd__conb_1
XFILLER_0_173_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_116_ counter\[4\] counter\[5\] _089_ VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__nand3_1
XFILLER_0_81_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_972 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_71 VGND VGND VPWR VPWR riscv_pipeline_top_71/HI M_AXI_AWADDR[24]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_82 VGND VGND VPWR VPWR riscv_pipeline_top_82/HI M_AXI_WDATA[2]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_60 VGND VGND VPWR VPWR riscv_pipeline_top_60/HI M_AXI_AWADDR[13]
+ sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_93 VGND VGND VPWR VPWR riscv_pipeline_top_93/HI M_AXI_WDATA[13]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_155_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_201_ clknet_1_1__leaf_clk _012_ net11 VGND VGND VPWR VPWR counter\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_132_ net128 _042_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xriscv_pipeline_top_119 VGND VGND VPWR VPWR riscv_pipeline_top_119/HI led[4] sky130_fd_sc_hd__conb_1
Xriscv_pipeline_top_108 VGND VGND VPWR VPWR riscv_pipeline_top_108/HI M_AXI_WDATA[28]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_173_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_115_ net139 _089_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__xor2_1
XFILLER_0_80_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_984 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
.ends

