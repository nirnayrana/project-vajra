module vajra_caravel_soc (wb_clk_i,
    wb_rst_i,
    io_in,
    io_oeb,
    io_out);
 input wb_clk_i;
 input wb_rst_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;

 wire _08226_;
 wire _71933_;
 wire _71934_;
 wire _71935_;
 wire _71936_;
 wire _71937_;
 wire _71938_;
 wire _71939_;
 wire _71940_;
 wire _71941_;
 wire _71942_;
 wire _71943_;
 wire _71944_;
 wire _71945_;
 wire _71946_;
 wire _71947_;
 wire _71948_;
 wire _71949_;
 wire _71950_;
 wire _71951_;
 wire _71952_;
 wire _71953_;
 wire _71954_;
 wire _71955_;
 wire \u_cpu.ALU.ALUResult[0] ;
 wire \u_cpu.ALU.ALUResult[10] ;
 wire \u_cpu.ALU.ALUResult[11] ;
 wire \u_cpu.ALU.ALUResult[12] ;
 wire \u_cpu.ALU.ALUResult[13] ;
 wire \u_cpu.ALU.ALUResult[14] ;
 wire \u_cpu.ALU.ALUResult[15] ;
 wire \u_cpu.ALU.ALUResult[16] ;
 wire \u_cpu.ALU.ALUResult[17] ;
 wire \u_cpu.ALU.ALUResult[18] ;
 wire \u_cpu.ALU.ALUResult[19] ;
 wire \u_cpu.ALU.ALUResult[1] ;
 wire \u_cpu.ALU.ALUResult[20] ;
 wire \u_cpu.ALU.ALUResult[21] ;
 wire \u_cpu.ALU.ALUResult[22] ;
 wire \u_cpu.ALU.ALUResult[23] ;
 wire \u_cpu.ALU.ALUResult[24] ;
 wire \u_cpu.ALU.ALUResult[25] ;
 wire \u_cpu.ALU.ALUResult[26] ;
 wire \u_cpu.ALU.ALUResult[27] ;
 wire \u_cpu.ALU.ALUResult[28] ;
 wire \u_cpu.ALU.ALUResult[29] ;
 wire \u_cpu.ALU.ALUResult[2] ;
 wire \u_cpu.ALU.ALUResult[30] ;
 wire \u_cpu.ALU.ALUResult[31] ;
 wire \u_cpu.ALU.ALUResult[3] ;
 wire \u_cpu.ALU.ALUResult[4] ;
 wire \u_cpu.ALU.ALUResult[5] ;
 wire \u_cpu.ALU.ALUResult[6] ;
 wire \u_cpu.ALU.ALUResult[7] ;
 wire \u_cpu.ALU.ALUResult[8] ;
 wire \u_cpu.ALU.ALUResult[9] ;
 wire \u_cpu.ALU.Product_Wallace[0] ;
 wire \u_cpu.ALU.Product_Wallace[10] ;
 wire \u_cpu.ALU.Product_Wallace[11] ;
 wire \u_cpu.ALU.Product_Wallace[12] ;
 wire \u_cpu.ALU.Product_Wallace[13] ;
 wire \u_cpu.ALU.Product_Wallace[14] ;
 wire \u_cpu.ALU.Product_Wallace[15] ;
 wire \u_cpu.ALU.Product_Wallace[16] ;
 wire \u_cpu.ALU.Product_Wallace[17] ;
 wire \u_cpu.ALU.Product_Wallace[18] ;
 wire \u_cpu.ALU.Product_Wallace[19] ;
 wire \u_cpu.ALU.Product_Wallace[1] ;
 wire \u_cpu.ALU.Product_Wallace[20] ;
 wire \u_cpu.ALU.Product_Wallace[21] ;
 wire \u_cpu.ALU.Product_Wallace[22] ;
 wire \u_cpu.ALU.Product_Wallace[23] ;
 wire \u_cpu.ALU.Product_Wallace[24] ;
 wire \u_cpu.ALU.Product_Wallace[25] ;
 wire \u_cpu.ALU.Product_Wallace[26] ;
 wire \u_cpu.ALU.Product_Wallace[27] ;
 wire \u_cpu.ALU.Product_Wallace[28] ;
 wire \u_cpu.ALU.Product_Wallace[29] ;
 wire \u_cpu.ALU.Product_Wallace[2] ;
 wire \u_cpu.ALU.Product_Wallace[30] ;
 wire \u_cpu.ALU.Product_Wallace[31] ;
 wire \u_cpu.ALU.Product_Wallace[3] ;
 wire \u_cpu.ALU.Product_Wallace[4] ;
 wire \u_cpu.ALU.Product_Wallace[5] ;
 wire \u_cpu.ALU.Product_Wallace[6] ;
 wire \u_cpu.ALU.Product_Wallace[7] ;
 wire \u_cpu.ALU.Product_Wallace[8] ;
 wire \u_cpu.ALU.Product_Wallace[9] ;
 wire \u_cpu.ALU.SrcA[0] ;
 wire \u_cpu.ALU.SrcA[10] ;
 wire \u_cpu.ALU.SrcA[11] ;
 wire \u_cpu.ALU.SrcA[12] ;
 wire \u_cpu.ALU.SrcA[13] ;
 wire \u_cpu.ALU.SrcA[14] ;
 wire \u_cpu.ALU.SrcA[15] ;
 wire \u_cpu.ALU.SrcA[16] ;
 wire \u_cpu.ALU.SrcA[17] ;
 wire \u_cpu.ALU.SrcA[18] ;
 wire \u_cpu.ALU.SrcA[19] ;
 wire \u_cpu.ALU.SrcA[1] ;
 wire \u_cpu.ALU.SrcA[20] ;
 wire \u_cpu.ALU.SrcA[21] ;
 wire \u_cpu.ALU.SrcA[22] ;
 wire \u_cpu.ALU.SrcA[23] ;
 wire \u_cpu.ALU.SrcA[24] ;
 wire \u_cpu.ALU.SrcA[25] ;
 wire \u_cpu.ALU.SrcA[26] ;
 wire \u_cpu.ALU.SrcA[27] ;
 wire \u_cpu.ALU.SrcA[28] ;
 wire \u_cpu.ALU.SrcA[29] ;
 wire \u_cpu.ALU.SrcA[2] ;
 wire \u_cpu.ALU.SrcA[30] ;
 wire \u_cpu.ALU.SrcA[31] ;
 wire \u_cpu.ALU.SrcA[3] ;
 wire \u_cpu.ALU.SrcA[4] ;
 wire \u_cpu.ALU.SrcA[5] ;
 wire \u_cpu.ALU.SrcA[6] ;
 wire \u_cpu.ALU.SrcA[7] ;
 wire \u_cpu.ALU.SrcA[8] ;
 wire \u_cpu.ALU.SrcA[9] ;
 wire \u_cpu.ALU.SrcB[0] ;
 wire \u_cpu.ALU.SrcB[10] ;
 wire \u_cpu.ALU.SrcB[11] ;
 wire \u_cpu.ALU.SrcB[12] ;
 wire \u_cpu.ALU.SrcB[13] ;
 wire \u_cpu.ALU.SrcB[14] ;
 wire \u_cpu.ALU.SrcB[15] ;
 wire \u_cpu.ALU.SrcB[16] ;
 wire \u_cpu.ALU.SrcB[17] ;
 wire \u_cpu.ALU.SrcB[18] ;
 wire \u_cpu.ALU.SrcB[19] ;
 wire \u_cpu.ALU.SrcB[1] ;
 wire \u_cpu.ALU.SrcB[20] ;
 wire \u_cpu.ALU.SrcB[21] ;
 wire \u_cpu.ALU.SrcB[22] ;
 wire \u_cpu.ALU.SrcB[23] ;
 wire \u_cpu.ALU.SrcB[24] ;
 wire \u_cpu.ALU.SrcB[25] ;
 wire \u_cpu.ALU.SrcB[26] ;
 wire \u_cpu.ALU.SrcB[27] ;
 wire \u_cpu.ALU.SrcB[28] ;
 wire \u_cpu.ALU.SrcB[29] ;
 wire \u_cpu.ALU.SrcB[2] ;
 wire \u_cpu.ALU.SrcB[30] ;
 wire \u_cpu.ALU.SrcB[31] ;
 wire \u_cpu.ALU.SrcB[3] ;
 wire \u_cpu.ALU.SrcB[4] ;
 wire \u_cpu.ALU.SrcB[5] ;
 wire \u_cpu.ALU.SrcB[6] ;
 wire \u_cpu.ALU.SrcB[7] ;
 wire \u_cpu.ALU.SrcB[8] ;
 wire \u_cpu.ALU.SrcB[9] ;
 wire \u_cpu.ALU._0000_ ;
 wire \u_cpu.ALU._0001_ ;
 wire \u_cpu.ALU._0002_ ;
 wire \u_cpu.ALU._0003_ ;
 wire \u_cpu.ALU._0004_ ;
 wire \u_cpu.ALU._0005_ ;
 wire \u_cpu.ALU._0006_ ;
 wire \u_cpu.ALU._0007_ ;
 wire \u_cpu.ALU._0008_ ;
 wire \u_cpu.ALU._0009_ ;
 wire \u_cpu.ALU._0010_ ;
 wire \u_cpu.ALU._0011_ ;
 wire \u_cpu.ALU._0012_ ;
 wire \u_cpu.ALU._0013_ ;
 wire \u_cpu.ALU._0014_ ;
 wire \u_cpu.ALU._0015_ ;
 wire \u_cpu.ALU._0016_ ;
 wire \u_cpu.ALU._0017_ ;
 wire \u_cpu.ALU._0018_ ;
 wire \u_cpu.ALU._0019_ ;
 wire \u_cpu.ALU._0020_ ;
 wire \u_cpu.ALU._0021_ ;
 wire \u_cpu.ALU._0022_ ;
 wire \u_cpu.ALU._0023_ ;
 wire \u_cpu.ALU._0024_ ;
 wire \u_cpu.ALU._0025_ ;
 wire \u_cpu.ALU._0026_ ;
 wire \u_cpu.ALU._0027_ ;
 wire \u_cpu.ALU._0028_ ;
 wire \u_cpu.ALU._0029_ ;
 wire \u_cpu.ALU._0030_ ;
 wire \u_cpu.ALU._0031_ ;
 wire \u_cpu.ALU._0032_ ;
 wire \u_cpu.ALU._0033_ ;
 wire \u_cpu.ALU._0034_ ;
 wire \u_cpu.ALU._0035_ ;
 wire \u_cpu.ALU._0036_ ;
 wire \u_cpu.ALU._0037_ ;
 wire \u_cpu.ALU._0038_ ;
 wire \u_cpu.ALU._0039_ ;
 wire \u_cpu.ALU._0040_ ;
 wire \u_cpu.ALU._0041_ ;
 wire \u_cpu.ALU._0042_ ;
 wire \u_cpu.ALU._0043_ ;
 wire \u_cpu.ALU._0044_ ;
 wire \u_cpu.ALU._0045_ ;
 wire \u_cpu.ALU._0046_ ;
 wire \u_cpu.ALU._0047_ ;
 wire \u_cpu.ALU._0048_ ;
 wire \u_cpu.ALU._0049_ ;
 wire \u_cpu.ALU._0050_ ;
 wire \u_cpu.ALU._0051_ ;
 wire \u_cpu.ALU._0052_ ;
 wire \u_cpu.ALU._0053_ ;
 wire \u_cpu.ALU._0054_ ;
 wire \u_cpu.ALU._0055_ ;
 wire \u_cpu.ALU._0056_ ;
 wire \u_cpu.ALU._0057_ ;
 wire \u_cpu.ALU._0058_ ;
 wire \u_cpu.ALU._0059_ ;
 wire \u_cpu.ALU._0060_ ;
 wire \u_cpu.ALU._0061_ ;
 wire \u_cpu.ALU._0062_ ;
 wire \u_cpu.ALU._0063_ ;
 wire \u_cpu.ALU._0064_ ;
 wire \u_cpu.ALU._0065_ ;
 wire \u_cpu.ALU._0066_ ;
 wire \u_cpu.ALU._0067_ ;
 wire \u_cpu.ALU._0068_ ;
 wire \u_cpu.ALU._0069_ ;
 wire \u_cpu.ALU._0070_ ;
 wire \u_cpu.ALU._0071_ ;
 wire \u_cpu.ALU._0072_ ;
 wire \u_cpu.ALU._0073_ ;
 wire \u_cpu.ALU._0074_ ;
 wire \u_cpu.ALU._0075_ ;
 wire \u_cpu.ALU._0076_ ;
 wire \u_cpu.ALU._0077_ ;
 wire \u_cpu.ALU._0078_ ;
 wire \u_cpu.ALU._0079_ ;
 wire \u_cpu.ALU._0080_ ;
 wire \u_cpu.ALU._0081_ ;
 wire \u_cpu.ALU._0082_ ;
 wire \u_cpu.ALU._0083_ ;
 wire \u_cpu.ALU._0084_ ;
 wire \u_cpu.ALU._0085_ ;
 wire \u_cpu.ALU._0086_ ;
 wire \u_cpu.ALU._0087_ ;
 wire \u_cpu.ALU._0088_ ;
 wire \u_cpu.ALU._0089_ ;
 wire \u_cpu.ALU._0090_ ;
 wire \u_cpu.ALU._0091_ ;
 wire \u_cpu.ALU._0092_ ;
 wire \u_cpu.ALU._0093_ ;
 wire \u_cpu.ALU._0094_ ;
 wire \u_cpu.ALU._0095_ ;
 wire \u_cpu.ALU._0096_ ;
 wire \u_cpu.ALU._0097_ ;
 wire \u_cpu.ALU._0098_ ;
 wire \u_cpu.ALU._0099_ ;
 wire \u_cpu.ALU._0100_ ;
 wire \u_cpu.ALU._0101_ ;
 wire \u_cpu.ALU._0102_ ;
 wire \u_cpu.ALU._0103_ ;
 wire \u_cpu.ALU._0104_ ;
 wire \u_cpu.ALU._0105_ ;
 wire \u_cpu.ALU._0106_ ;
 wire \u_cpu.ALU._0107_ ;
 wire \u_cpu.ALU._0108_ ;
 wire \u_cpu.ALU._0109_ ;
 wire \u_cpu.ALU._0110_ ;
 wire \u_cpu.ALU._0111_ ;
 wire \u_cpu.ALU._0112_ ;
 wire \u_cpu.ALU._0113_ ;
 wire \u_cpu.ALU._0114_ ;
 wire \u_cpu.ALU._0115_ ;
 wire \u_cpu.ALU._0116_ ;
 wire \u_cpu.ALU._0117_ ;
 wire \u_cpu.ALU._0118_ ;
 wire \u_cpu.ALU._0119_ ;
 wire \u_cpu.ALU._0120_ ;
 wire \u_cpu.ALU._0121_ ;
 wire \u_cpu.ALU._0122_ ;
 wire \u_cpu.ALU._0123_ ;
 wire \u_cpu.ALU._0124_ ;
 wire \u_cpu.ALU._0125_ ;
 wire \u_cpu.ALU._0126_ ;
 wire \u_cpu.ALU._0127_ ;
 wire \u_cpu.ALU._0128_ ;
 wire \u_cpu.ALU._0129_ ;
 wire \u_cpu.ALU._0130_ ;
 wire \u_cpu.ALU._0131_ ;
 wire \u_cpu.ALU._0132_ ;
 wire \u_cpu.ALU._0133_ ;
 wire \u_cpu.ALU._0134_ ;
 wire \u_cpu.ALU._0135_ ;
 wire \u_cpu.ALU._0136_ ;
 wire \u_cpu.ALU._0137_ ;
 wire \u_cpu.ALU._0138_ ;
 wire \u_cpu.ALU._0139_ ;
 wire \u_cpu.ALU._0140_ ;
 wire \u_cpu.ALU._0141_ ;
 wire \u_cpu.ALU._0142_ ;
 wire \u_cpu.ALU._0143_ ;
 wire \u_cpu.ALU._0144_ ;
 wire \u_cpu.ALU._0145_ ;
 wire \u_cpu.ALU._0146_ ;
 wire \u_cpu.ALU._0147_ ;
 wire \u_cpu.ALU._0148_ ;
 wire \u_cpu.ALU._0149_ ;
 wire \u_cpu.ALU._0150_ ;
 wire \u_cpu.ALU._0151_ ;
 wire \u_cpu.ALU._0152_ ;
 wire \u_cpu.ALU._0153_ ;
 wire \u_cpu.ALU._0154_ ;
 wire \u_cpu.ALU._0155_ ;
 wire \u_cpu.ALU._0156_ ;
 wire \u_cpu.ALU._0157_ ;
 wire \u_cpu.ALU._0158_ ;
 wire \u_cpu.ALU._0159_ ;
 wire \u_cpu.ALU._0160_ ;
 wire \u_cpu.ALU._0161_ ;
 wire \u_cpu.ALU._0162_ ;
 wire \u_cpu.ALU._0163_ ;
 wire \u_cpu.ALU._0164_ ;
 wire \u_cpu.ALU._0165_ ;
 wire \u_cpu.ALU._0166_ ;
 wire \u_cpu.ALU._0167_ ;
 wire \u_cpu.ALU._0168_ ;
 wire \u_cpu.ALU._0169_ ;
 wire \u_cpu.ALU._0170_ ;
 wire \u_cpu.ALU._0171_ ;
 wire \u_cpu.ALU._0172_ ;
 wire \u_cpu.ALU._0173_ ;
 wire \u_cpu.ALU._0174_ ;
 wire \u_cpu.ALU._0175_ ;
 wire \u_cpu.ALU._0176_ ;
 wire \u_cpu.ALU._0177_ ;
 wire \u_cpu.ALU._0178_ ;
 wire \u_cpu.ALU._0179_ ;
 wire \u_cpu.ALU._0180_ ;
 wire \u_cpu.ALU._0181_ ;
 wire \u_cpu.ALU._0182_ ;
 wire \u_cpu.ALU._0183_ ;
 wire \u_cpu.ALU._0184_ ;
 wire \u_cpu.ALU._0185_ ;
 wire \u_cpu.ALU._0186_ ;
 wire \u_cpu.ALU._0187_ ;
 wire \u_cpu.ALU._0188_ ;
 wire \u_cpu.ALU._0189_ ;
 wire \u_cpu.ALU._0190_ ;
 wire \u_cpu.ALU._0191_ ;
 wire \u_cpu.ALU._0192_ ;
 wire \u_cpu.ALU._0193_ ;
 wire \u_cpu.ALU._0194_ ;
 wire \u_cpu.ALU._0195_ ;
 wire \u_cpu.ALU._0196_ ;
 wire \u_cpu.ALU._0197_ ;
 wire \u_cpu.ALU._0198_ ;
 wire \u_cpu.ALU._0199_ ;
 wire \u_cpu.ALU._0200_ ;
 wire \u_cpu.ALU._0201_ ;
 wire \u_cpu.ALU._0202_ ;
 wire \u_cpu.ALU._0203_ ;
 wire \u_cpu.ALU._0204_ ;
 wire \u_cpu.ALU._0205_ ;
 wire \u_cpu.ALU._0206_ ;
 wire \u_cpu.ALU._0207_ ;
 wire \u_cpu.ALU._0208_ ;
 wire \u_cpu.ALU._0209_ ;
 wire \u_cpu.ALU._0210_ ;
 wire \u_cpu.ALU._0211_ ;
 wire \u_cpu.ALU._0212_ ;
 wire \u_cpu.ALU._0213_ ;
 wire \u_cpu.ALU._0214_ ;
 wire \u_cpu.ALU._0215_ ;
 wire \u_cpu.ALU._0216_ ;
 wire \u_cpu.ALU._0217_ ;
 wire \u_cpu.ALU._0218_ ;
 wire \u_cpu.ALU._0219_ ;
 wire \u_cpu.ALU._0220_ ;
 wire \u_cpu.ALU._0221_ ;
 wire \u_cpu.ALU._0222_ ;
 wire \u_cpu.ALU._0223_ ;
 wire \u_cpu.ALU._0224_ ;
 wire \u_cpu.ALU._0225_ ;
 wire \u_cpu.ALU._0226_ ;
 wire \u_cpu.ALU._0227_ ;
 wire \u_cpu.ALU._0228_ ;
 wire \u_cpu.ALU._0229_ ;
 wire \u_cpu.ALU._0230_ ;
 wire \u_cpu.ALU._0231_ ;
 wire \u_cpu.ALU._0232_ ;
 wire \u_cpu.ALU._0233_ ;
 wire \u_cpu.ALU._0234_ ;
 wire \u_cpu.ALU._0235_ ;
 wire \u_cpu.ALU._0236_ ;
 wire \u_cpu.ALU._0237_ ;
 wire \u_cpu.ALU._0238_ ;
 wire \u_cpu.ALU._0239_ ;
 wire \u_cpu.ALU._0240_ ;
 wire \u_cpu.ALU._0241_ ;
 wire \u_cpu.ALU._0242_ ;
 wire \u_cpu.ALU._0243_ ;
 wire \u_cpu.ALU._0244_ ;
 wire \u_cpu.ALU._0245_ ;
 wire \u_cpu.ALU._0246_ ;
 wire \u_cpu.ALU._0247_ ;
 wire \u_cpu.ALU._0248_ ;
 wire \u_cpu.ALU._0249_ ;
 wire \u_cpu.ALU._0250_ ;
 wire \u_cpu.ALU._0251_ ;
 wire \u_cpu.ALU._0252_ ;
 wire \u_cpu.ALU._0253_ ;
 wire \u_cpu.ALU._0254_ ;
 wire \u_cpu.ALU._0255_ ;
 wire \u_cpu.ALU._0256_ ;
 wire \u_cpu.ALU._0257_ ;
 wire \u_cpu.ALU._0258_ ;
 wire \u_cpu.ALU._0259_ ;
 wire \u_cpu.ALU._0260_ ;
 wire \u_cpu.ALU._0261_ ;
 wire \u_cpu.ALU._0262_ ;
 wire \u_cpu.ALU._0263_ ;
 wire \u_cpu.ALU._0264_ ;
 wire \u_cpu.ALU._0265_ ;
 wire \u_cpu.ALU._0266_ ;
 wire \u_cpu.ALU._0267_ ;
 wire \u_cpu.ALU._0268_ ;
 wire \u_cpu.ALU._0269_ ;
 wire \u_cpu.ALU._0270_ ;
 wire \u_cpu.ALU._0271_ ;
 wire \u_cpu.ALU._0272_ ;
 wire \u_cpu.ALU._0273_ ;
 wire \u_cpu.ALU._0274_ ;
 wire \u_cpu.ALU._0275_ ;
 wire \u_cpu.ALU._0276_ ;
 wire \u_cpu.ALU._0277_ ;
 wire \u_cpu.ALU._0278_ ;
 wire \u_cpu.ALU._0279_ ;
 wire \u_cpu.ALU._0280_ ;
 wire \u_cpu.ALU._0281_ ;
 wire \u_cpu.ALU._0282_ ;
 wire \u_cpu.ALU._0283_ ;
 wire \u_cpu.ALU._0284_ ;
 wire \u_cpu.ALU._0285_ ;
 wire \u_cpu.ALU._0286_ ;
 wire \u_cpu.ALU._0287_ ;
 wire \u_cpu.ALU._0288_ ;
 wire \u_cpu.ALU._0289_ ;
 wire \u_cpu.ALU._0290_ ;
 wire \u_cpu.ALU._0291_ ;
 wire \u_cpu.ALU._0292_ ;
 wire \u_cpu.ALU._0293_ ;
 wire \u_cpu.ALU._0294_ ;
 wire \u_cpu.ALU._0295_ ;
 wire \u_cpu.ALU._0296_ ;
 wire \u_cpu.ALU._0297_ ;
 wire \u_cpu.ALU._0298_ ;
 wire \u_cpu.ALU._0299_ ;
 wire \u_cpu.ALU._0300_ ;
 wire \u_cpu.ALU._0301_ ;
 wire \u_cpu.ALU._0302_ ;
 wire \u_cpu.ALU._0303_ ;
 wire \u_cpu.ALU._0304_ ;
 wire \u_cpu.ALU._0305_ ;
 wire \u_cpu.ALU._0306_ ;
 wire \u_cpu.ALU._0307_ ;
 wire \u_cpu.ALU._0308_ ;
 wire \u_cpu.ALU._0309_ ;
 wire \u_cpu.ALU._0310_ ;
 wire \u_cpu.ALU._0311_ ;
 wire \u_cpu.ALU._0312_ ;
 wire \u_cpu.ALU._0313_ ;
 wire \u_cpu.ALU._0314_ ;
 wire \u_cpu.ALU._0315_ ;
 wire \u_cpu.ALU._0316_ ;
 wire \u_cpu.ALU._0317_ ;
 wire \u_cpu.ALU._0318_ ;
 wire \u_cpu.ALU._0319_ ;
 wire \u_cpu.ALU._0320_ ;
 wire \u_cpu.ALU._0321_ ;
 wire \u_cpu.ALU._0322_ ;
 wire \u_cpu.ALU._0323_ ;
 wire \u_cpu.ALU._0324_ ;
 wire \u_cpu.ALU._0325_ ;
 wire \u_cpu.ALU._0326_ ;
 wire \u_cpu.ALU._0327_ ;
 wire \u_cpu.ALU._0328_ ;
 wire \u_cpu.ALU._0329_ ;
 wire \u_cpu.ALU._0330_ ;
 wire \u_cpu.ALU._0331_ ;
 wire \u_cpu.ALU._0332_ ;
 wire \u_cpu.ALU._0333_ ;
 wire \u_cpu.ALU._0334_ ;
 wire \u_cpu.ALU._0335_ ;
 wire \u_cpu.ALU._0336_ ;
 wire \u_cpu.ALU._0337_ ;
 wire \u_cpu.ALU._0338_ ;
 wire \u_cpu.ALU._0339_ ;
 wire \u_cpu.ALU._0340_ ;
 wire \u_cpu.ALU._0341_ ;
 wire \u_cpu.ALU._0342_ ;
 wire \u_cpu.ALU._0343_ ;
 wire \u_cpu.ALU._0344_ ;
 wire \u_cpu.ALU._0345_ ;
 wire \u_cpu.ALU._0346_ ;
 wire \u_cpu.ALU._0347_ ;
 wire \u_cpu.ALU._0348_ ;
 wire \u_cpu.ALU._0349_ ;
 wire \u_cpu.ALU._0350_ ;
 wire \u_cpu.ALU._0351_ ;
 wire \u_cpu.ALU._0352_ ;
 wire \u_cpu.ALU._0353_ ;
 wire \u_cpu.ALU._0354_ ;
 wire \u_cpu.ALU._0355_ ;
 wire \u_cpu.ALU._0356_ ;
 wire \u_cpu.ALU._0357_ ;
 wire \u_cpu.ALU._0358_ ;
 wire \u_cpu.ALU._0359_ ;
 wire \u_cpu.ALU._0360_ ;
 wire \u_cpu.ALU._0361_ ;
 wire \u_cpu.ALU._0362_ ;
 wire \u_cpu.ALU._0363_ ;
 wire \u_cpu.ALU._0364_ ;
 wire \u_cpu.ALU._0365_ ;
 wire \u_cpu.ALU._0366_ ;
 wire \u_cpu.ALU._0367_ ;
 wire \u_cpu.ALU._0368_ ;
 wire \u_cpu.ALU._0369_ ;
 wire \u_cpu.ALU._0370_ ;
 wire \u_cpu.ALU._0371_ ;
 wire \u_cpu.ALU._0372_ ;
 wire \u_cpu.ALU._0373_ ;
 wire \u_cpu.ALU._0374_ ;
 wire \u_cpu.ALU._0375_ ;
 wire \u_cpu.ALU._0376_ ;
 wire \u_cpu.ALU._0377_ ;
 wire \u_cpu.ALU._0378_ ;
 wire \u_cpu.ALU._0379_ ;
 wire \u_cpu.ALU._0380_ ;
 wire \u_cpu.ALU._0381_ ;
 wire \u_cpu.ALU._0382_ ;
 wire \u_cpu.ALU._0383_ ;
 wire \u_cpu.ALU._0384_ ;
 wire \u_cpu.ALU._0385_ ;
 wire \u_cpu.ALU._0386_ ;
 wire \u_cpu.ALU._0387_ ;
 wire \u_cpu.ALU._0388_ ;
 wire \u_cpu.ALU._0389_ ;
 wire \u_cpu.ALU._0390_ ;
 wire \u_cpu.ALU._0391_ ;
 wire \u_cpu.ALU._0392_ ;
 wire \u_cpu.ALU._0393_ ;
 wire \u_cpu.ALU._0394_ ;
 wire \u_cpu.ALU._0395_ ;
 wire \u_cpu.ALU._0396_ ;
 wire \u_cpu.ALU._0397_ ;
 wire \u_cpu.ALU._0398_ ;
 wire \u_cpu.ALU._0399_ ;
 wire \u_cpu.ALU._0400_ ;
 wire \u_cpu.ALU._0401_ ;
 wire \u_cpu.ALU._0402_ ;
 wire \u_cpu.ALU._0403_ ;
 wire \u_cpu.ALU._0404_ ;
 wire \u_cpu.ALU._0405_ ;
 wire \u_cpu.ALU._0406_ ;
 wire \u_cpu.ALU._0407_ ;
 wire \u_cpu.ALU._0408_ ;
 wire \u_cpu.ALU._0409_ ;
 wire \u_cpu.ALU._0410_ ;
 wire \u_cpu.ALU._0411_ ;
 wire \u_cpu.ALU._0412_ ;
 wire \u_cpu.ALU._0413_ ;
 wire \u_cpu.ALU._0414_ ;
 wire \u_cpu.ALU._0415_ ;
 wire \u_cpu.ALU._0416_ ;
 wire \u_cpu.ALU._0417_ ;
 wire \u_cpu.ALU._0418_ ;
 wire \u_cpu.ALU._0419_ ;
 wire \u_cpu.ALU._0420_ ;
 wire \u_cpu.ALU._0421_ ;
 wire \u_cpu.ALU._0422_ ;
 wire \u_cpu.ALU._0423_ ;
 wire \u_cpu.ALU._0424_ ;
 wire \u_cpu.ALU._0425_ ;
 wire \u_cpu.ALU._0426_ ;
 wire \u_cpu.ALU._0427_ ;
 wire \u_cpu.ALU._0428_ ;
 wire \u_cpu.ALU._0429_ ;
 wire \u_cpu.ALU._0430_ ;
 wire \u_cpu.ALU._0431_ ;
 wire \u_cpu.ALU._0432_ ;
 wire \u_cpu.ALU._0433_ ;
 wire \u_cpu.ALU._0434_ ;
 wire \u_cpu.ALU._0435_ ;
 wire \u_cpu.ALU._0436_ ;
 wire \u_cpu.ALU._0437_ ;
 wire \u_cpu.ALU._0438_ ;
 wire \u_cpu.ALU._0439_ ;
 wire \u_cpu.ALU._0440_ ;
 wire \u_cpu.ALU._0441_ ;
 wire \u_cpu.ALU._0442_ ;
 wire \u_cpu.ALU._0443_ ;
 wire \u_cpu.ALU._0444_ ;
 wire \u_cpu.ALU._0445_ ;
 wire \u_cpu.ALU._0446_ ;
 wire \u_cpu.ALU._0447_ ;
 wire \u_cpu.ALU._0448_ ;
 wire \u_cpu.ALU._0449_ ;
 wire \u_cpu.ALU._0450_ ;
 wire \u_cpu.ALU._0451_ ;
 wire \u_cpu.ALU._0452_ ;
 wire \u_cpu.ALU._0453_ ;
 wire \u_cpu.ALU._0454_ ;
 wire \u_cpu.ALU._0455_ ;
 wire \u_cpu.ALU._0456_ ;
 wire \u_cpu.ALU._0457_ ;
 wire \u_cpu.ALU._0458_ ;
 wire \u_cpu.ALU._0459_ ;
 wire \u_cpu.ALU._0460_ ;
 wire \u_cpu.ALU._0461_ ;
 wire \u_cpu.ALU._0462_ ;
 wire \u_cpu.ALU._0463_ ;
 wire \u_cpu.ALU._0464_ ;
 wire \u_cpu.ALU._0465_ ;
 wire \u_cpu.ALU._0466_ ;
 wire \u_cpu.ALU._0467_ ;
 wire \u_cpu.ALU._0468_ ;
 wire \u_cpu.ALU._0469_ ;
 wire \u_cpu.ALU._0470_ ;
 wire \u_cpu.ALU._0471_ ;
 wire \u_cpu.ALU._0472_ ;
 wire \u_cpu.ALU._0473_ ;
 wire \u_cpu.ALU._0474_ ;
 wire \u_cpu.ALU._0475_ ;
 wire \u_cpu.ALU._0476_ ;
 wire \u_cpu.ALU._0477_ ;
 wire \u_cpu.ALU._0478_ ;
 wire \u_cpu.ALU._0479_ ;
 wire \u_cpu.ALU._0480_ ;
 wire \u_cpu.ALU._0481_ ;
 wire \u_cpu.ALU._0482_ ;
 wire \u_cpu.ALU._0483_ ;
 wire \u_cpu.ALU._0484_ ;
 wire \u_cpu.ALU._0485_ ;
 wire \u_cpu.ALU._0486_ ;
 wire \u_cpu.ALU._0487_ ;
 wire \u_cpu.ALU._0488_ ;
 wire \u_cpu.ALU._0489_ ;
 wire \u_cpu.ALU._0490_ ;
 wire \u_cpu.ALU._0491_ ;
 wire \u_cpu.ALU._0492_ ;
 wire \u_cpu.ALU._0493_ ;
 wire \u_cpu.ALU._0494_ ;
 wire \u_cpu.ALU._0495_ ;
 wire \u_cpu.ALU._0496_ ;
 wire \u_cpu.ALU._0507_ ;
 wire \u_cpu.ALU._0515_ ;
 wire \u_cpu.ALU._0516_ ;
 wire \u_cpu.ALU._0517_ ;
 wire \u_cpu.ALU._0518_ ;
 wire \u_cpu.ALU._0519_ ;
 wire \u_cpu.ALU._0520_ ;
 wire \u_cpu.ALU._0521_ ;
 wire \u_cpu.ALU._0522_ ;
 wire \u_cpu.ALU._0523_ ;
 wire \u_cpu.ALU._0524_ ;
 wire \u_cpu.ALU._0525_ ;
 wire \u_cpu.ALU._0526_ ;
 wire \u_cpu.ALU._0527_ ;
 wire \u_cpu.ALU._0528_ ;
 wire \u_cpu.ALU._0529_ ;
 wire \u_cpu.ALU._0530_ ;
 wire \u_cpu.ALU._0531_ ;
 wire \u_cpu.ALU._0532_ ;
 wire \u_cpu.ALU._0533_ ;
 wire \u_cpu.ALU._0534_ ;
 wire \u_cpu.ALU._0535_ ;
 wire \u_cpu.ALU._0536_ ;
 wire \u_cpu.ALU._0537_ ;
 wire \u_cpu.ALU._0538_ ;
 wire \u_cpu.ALU._0539_ ;
 wire \u_cpu.ALU._0540_ ;
 wire \u_cpu.ALU._0541_ ;
 wire \u_cpu.ALU._0542_ ;
 wire \u_cpu.ALU._0543_ ;
 wire \u_cpu.ALU._0544_ ;
 wire \u_cpu.ALU._0545_ ;
 wire \u_cpu.ALU._0546_ ;
 wire \u_cpu.ALU._0547_ ;
 wire \u_cpu.ALU._0548_ ;
 wire \u_cpu.ALU._0549_ ;
 wire \u_cpu.ALU._0550_ ;
 wire \u_cpu.ALU._0551_ ;
 wire \u_cpu.ALU._0552_ ;
 wire \u_cpu.ALU._0553_ ;
 wire \u_cpu.ALU._0554_ ;
 wire \u_cpu.ALU._0555_ ;
 wire \u_cpu.ALU._0556_ ;
 wire \u_cpu.ALU._0557_ ;
 wire \u_cpu.ALU._0558_ ;
 wire \u_cpu.ALU._0559_ ;
 wire \u_cpu.ALU._0560_ ;
 wire \u_cpu.ALU._0561_ ;
 wire \u_cpu.ALU._0562_ ;
 wire \u_cpu.ALU._0563_ ;
 wire \u_cpu.ALU._0564_ ;
 wire \u_cpu.ALU._0565_ ;
 wire \u_cpu.ALU._0566_ ;
 wire \u_cpu.ALU._0567_ ;
 wire \u_cpu.ALU._0568_ ;
 wire \u_cpu.ALU._0569_ ;
 wire \u_cpu.ALU._0570_ ;
 wire \u_cpu.ALU._0571_ ;
 wire \u_cpu.ALU._0572_ ;
 wire \u_cpu.ALU._0573_ ;
 wire \u_cpu.ALU._0574_ ;
 wire \u_cpu.ALU._0575_ ;
 wire \u_cpu.ALU._0576_ ;
 wire \u_cpu.ALU._0577_ ;
 wire \u_cpu.ALU._0578_ ;
 wire \u_cpu.ALU._0579_ ;
 wire \u_cpu.ALU._0580_ ;
 wire \u_cpu.ALU._0581_ ;
 wire \u_cpu.ALU._0582_ ;
 wire \u_cpu.ALU._0583_ ;
 wire \u_cpu.ALU._0584_ ;
 wire \u_cpu.ALU._0585_ ;
 wire \u_cpu.ALU._0586_ ;
 wire \u_cpu.ALU._0587_ ;
 wire \u_cpu.ALU._0588_ ;
 wire \u_cpu.ALU._0589_ ;
 wire \u_cpu.ALU._0590_ ;
 wire \u_cpu.ALU._0591_ ;
 wire \u_cpu.ALU._0592_ ;
 wire \u_cpu.ALU._0593_ ;
 wire \u_cpu.ALU._0594_ ;
 wire \u_cpu.ALU._0595_ ;
 wire \u_cpu.ALU._0596_ ;
 wire \u_cpu.ALU._0597_ ;
 wire \u_cpu.ALU._0598_ ;
 wire \u_cpu.ALU._0599_ ;
 wire \u_cpu.ALU._0600_ ;
 wire \u_cpu.ALU._0601_ ;
 wire \u_cpu.ALU._0602_ ;
 wire \u_cpu.ALU._0603_ ;
 wire \u_cpu.ALU._0604_ ;
 wire \u_cpu.ALU._0605_ ;
 wire \u_cpu.ALU._0606_ ;
 wire \u_cpu.ALU._0607_ ;
 wire \u_cpu.ALU._0608_ ;
 wire \u_cpu.ALU._0609_ ;
 wire \u_cpu.ALU._0610_ ;
 wire \u_cpu.ALU._0611_ ;
 wire \u_cpu.ALU._0612_ ;
 wire \u_cpu.ALU._0613_ ;
 wire \u_cpu.ALU._0614_ ;
 wire \u_cpu.ALU._0615_ ;
 wire \u_cpu.ALU._0616_ ;
 wire \u_cpu.ALU._0617_ ;
 wire \u_cpu.ALU._0618_ ;
 wire \u_cpu.ALU._0619_ ;
 wire \u_cpu.ALU._0620_ ;
 wire \u_cpu.ALU._0621_ ;
 wire \u_cpu.ALU._0622_ ;
 wire \u_cpu.ALU._0623_ ;
 wire \u_cpu.ALU._0624_ ;
 wire \u_cpu.ALU._0625_ ;
 wire \u_cpu.ALU._0626_ ;
 wire \u_cpu.ALU._0627_ ;
 wire \u_cpu.ALU._0628_ ;
 wire \u_cpu.ALU._0629_ ;
 wire \u_cpu.ALU._0630_ ;
 wire \u_cpu.ALU._0631_ ;
 wire \u_cpu.ALU._0632_ ;
 wire \u_cpu.ALU._0633_ ;
 wire \u_cpu.ALU._0634_ ;
 wire \u_cpu.ALU._0635_ ;
 wire \u_cpu.ALU._0636_ ;
 wire \u_cpu.ALU._0637_ ;
 wire \u_cpu.ALU._0638_ ;
 wire \u_cpu.ALU._0639_ ;
 wire \u_cpu.ALU._0640_ ;
 wire \u_cpu.ALU._0641_ ;
 wire \u_cpu.ALU._0642_ ;
 wire \u_cpu.ALU._0643_ ;
 wire \u_cpu.ALU._0644_ ;
 wire \u_cpu.ALU._0645_ ;
 wire \u_cpu.ALU._0646_ ;
 wire \u_cpu.ALU._0647_ ;
 wire \u_cpu.ALU._0648_ ;
 wire \u_cpu.ALU._0649_ ;
 wire \u_cpu.ALU._0650_ ;
 wire \u_cpu.ALU._0651_ ;
 wire \u_cpu.ALU._0652_ ;
 wire \u_cpu.ALU._0653_ ;
 wire \u_cpu.ALU._0654_ ;
 wire \u_cpu.ALU._0655_ ;
 wire \u_cpu.ALU._0656_ ;
 wire \u_cpu.ALU._0657_ ;
 wire \u_cpu.ALU._0658_ ;
 wire \u_cpu.ALU._0659_ ;
 wire \u_cpu.ALU._0660_ ;
 wire \u_cpu.ALU._0661_ ;
 wire \u_cpu.ALU._0662_ ;
 wire \u_cpu.ALU._0663_ ;
 wire \u_cpu.ALU._0664_ ;
 wire \u_cpu.ALU._0665_ ;
 wire \u_cpu.ALU._0666_ ;
 wire \u_cpu.ALU._0667_ ;
 wire \u_cpu.ALU._0668_ ;
 wire \u_cpu.ALU._0669_ ;
 wire \u_cpu.ALU._0670_ ;
 wire \u_cpu.ALU._0671_ ;
 wire \u_cpu.ALU._0672_ ;
 wire \u_cpu.ALU._0673_ ;
 wire \u_cpu.ALU._0674_ ;
 wire \u_cpu.ALU._0675_ ;
 wire \u_cpu.ALU._0676_ ;
 wire \u_cpu.ALU._0677_ ;
 wire \u_cpu.ALU._0678_ ;
 wire \u_cpu.ALU._0679_ ;
 wire \u_cpu.ALU._0680_ ;
 wire \u_cpu.ALU._0681_ ;
 wire \u_cpu.ALU._0682_ ;
 wire \u_cpu.ALU._0683_ ;
 wire \u_cpu.ALU._0684_ ;
 wire \u_cpu.ALU._0685_ ;
 wire \u_cpu.ALU._0686_ ;
 wire \u_cpu.ALU._0687_ ;
 wire \u_cpu.ALU._0688_ ;
 wire \u_cpu.ALU._0689_ ;
 wire \u_cpu.ALU._0690_ ;
 wire \u_cpu.ALU._0691_ ;
 wire \u_cpu.ALU._0692_ ;
 wire \u_cpu.ALU._0693_ ;
 wire \u_cpu.ALU._0694_ ;
 wire \u_cpu.ALU._0695_ ;
 wire \u_cpu.ALU._0696_ ;
 wire \u_cpu.ALU._0697_ ;
 wire \u_cpu.ALU._0698_ ;
 wire \u_cpu.ALU._0699_ ;
 wire \u_cpu.ALU._0700_ ;
 wire \u_cpu.ALU._0701_ ;
 wire \u_cpu.ALU._0702_ ;
 wire \u_cpu.ALU._0703_ ;
 wire \u_cpu.ALU._0704_ ;
 wire \u_cpu.ALU._0705_ ;
 wire \u_cpu.ALU._0706_ ;
 wire \u_cpu.ALU._0707_ ;
 wire \u_cpu.ALU._0708_ ;
 wire \u_cpu.ALU._0709_ ;
 wire \u_cpu.ALU._0710_ ;
 wire \u_cpu.ALU._0711_ ;
 wire \u_cpu.ALU._0712_ ;
 wire \u_cpu.ALU._0713_ ;
 wire \u_cpu.ALU._0714_ ;
 wire \u_cpu.ALU._0715_ ;
 wire \u_cpu.ALU._0716_ ;
 wire \u_cpu.ALU._0717_ ;
 wire \u_cpu.ALU._0718_ ;
 wire \u_cpu.ALU._0719_ ;
 wire \u_cpu.ALU._0720_ ;
 wire \u_cpu.ALU._0721_ ;
 wire \u_cpu.ALU._0722_ ;
 wire \u_cpu.ALU._0723_ ;
 wire \u_cpu.ALU._0724_ ;
 wire \u_cpu.ALU._0725_ ;
 wire \u_cpu.ALU._0726_ ;
 wire \u_cpu.ALU._0727_ ;
 wire \u_cpu.ALU._0728_ ;
 wire \u_cpu.ALU._0729_ ;
 wire \u_cpu.ALU._0730_ ;
 wire \u_cpu.ALU._0731_ ;
 wire \u_cpu.ALU._0732_ ;
 wire \u_cpu.ALU._0733_ ;
 wire \u_cpu.ALU._0734_ ;
 wire \u_cpu.ALU._0735_ ;
 wire \u_cpu.ALU._0736_ ;
 wire \u_cpu.ALU._0737_ ;
 wire \u_cpu.ALU._0738_ ;
 wire \u_cpu.ALU._0739_ ;
 wire \u_cpu.ALU._0740_ ;
 wire \u_cpu.ALU._0741_ ;
 wire \u_cpu.ALU._0742_ ;
 wire \u_cpu.ALU._0743_ ;
 wire \u_cpu.ALU._0744_ ;
 wire \u_cpu.ALU._0745_ ;
 wire \u_cpu.ALU._0746_ ;
 wire \u_cpu.ALU._0747_ ;
 wire \u_cpu.ALU._0748_ ;
 wire \u_cpu.ALU._0749_ ;
 wire \u_cpu.ALU._0750_ ;
 wire \u_cpu.ALU._0751_ ;
 wire \u_cpu.ALU._0752_ ;
 wire \u_cpu.ALU._0753_ ;
 wire \u_cpu.ALU._0754_ ;
 wire \u_cpu.ALU._0755_ ;
 wire \u_cpu.ALU._0756_ ;
 wire \u_cpu.ALU._0757_ ;
 wire \u_cpu.ALU._0758_ ;
 wire \u_cpu.ALU._0759_ ;
 wire \u_cpu.ALU._0760_ ;
 wire \u_cpu.ALU._0761_ ;
 wire \u_cpu.ALU._0762_ ;
 wire \u_cpu.ALU._0763_ ;
 wire \u_cpu.ALU._0764_ ;
 wire \u_cpu.ALU._0765_ ;
 wire \u_cpu.ALU._0766_ ;
 wire \u_cpu.ALU._0767_ ;
 wire \u_cpu.ALU._0768_ ;
 wire \u_cpu.ALU._0769_ ;
 wire \u_cpu.ALU._0770_ ;
 wire \u_cpu.ALU._0771_ ;
 wire \u_cpu.ALU._0772_ ;
 wire \u_cpu.ALU._0773_ ;
 wire \u_cpu.ALU._0774_ ;
 wire \u_cpu.ALU._0775_ ;
 wire \u_cpu.ALU._0776_ ;
 wire \u_cpu.ALU._0777_ ;
 wire \u_cpu.ALU._0778_ ;
 wire \u_cpu.ALU._0779_ ;
 wire \u_cpu.ALU._0780_ ;
 wire \u_cpu.ALU._0781_ ;
 wire \u_cpu.ALU._0782_ ;
 wire \u_cpu.ALU._0783_ ;
 wire \u_cpu.ALU._0784_ ;
 wire \u_cpu.ALU._0785_ ;
 wire \u_cpu.ALU._0786_ ;
 wire \u_cpu.ALU._0787_ ;
 wire \u_cpu.ALU._0788_ ;
 wire \u_cpu.ALU._0789_ ;
 wire \u_cpu.ALU._0790_ ;
 wire \u_cpu.ALU._0791_ ;
 wire \u_cpu.ALU._0792_ ;
 wire \u_cpu.ALU._0793_ ;
 wire \u_cpu.ALU._0794_ ;
 wire \u_cpu.ALU._0795_ ;
 wire \u_cpu.ALU._0796_ ;
 wire \u_cpu.ALU._0797_ ;
 wire \u_cpu.ALU._0798_ ;
 wire \u_cpu.ALU._0799_ ;
 wire \u_cpu.ALU._0800_ ;
 wire \u_cpu.ALU._0801_ ;
 wire \u_cpu.ALU._0802_ ;
 wire \u_cpu.ALU._0803_ ;
 wire \u_cpu.ALU._0804_ ;
 wire \u_cpu.ALU._0805_ ;
 wire \u_cpu.ALU._0806_ ;
 wire \u_cpu.ALU._0807_ ;
 wire \u_cpu.ALU._0808_ ;
 wire \u_cpu.ALU._0809_ ;
 wire \u_cpu.ALU._0810_ ;
 wire \u_cpu.ALU._0811_ ;
 wire \u_cpu.ALU._0812_ ;
 wire \u_cpu.ALU._0813_ ;
 wire \u_cpu.ALU._0814_ ;
 wire \u_cpu.ALU._0815_ ;
 wire \u_cpu.ALU._0816_ ;
 wire \u_cpu.ALU._0817_ ;
 wire \u_cpu.ALU._0818_ ;
 wire \u_cpu.ALU._0819_ ;
 wire \u_cpu.ALU._0820_ ;
 wire \u_cpu.ALU._0821_ ;
 wire \u_cpu.ALU._0822_ ;
 wire \u_cpu.ALU._0823_ ;
 wire \u_cpu.ALU._0824_ ;
 wire \u_cpu.ALU._0825_ ;
 wire \u_cpu.ALU._0826_ ;
 wire \u_cpu.ALU._0827_ ;
 wire \u_cpu.ALU._0828_ ;
 wire \u_cpu.ALU._0829_ ;
 wire \u_cpu.ALU._0830_ ;
 wire \u_cpu.ALU._0831_ ;
 wire \u_cpu.ALU._0832_ ;
 wire \u_cpu.ALU._0833_ ;
 wire \u_cpu.ALU._0834_ ;
 wire \u_cpu.ALU._0835_ ;
 wire \u_cpu.ALU._0836_ ;
 wire \u_cpu.ALU._0837_ ;
 wire \u_cpu.ALU._0838_ ;
 wire \u_cpu.ALU._0839_ ;
 wire \u_cpu.ALU._0840_ ;
 wire \u_cpu.ALU._0841_ ;
 wire \u_cpu.ALU._0842_ ;
 wire \u_cpu.ALU._0843_ ;
 wire \u_cpu.ALU._0844_ ;
 wire \u_cpu.ALU._0845_ ;
 wire \u_cpu.ALU._0846_ ;
 wire \u_cpu.ALU._0847_ ;
 wire \u_cpu.ALU._0848_ ;
 wire \u_cpu.ALU._0849_ ;
 wire \u_cpu.ALU._0850_ ;
 wire \u_cpu.ALU._0851_ ;
 wire \u_cpu.ALU._0852_ ;
 wire \u_cpu.ALU._0853_ ;
 wire \u_cpu.ALU._0854_ ;
 wire \u_cpu.ALU._0855_ ;
 wire \u_cpu.ALU._0856_ ;
 wire \u_cpu.ALU._0857_ ;
 wire \u_cpu.ALU._0858_ ;
 wire \u_cpu.ALU._0859_ ;
 wire \u_cpu.ALU._0860_ ;
 wire \u_cpu.ALU._0861_ ;
 wire \u_cpu.ALU._0862_ ;
 wire \u_cpu.ALU._0863_ ;
 wire \u_cpu.ALU._0864_ ;
 wire \u_cpu.ALU._0865_ ;
 wire \u_cpu.ALU._0866_ ;
 wire \u_cpu.ALU._0867_ ;
 wire \u_cpu.ALU._0868_ ;
 wire \u_cpu.ALU._0869_ ;
 wire \u_cpu.ALU._0870_ ;
 wire \u_cpu.ALU._0871_ ;
 wire \u_cpu.ALU._0872_ ;
 wire \u_cpu.ALU._0873_ ;
 wire \u_cpu.ALU._0874_ ;
 wire \u_cpu.ALU._0875_ ;
 wire \u_cpu.ALU._0876_ ;
 wire \u_cpu.ALU._0877_ ;
 wire \u_cpu.ALU._0878_ ;
 wire \u_cpu.ALU._0879_ ;
 wire \u_cpu.ALU._0880_ ;
 wire \u_cpu.ALU._0881_ ;
 wire \u_cpu.ALU._0882_ ;
 wire \u_cpu.ALU._0883_ ;
 wire \u_cpu.ALU._0884_ ;
 wire \u_cpu.ALU._0885_ ;
 wire \u_cpu.ALU._0886_ ;
 wire \u_cpu.ALU._0887_ ;
 wire \u_cpu.ALU._0888_ ;
 wire \u_cpu.ALU._0889_ ;
 wire \u_cpu.ALU._0890_ ;
 wire \u_cpu.ALU._0891_ ;
 wire \u_cpu.ALU._0892_ ;
 wire \u_cpu.ALU._0893_ ;
 wire \u_cpu.ALU._0894_ ;
 wire \u_cpu.ALU._0895_ ;
 wire \u_cpu.ALU._0896_ ;
 wire \u_cpu.ALU._0897_ ;
 wire \u_cpu.ALU._0898_ ;
 wire \u_cpu.ALU._0899_ ;
 wire \u_cpu.ALU._0900_ ;
 wire \u_cpu.ALU._0901_ ;
 wire \u_cpu.ALU._0902_ ;
 wire \u_cpu.ALU._0903_ ;
 wire \u_cpu.ALU._0904_ ;
 wire \u_cpu.ALU._0905_ ;
 wire \u_cpu.ALU._0906_ ;
 wire \u_cpu.ALU._0907_ ;
 wire \u_cpu.ALU._0908_ ;
 wire \u_cpu.ALU._0909_ ;
 wire \u_cpu.ALU._0910_ ;
 wire \u_cpu.ALU._0911_ ;
 wire \u_cpu.ALU._0912_ ;
 wire \u_cpu.ALU._0913_ ;
 wire \u_cpu.ALU._0914_ ;
 wire \u_cpu.ALU._0915_ ;
 wire \u_cpu.ALU._0916_ ;
 wire \u_cpu.ALU._0917_ ;
 wire \u_cpu.ALU._0918_ ;
 wire \u_cpu.ALU._0919_ ;
 wire \u_cpu.ALU._0920_ ;
 wire \u_cpu.ALU._0921_ ;
 wire \u_cpu.ALU._0922_ ;
 wire \u_cpu.ALU._0923_ ;
 wire \u_cpu.ALU._0924_ ;
 wire \u_cpu.ALU._0925_ ;
 wire \u_cpu.ALU._0926_ ;
 wire \u_cpu.ALU._0927_ ;
 wire \u_cpu.ALU._0928_ ;
 wire \u_cpu.ALU._0929_ ;
 wire \u_cpu.ALU._0930_ ;
 wire \u_cpu.ALU._0931_ ;
 wire \u_cpu.ALU._0932_ ;
 wire \u_cpu.ALU._0933_ ;
 wire \u_cpu.ALU._0934_ ;
 wire \u_cpu.ALU._0935_ ;
 wire \u_cpu.ALU._0936_ ;
 wire \u_cpu.ALU._0937_ ;
 wire \u_cpu.ALU._0938_ ;
 wire \u_cpu.ALU._0939_ ;
 wire \u_cpu.ALU._0940_ ;
 wire \u_cpu.ALU._0941_ ;
 wire \u_cpu.ALU._0942_ ;
 wire \u_cpu.ALU._0943_ ;
 wire \u_cpu.ALU._0944_ ;
 wire \u_cpu.ALU._0945_ ;
 wire \u_cpu.ALU._0946_ ;
 wire \u_cpu.ALU._0947_ ;
 wire \u_cpu.ALU._0948_ ;
 wire \u_cpu.ALU._0949_ ;
 wire \u_cpu.ALU._0950_ ;
 wire \u_cpu.ALU._0951_ ;
 wire \u_cpu.ALU._0952_ ;
 wire \u_cpu.ALU._0953_ ;
 wire \u_cpu.ALU._0954_ ;
 wire \u_cpu.ALU._0955_ ;
 wire \u_cpu.ALU._0956_ ;
 wire \u_cpu.ALU._0957_ ;
 wire \u_cpu.ALU._0958_ ;
 wire \u_cpu.ALU._0959_ ;
 wire \u_cpu.ALU._0960_ ;
 wire \u_cpu.ALU._0961_ ;
 wire \u_cpu.ALU._0962_ ;
 wire \u_cpu.ALU._0963_ ;
 wire \u_cpu.ALU._0964_ ;
 wire \u_cpu.ALU._0965_ ;
 wire \u_cpu.ALU._0966_ ;
 wire \u_cpu.ALU._0967_ ;
 wire \u_cpu.ALU._0968_ ;
 wire \u_cpu.ALU._0969_ ;
 wire \u_cpu.ALU._0970_ ;
 wire \u_cpu.ALU._0971_ ;
 wire \u_cpu.ALU._0972_ ;
 wire \u_cpu.ALU._0973_ ;
 wire \u_cpu.ALU._0974_ ;
 wire \u_cpu.ALU._0975_ ;
 wire \u_cpu.ALU._0976_ ;
 wire \u_cpu.ALU._0977_ ;
 wire \u_cpu.ALU._0978_ ;
 wire \u_cpu.ALU._0979_ ;
 wire \u_cpu.ALU._0980_ ;
 wire \u_cpu.ALU._0981_ ;
 wire \u_cpu.ALU._0982_ ;
 wire \u_cpu.ALU._0983_ ;
 wire \u_cpu.ALU._0984_ ;
 wire \u_cpu.ALU._0985_ ;
 wire \u_cpu.ALU._0986_ ;
 wire \u_cpu.ALU._0987_ ;
 wire \u_cpu.ALU._0988_ ;
 wire \u_cpu.ALU._0989_ ;
 wire \u_cpu.ALU._0990_ ;
 wire \u_cpu.ALU._0991_ ;
 wire \u_cpu.ALU._0992_ ;
 wire \u_cpu.ALU._0993_ ;
 wire \u_cpu.ALU._0994_ ;
 wire \u_cpu.ALU._0995_ ;
 wire \u_cpu.ALU._0996_ ;
 wire \u_cpu.ALU._0997_ ;
 wire \u_cpu.ALU._0998_ ;
 wire \u_cpu.ALU._0999_ ;
 wire \u_cpu.ALU._1000_ ;
 wire \u_cpu.ALU._1001_ ;
 wire \u_cpu.ALU._1002_ ;
 wire \u_cpu.ALU._1003_ ;
 wire \u_cpu.ALU._1004_ ;
 wire \u_cpu.ALU._1005_ ;
 wire \u_cpu.ALU._1006_ ;
 wire \u_cpu.ALU._1007_ ;
 wire \u_cpu.ALU._1008_ ;
 wire \u_cpu.ALU._1009_ ;
 wire \u_cpu.ALU._1010_ ;
 wire \u_cpu.ALU._1011_ ;
 wire \u_cpu.ALU._1012_ ;
 wire \u_cpu.ALU._1013_ ;
 wire \u_cpu.ALU._1014_ ;
 wire \u_cpu.ALU._1015_ ;
 wire \u_cpu.ALU._1016_ ;
 wire \u_cpu.ALU._1017_ ;
 wire \u_cpu.ALU._1018_ ;
 wire \u_cpu.ALU._1019_ ;
 wire \u_cpu.ALU._1020_ ;
 wire \u_cpu.ALU._1021_ ;
 wire \u_cpu.ALU._1022_ ;
 wire \u_cpu.ALU._1023_ ;
 wire \u_cpu.ALU._1024_ ;
 wire \u_cpu.ALU._1025_ ;
 wire \u_cpu.ALU._1026_ ;
 wire \u_cpu.ALU._1027_ ;
 wire \u_cpu.ALU._1028_ ;
 wire \u_cpu.ALU._1029_ ;
 wire \u_cpu.ALU._1030_ ;
 wire \u_cpu.ALU._1031_ ;
 wire \u_cpu.ALU._1032_ ;
 wire \u_cpu.ALU._1033_ ;
 wire \u_cpu.ALU._1034_ ;
 wire \u_cpu.ALU._1035_ ;
 wire \u_cpu.ALU._1036_ ;
 wire \u_cpu.ALU._1037_ ;
 wire \u_cpu.ALU._1038_ ;
 wire \u_cpu.ALU._1039_ ;
 wire \u_cpu.ALU._1040_ ;
 wire \u_cpu.ALU._1041_ ;
 wire \u_cpu.ALU._1042_ ;
 wire \u_cpu.ALU._1043_ ;
 wire \u_cpu.ALU._1044_ ;
 wire \u_cpu.ALU._1045_ ;
 wire \u_cpu.ALU._1046_ ;
 wire \u_cpu.ALU._1047_ ;
 wire \u_cpu.ALU._1048_ ;
 wire \u_cpu.ALU._1049_ ;
 wire \u_cpu.ALU._1050_ ;
 wire \u_cpu.ALU._1051_ ;
 wire \u_cpu.ALU._1052_ ;
 wire \u_cpu.ALU._1053_ ;
 wire \u_cpu.ALU._1054_ ;
 wire \u_cpu.ALU._1055_ ;
 wire \u_cpu.ALU._1056_ ;
 wire \u_cpu.ALU._1057_ ;
 wire \u_cpu.ALU._1058_ ;
 wire \u_cpu.ALU._1059_ ;
 wire \u_cpu.ALU._1060_ ;
 wire \u_cpu.ALU._1061_ ;
 wire \u_cpu.ALU._1062_ ;
 wire \u_cpu.ALU._1063_ ;
 wire \u_cpu.ALU._1064_ ;
 wire \u_cpu.ALU._1065_ ;
 wire \u_cpu.ALU._1066_ ;
 wire \u_cpu.ALU._1067_ ;
 wire \u_cpu.ALU._1068_ ;
 wire \u_cpu.ALU._1069_ ;
 wire \u_cpu.ALU._1070_ ;
 wire \u_cpu.ALU._1071_ ;
 wire \u_cpu.ALU._1072_ ;
 wire \u_cpu.ALU._1073_ ;
 wire \u_cpu.ALU._1074_ ;
 wire \u_cpu.ALU._1075_ ;
 wire \u_cpu.ALU._1076_ ;
 wire \u_cpu.ALU._1077_ ;
 wire \u_cpu.ALU._1078_ ;
 wire \u_cpu.ALU._1079_ ;
 wire \u_cpu.ALU._1080_ ;
 wire \u_cpu.ALU._1081_ ;
 wire \u_cpu.ALU._1082_ ;
 wire \u_cpu.ALU._1083_ ;
 wire \u_cpu.ALU._1084_ ;
 wire \u_cpu.ALU._1085_ ;
 wire \u_cpu.ALU._1086_ ;
 wire \u_cpu.ALU._1087_ ;
 wire \u_cpu.ALU._1088_ ;
 wire \u_cpu.ALU._1089_ ;
 wire \u_cpu.ALU._1090_ ;
 wire \u_cpu.ALU._1091_ ;
 wire \u_cpu.ALU._1092_ ;
 wire \u_cpu.ALU._1093_ ;
 wire \u_cpu.ALU._1094_ ;
 wire \u_cpu.ALU._1095_ ;
 wire \u_cpu.ALU._1096_ ;
 wire \u_cpu.ALU._1097_ ;
 wire \u_cpu.ALU._1098_ ;
 wire \u_cpu.ALU._1099_ ;
 wire \u_cpu.ALU._1100_ ;
 wire \u_cpu.ALU._1101_ ;
 wire \u_cpu.ALU._1102_ ;
 wire \u_cpu.ALU._1103_ ;
 wire \u_cpu.ALU._1104_ ;
 wire \u_cpu.ALU._1105_ ;
 wire \u_cpu.ALU._1106_ ;
 wire \u_cpu.ALU._1107_ ;
 wire \u_cpu.ALU._1108_ ;
 wire \u_cpu.ALU._1109_ ;
 wire \u_cpu.ALU._1110_ ;
 wire \u_cpu.ALU._1111_ ;
 wire \u_cpu.ALU._1112_ ;
 wire \u_cpu.ALU._1113_ ;
 wire \u_cpu.ALU._1114_ ;
 wire \u_cpu.ALU._1115_ ;
 wire \u_cpu.ALU._1116_ ;
 wire \u_cpu.ALU._1117_ ;
 wire \u_cpu.ALU._1118_ ;
 wire \u_cpu.ALU._1119_ ;
 wire \u_cpu.ALU._1120_ ;
 wire \u_cpu.ALU._1121_ ;
 wire \u_cpu.ALU._1122_ ;
 wire \u_cpu.ALU._1123_ ;
 wire \u_cpu.ALU._1124_ ;
 wire \u_cpu.ALU._1125_ ;
 wire \u_cpu.ALU._1126_ ;
 wire \u_cpu.ALU._1127_ ;
 wire \u_cpu.ALU._1128_ ;
 wire \u_cpu.ALU._1129_ ;
 wire \u_cpu.ALU._1130_ ;
 wire \u_cpu.ALU._1131_ ;
 wire \u_cpu.ALU._1132_ ;
 wire \u_cpu.ALU._1133_ ;
 wire \u_cpu.ALU._1134_ ;
 wire \u_cpu.ALU._1135_ ;
 wire \u_cpu.ALU._1136_ ;
 wire \u_cpu.ALU._1137_ ;
 wire \u_cpu.ALU._1138_ ;
 wire \u_cpu.ALU._1139_ ;
 wire \u_cpu.ALU._1140_ ;
 wire \u_cpu.ALU._1141_ ;
 wire \u_cpu.ALU._1142_ ;
 wire \u_cpu.ALU._1143_ ;
 wire \u_cpu.ALU._1144_ ;
 wire \u_cpu.ALU._1145_ ;
 wire \u_cpu.ALU._1146_ ;
 wire \u_cpu.ALU._1147_ ;
 wire \u_cpu.ALU._1148_ ;
 wire \u_cpu.ALU._1149_ ;
 wire \u_cpu.ALU._1150_ ;
 wire \u_cpu.ALU._1151_ ;
 wire \u_cpu.ALU._1152_ ;
 wire \u_cpu.ALU._1153_ ;
 wire \u_cpu.ALU._1154_ ;
 wire \u_cpu.ALU._1155_ ;
 wire \u_cpu.ALU._1156_ ;
 wire \u_cpu.ALU._1157_ ;
 wire \u_cpu.ALU._1158_ ;
 wire \u_cpu.ALU._1159_ ;
 wire \u_cpu.ALU._1160_ ;
 wire \u_cpu.ALU._1161_ ;
 wire \u_cpu.ALU._1162_ ;
 wire \u_cpu.ALU._1163_ ;
 wire \u_cpu.ALU._1164_ ;
 wire \u_cpu.ALU._1165_ ;
 wire \u_cpu.ALU._1166_ ;
 wire \u_cpu.ALU._1167_ ;
 wire \u_cpu.ALU._1168_ ;
 wire \u_cpu.ALU._1169_ ;
 wire \u_cpu.ALU._1170_ ;
 wire \u_cpu.ALU._1171_ ;
 wire \u_cpu.ALU._1172_ ;
 wire \u_cpu.ALU._1173_ ;
 wire \u_cpu.ALU._1174_ ;
 wire \u_cpu.ALU._1175_ ;
 wire \u_cpu.ALU._1176_ ;
 wire \u_cpu.ALU._1177_ ;
 wire \u_cpu.ALU._1178_ ;
 wire \u_cpu.ALU._1179_ ;
 wire \u_cpu.ALU._1180_ ;
 wire \u_cpu.ALU._1181_ ;
 wire \u_cpu.ALU._1182_ ;
 wire \u_cpu.ALU._1183_ ;
 wire \u_cpu.ALU._1184_ ;
 wire \u_cpu.ALU._1185_ ;
 wire \u_cpu.ALU._1186_ ;
 wire \u_cpu.ALU._1187_ ;
 wire \u_cpu.ALU._1188_ ;
 wire \u_cpu.ALU._1189_ ;
 wire \u_cpu.ALU._1190_ ;
 wire \u_cpu.ALU._1191_ ;
 wire \u_cpu.ALU._1192_ ;
 wire \u_cpu.ALU._1193_ ;
 wire \u_cpu.ALU._1194_ ;
 wire \u_cpu.ALU._1195_ ;
 wire \u_cpu.ALU._1196_ ;
 wire \u_cpu.ALU._1197_ ;
 wire \u_cpu.ALU._1198_ ;
 wire \u_cpu.ALU._1199_ ;
 wire \u_cpu.ALU._1200_ ;
 wire \u_cpu.ALU._1201_ ;
 wire \u_cpu.ALU._1202_ ;
 wire \u_cpu.ALU._1203_ ;
 wire \u_cpu.ALU._1204_ ;
 wire \u_cpu.ALU._1205_ ;
 wire \u_cpu.ALU._1206_ ;
 wire \u_cpu.ALU._1207_ ;
 wire \u_cpu.ALU._1208_ ;
 wire \u_cpu.ALU._1209_ ;
 wire \u_cpu.ALU._1210_ ;
 wire \u_cpu.ALU._1211_ ;
 wire \u_cpu.ALU._1212_ ;
 wire \u_cpu.ALU._1213_ ;
 wire \u_cpu.ALU._1214_ ;
 wire \u_cpu.ALU._1215_ ;
 wire \u_cpu.ALU._1216_ ;
 wire \u_cpu.ALU._1217_ ;
 wire \u_cpu.ALU._1218_ ;
 wire \u_cpu.ALU._1219_ ;
 wire \u_cpu.ALU._1220_ ;
 wire \u_cpu.ALU._1221_ ;
 wire \u_cpu.ALU._1222_ ;
 wire \u_cpu.ALU._1223_ ;
 wire \u_cpu.ALU._1224_ ;
 wire \u_cpu.ALU._1225_ ;
 wire \u_cpu.ALU._1226_ ;
 wire \u_cpu.ALU._1227_ ;
 wire \u_cpu.ALU._1228_ ;
 wire \u_cpu.ALU._1229_ ;
 wire \u_cpu.ALU._1230_ ;
 wire \u_cpu.ALU._1231_ ;
 wire \u_cpu.ALU._1232_ ;
 wire \u_cpu.ALU._1233_ ;
 wire \u_cpu.ALU._1234_ ;
 wire \u_cpu.ALU._1235_ ;
 wire \u_cpu.ALU._1236_ ;
 wire \u_cpu.ALU._1237_ ;
 wire \u_cpu.ALU._1238_ ;
 wire \u_cpu.ALU._1239_ ;
 wire \u_cpu.ALU._1240_ ;
 wire \u_cpu.ALU._1241_ ;
 wire \u_cpu.ALU._1242_ ;
 wire \u_cpu.ALU._1243_ ;
 wire \u_cpu.ALU._1244_ ;
 wire \u_cpu.ALU._1245_ ;
 wire \u_cpu.ALU._1246_ ;
 wire \u_cpu.ALU._1247_ ;
 wire \u_cpu.ALU._1248_ ;
 wire \u_cpu.ALU._1249_ ;
 wire \u_cpu.ALU._1250_ ;
 wire \u_cpu.ALU._1251_ ;
 wire \u_cpu.ALU._1252_ ;
 wire \u_cpu.ALU._1253_ ;
 wire \u_cpu.ALU._1254_ ;
 wire \u_cpu.ALU._1255_ ;
 wire \u_cpu.ALU._1256_ ;
 wire \u_cpu.ALU._1257_ ;
 wire \u_cpu.ALU._1258_ ;
 wire \u_cpu.ALU._1259_ ;
 wire \u_cpu.ALU._1260_ ;
 wire \u_cpu.ALU._1261_ ;
 wire \u_cpu.ALU._1262_ ;
 wire \u_cpu.ALU._1263_ ;
 wire \u_cpu.ALU._1264_ ;
 wire \u_cpu.ALU._1265_ ;
 wire \u_cpu.ALU._1266_ ;
 wire \u_cpu.ALU._1267_ ;
 wire \u_cpu.ALU._1268_ ;
 wire \u_cpu.ALU._1269_ ;
 wire \u_cpu.ALU._1270_ ;
 wire \u_cpu.ALU._1271_ ;
 wire \u_cpu.ALU._1272_ ;
 wire \u_cpu.ALU._1273_ ;
 wire \u_cpu.ALU._1274_ ;
 wire \u_cpu.ALU._1275_ ;
 wire \u_cpu.ALU._1276_ ;
 wire \u_cpu.ALU._1277_ ;
 wire \u_cpu.ALU._1278_ ;
 wire \u_cpu.ALU._1279_ ;
 wire \u_cpu.ALU._1280_ ;
 wire \u_cpu.ALU._1281_ ;
 wire \u_cpu.ALU._1282_ ;
 wire \u_cpu.ALU._1283_ ;
 wire \u_cpu.ALU._1284_ ;
 wire \u_cpu.ALU._1285_ ;
 wire \u_cpu.ALU._1286_ ;
 wire \u_cpu.ALU._1287_ ;
 wire \u_cpu.ALU._1288_ ;
 wire \u_cpu.ALU._1289_ ;
 wire \u_cpu.ALU._1290_ ;
 wire \u_cpu.ALU._1291_ ;
 wire \u_cpu.ALU._1292_ ;
 wire \u_cpu.ALU._1293_ ;
 wire \u_cpu.ALU._1294_ ;
 wire \u_cpu.ALU._1295_ ;
 wire \u_cpu.ALU._1296_ ;
 wire \u_cpu.ALU._1297_ ;
 wire \u_cpu.ALU._1298_ ;
 wire \u_cpu.ALU._1299_ ;
 wire \u_cpu.ALU._1300_ ;
 wire \u_cpu.ALU._1301_ ;
 wire \u_cpu.ALU._1302_ ;
 wire \u_cpu.ALU._1303_ ;
 wire \u_cpu.ALU._1304_ ;
 wire \u_cpu.ALU._1305_ ;
 wire \u_cpu.ALU._1306_ ;
 wire \u_cpu.ALU._1307_ ;
 wire \u_cpu.ALU._1308_ ;
 wire \u_cpu.ALU._1309_ ;
 wire \u_cpu.ALU._1310_ ;
 wire \u_cpu.ALU._1311_ ;
 wire \u_cpu.ALU._1312_ ;
 wire \u_cpu.ALU._1313_ ;
 wire \u_cpu.ALU._1314_ ;
 wire \u_cpu.ALU._1315_ ;
 wire \u_cpu.ALU._1316_ ;
 wire \u_cpu.ALU._1317_ ;
 wire \u_cpu.ALU._1318_ ;
 wire \u_cpu.ALU._1319_ ;
 wire \u_cpu.ALU._1320_ ;
 wire \u_cpu.ALU._1321_ ;
 wire \u_cpu.ALU._1322_ ;
 wire \u_cpu.ALU._1323_ ;
 wire \u_cpu.ALU._1324_ ;
 wire \u_cpu.ALU._1325_ ;
 wire \u_cpu.ALU._1326_ ;
 wire \u_cpu.ALU._1327_ ;
 wire \u_cpu.ALU._1328_ ;
 wire \u_cpu.ALU._1329_ ;
 wire \u_cpu.ALU._1330_ ;
 wire \u_cpu.ALU._1331_ ;
 wire \u_cpu.ALU._1332_ ;
 wire \u_cpu.ALU._1333_ ;
 wire \u_cpu.ALU._1334_ ;
 wire \u_cpu.ALU._1335_ ;
 wire \u_cpu.ALU._1336_ ;
 wire \u_cpu.ALU._1337_ ;
 wire \u_cpu.ALU._1338_ ;
 wire \u_cpu.ALU._1339_ ;
 wire \u_cpu.ALU._1340_ ;
 wire \u_cpu.ALU._1341_ ;
 wire \u_cpu.ALU._1342_ ;
 wire \u_cpu.ALU._1343_ ;
 wire \u_cpu.ALU._1344_ ;
 wire \u_cpu.ALU._1345_ ;
 wire \u_cpu.ALU._1346_ ;
 wire \u_cpu.ALU._1347_ ;
 wire \u_cpu.ALU._1348_ ;
 wire \u_cpu.ALU._1349_ ;
 wire \u_cpu.ALU._1350_ ;
 wire \u_cpu.ALU.u_wallace._0000_ ;
 wire \u_cpu.ALU.u_wallace._0001_ ;
 wire \u_cpu.ALU.u_wallace._0002_ ;
 wire \u_cpu.ALU.u_wallace._0003_ ;
 wire \u_cpu.ALU.u_wallace._0004_ ;
 wire \u_cpu.ALU.u_wallace._0005_ ;
 wire \u_cpu.ALU.u_wallace._0006_ ;
 wire \u_cpu.ALU.u_wallace._0007_ ;
 wire \u_cpu.ALU.u_wallace._0008_ ;
 wire \u_cpu.ALU.u_wallace._0009_ ;
 wire \u_cpu.ALU.u_wallace._0010_ ;
 wire \u_cpu.ALU.u_wallace._0011_ ;
 wire \u_cpu.ALU.u_wallace._0012_ ;
 wire \u_cpu.ALU.u_wallace._0013_ ;
 wire \u_cpu.ALU.u_wallace._0014_ ;
 wire \u_cpu.ALU.u_wallace._0015_ ;
 wire \u_cpu.ALU.u_wallace._0016_ ;
 wire \u_cpu.ALU.u_wallace._0017_ ;
 wire \u_cpu.ALU.u_wallace._0018_ ;
 wire \u_cpu.ALU.u_wallace._0019_ ;
 wire \u_cpu.ALU.u_wallace._0020_ ;
 wire \u_cpu.ALU.u_wallace._0021_ ;
 wire \u_cpu.ALU.u_wallace._0022_ ;
 wire \u_cpu.ALU.u_wallace._0023_ ;
 wire \u_cpu.ALU.u_wallace._0024_ ;
 wire \u_cpu.ALU.u_wallace._0025_ ;
 wire \u_cpu.ALU.u_wallace._0026_ ;
 wire \u_cpu.ALU.u_wallace._0027_ ;
 wire \u_cpu.ALU.u_wallace._0028_ ;
 wire \u_cpu.ALU.u_wallace._0029_ ;
 wire \u_cpu.ALU.u_wallace._0030_ ;
 wire \u_cpu.ALU.u_wallace._0031_ ;
 wire \u_cpu.ALU.u_wallace._0032_ ;
 wire \u_cpu.ALU.u_wallace._0033_ ;
 wire \u_cpu.ALU.u_wallace._0034_ ;
 wire \u_cpu.ALU.u_wallace._0035_ ;
 wire \u_cpu.ALU.u_wallace._0036_ ;
 wire \u_cpu.ALU.u_wallace._0037_ ;
 wire \u_cpu.ALU.u_wallace._0038_ ;
 wire \u_cpu.ALU.u_wallace._0039_ ;
 wire \u_cpu.ALU.u_wallace._0040_ ;
 wire \u_cpu.ALU.u_wallace._0041_ ;
 wire \u_cpu.ALU.u_wallace._0042_ ;
 wire \u_cpu.ALU.u_wallace._0043_ ;
 wire \u_cpu.ALU.u_wallace._0044_ ;
 wire \u_cpu.ALU.u_wallace._0045_ ;
 wire \u_cpu.ALU.u_wallace._0046_ ;
 wire \u_cpu.ALU.u_wallace._0047_ ;
 wire \u_cpu.ALU.u_wallace._0048_ ;
 wire \u_cpu.ALU.u_wallace._0049_ ;
 wire \u_cpu.ALU.u_wallace._0050_ ;
 wire \u_cpu.ALU.u_wallace._0051_ ;
 wire \u_cpu.ALU.u_wallace._0052_ ;
 wire \u_cpu.ALU.u_wallace._0053_ ;
 wire \u_cpu.ALU.u_wallace._0054_ ;
 wire \u_cpu.ALU.u_wallace._0055_ ;
 wire \u_cpu.ALU.u_wallace._0056_ ;
 wire \u_cpu.ALU.u_wallace._0057_ ;
 wire \u_cpu.ALU.u_wallace._0058_ ;
 wire \u_cpu.ALU.u_wallace._0059_ ;
 wire \u_cpu.ALU.u_wallace._0060_ ;
 wire \u_cpu.ALU.u_wallace._0061_ ;
 wire \u_cpu.ALU.u_wallace._0062_ ;
 wire \u_cpu.ALU.u_wallace._0063_ ;
 wire \u_cpu.ALU.u_wallace._0064_ ;
 wire \u_cpu.ALU.u_wallace._0065_ ;
 wire \u_cpu.ALU.u_wallace._0066_ ;
 wire \u_cpu.ALU.u_wallace._0067_ ;
 wire \u_cpu.ALU.u_wallace._0068_ ;
 wire \u_cpu.ALU.u_wallace._0069_ ;
 wire \u_cpu.ALU.u_wallace._0070_ ;
 wire \u_cpu.ALU.u_wallace._0071_ ;
 wire \u_cpu.ALU.u_wallace._0072_ ;
 wire \u_cpu.ALU.u_wallace._0073_ ;
 wire \u_cpu.ALU.u_wallace._0074_ ;
 wire \u_cpu.ALU.u_wallace._0075_ ;
 wire \u_cpu.ALU.u_wallace._0076_ ;
 wire \u_cpu.ALU.u_wallace._0077_ ;
 wire \u_cpu.ALU.u_wallace._0078_ ;
 wire \u_cpu.ALU.u_wallace._0079_ ;
 wire \u_cpu.ALU.u_wallace._0080_ ;
 wire \u_cpu.ALU.u_wallace._0081_ ;
 wire \u_cpu.ALU.u_wallace._0082_ ;
 wire \u_cpu.ALU.u_wallace._0083_ ;
 wire \u_cpu.ALU.u_wallace._0084_ ;
 wire \u_cpu.ALU.u_wallace._0085_ ;
 wire \u_cpu.ALU.u_wallace._0086_ ;
 wire \u_cpu.ALU.u_wallace._0087_ ;
 wire \u_cpu.ALU.u_wallace._0088_ ;
 wire \u_cpu.ALU.u_wallace._0089_ ;
 wire \u_cpu.ALU.u_wallace._0090_ ;
 wire \u_cpu.ALU.u_wallace._0091_ ;
 wire \u_cpu.ALU.u_wallace._0092_ ;
 wire \u_cpu.ALU.u_wallace._0093_ ;
 wire \u_cpu.ALU.u_wallace._0094_ ;
 wire \u_cpu.ALU.u_wallace._0095_ ;
 wire \u_cpu.ALU.u_wallace._0096_ ;
 wire \u_cpu.ALU.u_wallace._0097_ ;
 wire \u_cpu.ALU.u_wallace._0098_ ;
 wire \u_cpu.ALU.u_wallace._0099_ ;
 wire \u_cpu.ALU.u_wallace._0100_ ;
 wire \u_cpu.ALU.u_wallace._0101_ ;
 wire \u_cpu.ALU.u_wallace._0102_ ;
 wire \u_cpu.ALU.u_wallace._0103_ ;
 wire \u_cpu.ALU.u_wallace._0104_ ;
 wire \u_cpu.ALU.u_wallace._0105_ ;
 wire \u_cpu.ALU.u_wallace._0106_ ;
 wire \u_cpu.ALU.u_wallace._0107_ ;
 wire \u_cpu.ALU.u_wallace._0108_ ;
 wire \u_cpu.ALU.u_wallace._0109_ ;
 wire \u_cpu.ALU.u_wallace._0110_ ;
 wire \u_cpu.ALU.u_wallace._0111_ ;
 wire \u_cpu.ALU.u_wallace._0112_ ;
 wire \u_cpu.ALU.u_wallace._0113_ ;
 wire \u_cpu.ALU.u_wallace._0114_ ;
 wire \u_cpu.ALU.u_wallace._0115_ ;
 wire \u_cpu.ALU.u_wallace._0116_ ;
 wire \u_cpu.ALU.u_wallace._0117_ ;
 wire \u_cpu.ALU.u_wallace._0118_ ;
 wire \u_cpu.ALU.u_wallace._0119_ ;
 wire \u_cpu.ALU.u_wallace._0120_ ;
 wire \u_cpu.ALU.u_wallace._0121_ ;
 wire \u_cpu.ALU.u_wallace._0122_ ;
 wire \u_cpu.ALU.u_wallace._0123_ ;
 wire \u_cpu.ALU.u_wallace._0124_ ;
 wire \u_cpu.ALU.u_wallace._0125_ ;
 wire \u_cpu.ALU.u_wallace._0126_ ;
 wire \u_cpu.ALU.u_wallace._0127_ ;
 wire \u_cpu.ALU.u_wallace._0128_ ;
 wire \u_cpu.ALU.u_wallace._0129_ ;
 wire \u_cpu.ALU.u_wallace._0130_ ;
 wire \u_cpu.ALU.u_wallace._0131_ ;
 wire \u_cpu.ALU.u_wallace._0132_ ;
 wire \u_cpu.ALU.u_wallace._0133_ ;
 wire \u_cpu.ALU.u_wallace._0134_ ;
 wire \u_cpu.ALU.u_wallace._0135_ ;
 wire \u_cpu.ALU.u_wallace._0136_ ;
 wire \u_cpu.ALU.u_wallace._0137_ ;
 wire \u_cpu.ALU.u_wallace._0138_ ;
 wire \u_cpu.ALU.u_wallace._0139_ ;
 wire \u_cpu.ALU.u_wallace._0140_ ;
 wire \u_cpu.ALU.u_wallace._0141_ ;
 wire \u_cpu.ALU.u_wallace._0142_ ;
 wire \u_cpu.ALU.u_wallace._0143_ ;
 wire \u_cpu.ALU.u_wallace._0144_ ;
 wire \u_cpu.ALU.u_wallace._0145_ ;
 wire \u_cpu.ALU.u_wallace._0146_ ;
 wire \u_cpu.ALU.u_wallace._0147_ ;
 wire \u_cpu.ALU.u_wallace._0148_ ;
 wire \u_cpu.ALU.u_wallace._0149_ ;
 wire \u_cpu.ALU.u_wallace._0150_ ;
 wire \u_cpu.ALU.u_wallace._0151_ ;
 wire \u_cpu.ALU.u_wallace._0152_ ;
 wire \u_cpu.ALU.u_wallace._0153_ ;
 wire \u_cpu.ALU.u_wallace._0154_ ;
 wire \u_cpu.ALU.u_wallace._0155_ ;
 wire \u_cpu.ALU.u_wallace._0156_ ;
 wire \u_cpu.ALU.u_wallace._0157_ ;
 wire \u_cpu.ALU.u_wallace._0158_ ;
 wire \u_cpu.ALU.u_wallace._0159_ ;
 wire \u_cpu.ALU.u_wallace._0160_ ;
 wire \u_cpu.ALU.u_wallace._0161_ ;
 wire \u_cpu.ALU.u_wallace._0162_ ;
 wire \u_cpu.ALU.u_wallace._0163_ ;
 wire \u_cpu.ALU.u_wallace._0164_ ;
 wire \u_cpu.ALU.u_wallace._0165_ ;
 wire \u_cpu.ALU.u_wallace._0166_ ;
 wire \u_cpu.ALU.u_wallace._0167_ ;
 wire \u_cpu.ALU.u_wallace._0168_ ;
 wire \u_cpu.ALU.u_wallace._0169_ ;
 wire \u_cpu.ALU.u_wallace._0170_ ;
 wire \u_cpu.ALU.u_wallace._0171_ ;
 wire \u_cpu.ALU.u_wallace._0172_ ;
 wire \u_cpu.ALU.u_wallace._0173_ ;
 wire \u_cpu.ALU.u_wallace._0174_ ;
 wire \u_cpu.ALU.u_wallace._0175_ ;
 wire \u_cpu.ALU.u_wallace._0176_ ;
 wire \u_cpu.ALU.u_wallace._0177_ ;
 wire \u_cpu.ALU.u_wallace._0178_ ;
 wire \u_cpu.ALU.u_wallace._0179_ ;
 wire \u_cpu.ALU.u_wallace._0180_ ;
 wire \u_cpu.ALU.u_wallace._0181_ ;
 wire \u_cpu.ALU.u_wallace._0182_ ;
 wire \u_cpu.ALU.u_wallace._0183_ ;
 wire \u_cpu.ALU.u_wallace._0184_ ;
 wire \u_cpu.ALU.u_wallace._0185_ ;
 wire \u_cpu.ALU.u_wallace._0186_ ;
 wire \u_cpu.ALU.u_wallace._0187_ ;
 wire \u_cpu.ALU.u_wallace._0188_ ;
 wire \u_cpu.ALU.u_wallace._0189_ ;
 wire \u_cpu.ALU.u_wallace._0190_ ;
 wire \u_cpu.ALU.u_wallace._0191_ ;
 wire \u_cpu.ALU.u_wallace._0192_ ;
 wire \u_cpu.ALU.u_wallace._0193_ ;
 wire \u_cpu.ALU.u_wallace._0194_ ;
 wire \u_cpu.ALU.u_wallace._0195_ ;
 wire \u_cpu.ALU.u_wallace._0196_ ;
 wire \u_cpu.ALU.u_wallace._0197_ ;
 wire \u_cpu.ALU.u_wallace._0198_ ;
 wire \u_cpu.ALU.u_wallace._0199_ ;
 wire \u_cpu.ALU.u_wallace._0200_ ;
 wire \u_cpu.ALU.u_wallace._0201_ ;
 wire \u_cpu.ALU.u_wallace._0202_ ;
 wire \u_cpu.ALU.u_wallace._0203_ ;
 wire \u_cpu.ALU.u_wallace._0204_ ;
 wire \u_cpu.ALU.u_wallace._0205_ ;
 wire \u_cpu.ALU.u_wallace._0206_ ;
 wire \u_cpu.ALU.u_wallace._0207_ ;
 wire \u_cpu.ALU.u_wallace._0208_ ;
 wire \u_cpu.ALU.u_wallace._0209_ ;
 wire \u_cpu.ALU.u_wallace._0210_ ;
 wire \u_cpu.ALU.u_wallace._0211_ ;
 wire \u_cpu.ALU.u_wallace._0212_ ;
 wire \u_cpu.ALU.u_wallace._0213_ ;
 wire \u_cpu.ALU.u_wallace._0214_ ;
 wire \u_cpu.ALU.u_wallace._0215_ ;
 wire \u_cpu.ALU.u_wallace._0216_ ;
 wire \u_cpu.ALU.u_wallace._0217_ ;
 wire \u_cpu.ALU.u_wallace._0218_ ;
 wire \u_cpu.ALU.u_wallace._0219_ ;
 wire \u_cpu.ALU.u_wallace._0220_ ;
 wire \u_cpu.ALU.u_wallace._0221_ ;
 wire \u_cpu.ALU.u_wallace._0222_ ;
 wire \u_cpu.ALU.u_wallace._0223_ ;
 wire \u_cpu.ALU.u_wallace._0224_ ;
 wire \u_cpu.ALU.u_wallace._0225_ ;
 wire \u_cpu.ALU.u_wallace._0226_ ;
 wire \u_cpu.ALU.u_wallace._0227_ ;
 wire \u_cpu.ALU.u_wallace._0228_ ;
 wire \u_cpu.ALU.u_wallace._0229_ ;
 wire \u_cpu.ALU.u_wallace._0230_ ;
 wire \u_cpu.ALU.u_wallace._0231_ ;
 wire \u_cpu.ALU.u_wallace._0232_ ;
 wire \u_cpu.ALU.u_wallace._0233_ ;
 wire \u_cpu.ALU.u_wallace._0234_ ;
 wire \u_cpu.ALU.u_wallace._0235_ ;
 wire \u_cpu.ALU.u_wallace._0236_ ;
 wire \u_cpu.ALU.u_wallace._0237_ ;
 wire \u_cpu.ALU.u_wallace._0238_ ;
 wire \u_cpu.ALU.u_wallace._0239_ ;
 wire \u_cpu.ALU.u_wallace._0240_ ;
 wire \u_cpu.ALU.u_wallace._0241_ ;
 wire \u_cpu.ALU.u_wallace._0242_ ;
 wire \u_cpu.ALU.u_wallace._0243_ ;
 wire \u_cpu.ALU.u_wallace._0244_ ;
 wire \u_cpu.ALU.u_wallace._0245_ ;
 wire \u_cpu.ALU.u_wallace._0246_ ;
 wire \u_cpu.ALU.u_wallace._0247_ ;
 wire \u_cpu.ALU.u_wallace._0248_ ;
 wire \u_cpu.ALU.u_wallace._0249_ ;
 wire \u_cpu.ALU.u_wallace._0250_ ;
 wire \u_cpu.ALU.u_wallace._0251_ ;
 wire \u_cpu.ALU.u_wallace._0252_ ;
 wire \u_cpu.ALU.u_wallace._0253_ ;
 wire \u_cpu.ALU.u_wallace._0254_ ;
 wire \u_cpu.ALU.u_wallace._0255_ ;
 wire \u_cpu.ALU.u_wallace._0256_ ;
 wire \u_cpu.ALU.u_wallace._0257_ ;
 wire \u_cpu.ALU.u_wallace._0258_ ;
 wire \u_cpu.ALU.u_wallace._0259_ ;
 wire \u_cpu.ALU.u_wallace._0260_ ;
 wire \u_cpu.ALU.u_wallace._0261_ ;
 wire \u_cpu.ALU.u_wallace._0262_ ;
 wire \u_cpu.ALU.u_wallace._0263_ ;
 wire \u_cpu.ALU.u_wallace._0264_ ;
 wire \u_cpu.ALU.u_wallace._0265_ ;
 wire \u_cpu.ALU.u_wallace._0266_ ;
 wire \u_cpu.ALU.u_wallace._0267_ ;
 wire \u_cpu.ALU.u_wallace._0268_ ;
 wire \u_cpu.ALU.u_wallace._0269_ ;
 wire \u_cpu.ALU.u_wallace._0270_ ;
 wire \u_cpu.ALU.u_wallace._0271_ ;
 wire \u_cpu.ALU.u_wallace._0272_ ;
 wire \u_cpu.ALU.u_wallace._0273_ ;
 wire \u_cpu.ALU.u_wallace._0274_ ;
 wire \u_cpu.ALU.u_wallace._0275_ ;
 wire \u_cpu.ALU.u_wallace._0276_ ;
 wire \u_cpu.ALU.u_wallace._0277_ ;
 wire \u_cpu.ALU.u_wallace._0278_ ;
 wire \u_cpu.ALU.u_wallace._0279_ ;
 wire \u_cpu.ALU.u_wallace._0280_ ;
 wire \u_cpu.ALU.u_wallace._0281_ ;
 wire \u_cpu.ALU.u_wallace._0282_ ;
 wire \u_cpu.ALU.u_wallace._0283_ ;
 wire \u_cpu.ALU.u_wallace._0284_ ;
 wire \u_cpu.ALU.u_wallace._0285_ ;
 wire \u_cpu.ALU.u_wallace._0286_ ;
 wire \u_cpu.ALU.u_wallace._0287_ ;
 wire \u_cpu.ALU.u_wallace._0288_ ;
 wire \u_cpu.ALU.u_wallace._0289_ ;
 wire \u_cpu.ALU.u_wallace._0290_ ;
 wire \u_cpu.ALU.u_wallace._0291_ ;
 wire \u_cpu.ALU.u_wallace._0292_ ;
 wire \u_cpu.ALU.u_wallace._0293_ ;
 wire \u_cpu.ALU.u_wallace._0294_ ;
 wire \u_cpu.ALU.u_wallace._0295_ ;
 wire \u_cpu.ALU.u_wallace._0296_ ;
 wire \u_cpu.ALU.u_wallace._0297_ ;
 wire \u_cpu.ALU.u_wallace._0298_ ;
 wire \u_cpu.ALU.u_wallace._0299_ ;
 wire \u_cpu.ALU.u_wallace._0300_ ;
 wire \u_cpu.ALU.u_wallace._0301_ ;
 wire \u_cpu.ALU.u_wallace._0302_ ;
 wire \u_cpu.ALU.u_wallace._0303_ ;
 wire \u_cpu.ALU.u_wallace._0304_ ;
 wire \u_cpu.ALU.u_wallace._0305_ ;
 wire \u_cpu.ALU.u_wallace._0306_ ;
 wire \u_cpu.ALU.u_wallace._0307_ ;
 wire \u_cpu.ALU.u_wallace._0308_ ;
 wire \u_cpu.ALU.u_wallace._0309_ ;
 wire \u_cpu.ALU.u_wallace._0310_ ;
 wire \u_cpu.ALU.u_wallace._0311_ ;
 wire \u_cpu.ALU.u_wallace._0312_ ;
 wire \u_cpu.ALU.u_wallace._0313_ ;
 wire \u_cpu.ALU.u_wallace._0314_ ;
 wire \u_cpu.ALU.u_wallace._0315_ ;
 wire \u_cpu.ALU.u_wallace._0316_ ;
 wire \u_cpu.ALU.u_wallace._0317_ ;
 wire \u_cpu.ALU.u_wallace._0318_ ;
 wire \u_cpu.ALU.u_wallace._0319_ ;
 wire \u_cpu.ALU.u_wallace._0320_ ;
 wire \u_cpu.ALU.u_wallace._0321_ ;
 wire \u_cpu.ALU.u_wallace._0322_ ;
 wire \u_cpu.ALU.u_wallace._0323_ ;
 wire \u_cpu.ALU.u_wallace._0324_ ;
 wire \u_cpu.ALU.u_wallace._0325_ ;
 wire \u_cpu.ALU.u_wallace._0326_ ;
 wire \u_cpu.ALU.u_wallace._0327_ ;
 wire \u_cpu.ALU.u_wallace._0328_ ;
 wire \u_cpu.ALU.u_wallace._0329_ ;
 wire \u_cpu.ALU.u_wallace._0330_ ;
 wire \u_cpu.ALU.u_wallace._0331_ ;
 wire \u_cpu.ALU.u_wallace._0332_ ;
 wire \u_cpu.ALU.u_wallace._0333_ ;
 wire \u_cpu.ALU.u_wallace._0334_ ;
 wire \u_cpu.ALU.u_wallace._0335_ ;
 wire \u_cpu.ALU.u_wallace._0336_ ;
 wire \u_cpu.ALU.u_wallace._0337_ ;
 wire \u_cpu.ALU.u_wallace._0338_ ;
 wire \u_cpu.ALU.u_wallace._0339_ ;
 wire \u_cpu.ALU.u_wallace._0340_ ;
 wire \u_cpu.ALU.u_wallace._0341_ ;
 wire \u_cpu.ALU.u_wallace._0342_ ;
 wire \u_cpu.ALU.u_wallace._0343_ ;
 wire \u_cpu.ALU.u_wallace._0344_ ;
 wire \u_cpu.ALU.u_wallace._0345_ ;
 wire \u_cpu.ALU.u_wallace._0346_ ;
 wire \u_cpu.ALU.u_wallace._0347_ ;
 wire \u_cpu.ALU.u_wallace._0348_ ;
 wire \u_cpu.ALU.u_wallace._0349_ ;
 wire \u_cpu.ALU.u_wallace._0350_ ;
 wire \u_cpu.ALU.u_wallace._0351_ ;
 wire \u_cpu.ALU.u_wallace._0352_ ;
 wire \u_cpu.ALU.u_wallace._0353_ ;
 wire \u_cpu.ALU.u_wallace._0354_ ;
 wire \u_cpu.ALU.u_wallace._0355_ ;
 wire \u_cpu.ALU.u_wallace._0356_ ;
 wire \u_cpu.ALU.u_wallace._0357_ ;
 wire \u_cpu.ALU.u_wallace._0358_ ;
 wire \u_cpu.ALU.u_wallace._0359_ ;
 wire \u_cpu.ALU.u_wallace._0360_ ;
 wire \u_cpu.ALU.u_wallace._0361_ ;
 wire \u_cpu.ALU.u_wallace._0362_ ;
 wire \u_cpu.ALU.u_wallace._0363_ ;
 wire \u_cpu.ALU.u_wallace._0364_ ;
 wire \u_cpu.ALU.u_wallace._0365_ ;
 wire \u_cpu.ALU.u_wallace._0366_ ;
 wire \u_cpu.ALU.u_wallace._0367_ ;
 wire \u_cpu.ALU.u_wallace._0368_ ;
 wire \u_cpu.ALU.u_wallace._0369_ ;
 wire \u_cpu.ALU.u_wallace._0370_ ;
 wire \u_cpu.ALU.u_wallace._0371_ ;
 wire \u_cpu.ALU.u_wallace._0372_ ;
 wire \u_cpu.ALU.u_wallace._0373_ ;
 wire \u_cpu.ALU.u_wallace._0374_ ;
 wire \u_cpu.ALU.u_wallace._0375_ ;
 wire \u_cpu.ALU.u_wallace._0376_ ;
 wire \u_cpu.ALU.u_wallace._0377_ ;
 wire \u_cpu.ALU.u_wallace._0378_ ;
 wire \u_cpu.ALU.u_wallace._0379_ ;
 wire \u_cpu.ALU.u_wallace._0380_ ;
 wire \u_cpu.ALU.u_wallace._0381_ ;
 wire \u_cpu.ALU.u_wallace._0382_ ;
 wire \u_cpu.ALU.u_wallace._0383_ ;
 wire \u_cpu.ALU.u_wallace._0384_ ;
 wire \u_cpu.ALU.u_wallace._0385_ ;
 wire \u_cpu.ALU.u_wallace._0386_ ;
 wire \u_cpu.ALU.u_wallace._0387_ ;
 wire \u_cpu.ALU.u_wallace._0388_ ;
 wire \u_cpu.ALU.u_wallace._0389_ ;
 wire \u_cpu.ALU.u_wallace._0390_ ;
 wire \u_cpu.ALU.u_wallace._0391_ ;
 wire \u_cpu.ALU.u_wallace._0392_ ;
 wire \u_cpu.ALU.u_wallace._0393_ ;
 wire \u_cpu.ALU.u_wallace._0394_ ;
 wire \u_cpu.ALU.u_wallace._0395_ ;
 wire \u_cpu.ALU.u_wallace._0396_ ;
 wire \u_cpu.ALU.u_wallace._0397_ ;
 wire \u_cpu.ALU.u_wallace._0398_ ;
 wire \u_cpu.ALU.u_wallace._0399_ ;
 wire \u_cpu.ALU.u_wallace._0400_ ;
 wire \u_cpu.ALU.u_wallace._0401_ ;
 wire \u_cpu.ALU.u_wallace._0402_ ;
 wire \u_cpu.ALU.u_wallace._0403_ ;
 wire \u_cpu.ALU.u_wallace._0404_ ;
 wire \u_cpu.ALU.u_wallace._0405_ ;
 wire \u_cpu.ALU.u_wallace._0406_ ;
 wire \u_cpu.ALU.u_wallace._0407_ ;
 wire \u_cpu.ALU.u_wallace._0408_ ;
 wire \u_cpu.ALU.u_wallace._0409_ ;
 wire \u_cpu.ALU.u_wallace._0410_ ;
 wire \u_cpu.ALU.u_wallace._0411_ ;
 wire \u_cpu.ALU.u_wallace._0412_ ;
 wire \u_cpu.ALU.u_wallace._0413_ ;
 wire \u_cpu.ALU.u_wallace._0414_ ;
 wire \u_cpu.ALU.u_wallace._0415_ ;
 wire \u_cpu.ALU.u_wallace._0416_ ;
 wire \u_cpu.ALU.u_wallace._0417_ ;
 wire \u_cpu.ALU.u_wallace._0418_ ;
 wire \u_cpu.ALU.u_wallace._0419_ ;
 wire \u_cpu.ALU.u_wallace._0420_ ;
 wire \u_cpu.ALU.u_wallace._0421_ ;
 wire \u_cpu.ALU.u_wallace._0422_ ;
 wire \u_cpu.ALU.u_wallace._0423_ ;
 wire \u_cpu.ALU.u_wallace._0424_ ;
 wire \u_cpu.ALU.u_wallace._0425_ ;
 wire \u_cpu.ALU.u_wallace._0426_ ;
 wire \u_cpu.ALU.u_wallace._0427_ ;
 wire \u_cpu.ALU.u_wallace._0428_ ;
 wire \u_cpu.ALU.u_wallace._0429_ ;
 wire \u_cpu.ALU.u_wallace._0430_ ;
 wire \u_cpu.ALU.u_wallace._0431_ ;
 wire \u_cpu.ALU.u_wallace._0432_ ;
 wire \u_cpu.ALU.u_wallace._0433_ ;
 wire \u_cpu.ALU.u_wallace._0434_ ;
 wire \u_cpu.ALU.u_wallace._0435_ ;
 wire \u_cpu.ALU.u_wallace._0436_ ;
 wire \u_cpu.ALU.u_wallace._0437_ ;
 wire \u_cpu.ALU.u_wallace._0438_ ;
 wire \u_cpu.ALU.u_wallace._0439_ ;
 wire \u_cpu.ALU.u_wallace._0440_ ;
 wire \u_cpu.ALU.u_wallace._0441_ ;
 wire \u_cpu.ALU.u_wallace._0442_ ;
 wire \u_cpu.ALU.u_wallace._0443_ ;
 wire \u_cpu.ALU.u_wallace._0444_ ;
 wire \u_cpu.ALU.u_wallace._0445_ ;
 wire \u_cpu.ALU.u_wallace._0446_ ;
 wire \u_cpu.ALU.u_wallace._0447_ ;
 wire \u_cpu.ALU.u_wallace._0448_ ;
 wire \u_cpu.ALU.u_wallace._0449_ ;
 wire \u_cpu.ALU.u_wallace._0450_ ;
 wire \u_cpu.ALU.u_wallace._0451_ ;
 wire \u_cpu.ALU.u_wallace._0452_ ;
 wire \u_cpu.ALU.u_wallace._0453_ ;
 wire \u_cpu.ALU.u_wallace._0454_ ;
 wire \u_cpu.ALU.u_wallace._0455_ ;
 wire \u_cpu.ALU.u_wallace._0456_ ;
 wire \u_cpu.ALU.u_wallace._0457_ ;
 wire \u_cpu.ALU.u_wallace._0458_ ;
 wire \u_cpu.ALU.u_wallace._0459_ ;
 wire \u_cpu.ALU.u_wallace._0460_ ;
 wire \u_cpu.ALU.u_wallace._0461_ ;
 wire \u_cpu.ALU.u_wallace._0462_ ;
 wire \u_cpu.ALU.u_wallace._0463_ ;
 wire \u_cpu.ALU.u_wallace._0464_ ;
 wire \u_cpu.ALU.u_wallace._0465_ ;
 wire \u_cpu.ALU.u_wallace._0466_ ;
 wire \u_cpu.ALU.u_wallace._0467_ ;
 wire \u_cpu.ALU.u_wallace._0468_ ;
 wire \u_cpu.ALU.u_wallace._0469_ ;
 wire \u_cpu.ALU.u_wallace._0470_ ;
 wire \u_cpu.ALU.u_wallace._0471_ ;
 wire \u_cpu.ALU.u_wallace._0472_ ;
 wire \u_cpu.ALU.u_wallace._0473_ ;
 wire \u_cpu.ALU.u_wallace._0474_ ;
 wire \u_cpu.ALU.u_wallace._0475_ ;
 wire \u_cpu.ALU.u_wallace._0476_ ;
 wire \u_cpu.ALU.u_wallace._0477_ ;
 wire \u_cpu.ALU.u_wallace._0478_ ;
 wire \u_cpu.ALU.u_wallace._0479_ ;
 wire \u_cpu.ALU.u_wallace._0480_ ;
 wire \u_cpu.ALU.u_wallace._0481_ ;
 wire \u_cpu.ALU.u_wallace._0482_ ;
 wire \u_cpu.ALU.u_wallace._0483_ ;
 wire \u_cpu.ALU.u_wallace._0484_ ;
 wire \u_cpu.ALU.u_wallace._0485_ ;
 wire \u_cpu.ALU.u_wallace._0486_ ;
 wire \u_cpu.ALU.u_wallace._0487_ ;
 wire \u_cpu.ALU.u_wallace._0488_ ;
 wire \u_cpu.ALU.u_wallace._0489_ ;
 wire \u_cpu.ALU.u_wallace._0490_ ;
 wire \u_cpu.ALU.u_wallace._0491_ ;
 wire \u_cpu.ALU.u_wallace._0492_ ;
 wire \u_cpu.ALU.u_wallace._0493_ ;
 wire \u_cpu.ALU.u_wallace._0494_ ;
 wire \u_cpu.ALU.u_wallace._0495_ ;
 wire \u_cpu.ALU.u_wallace._0496_ ;
 wire \u_cpu.ALU.u_wallace._0497_ ;
 wire \u_cpu.ALU.u_wallace._0498_ ;
 wire \u_cpu.ALU.u_wallace._0499_ ;
 wire \u_cpu.ALU.u_wallace._0500_ ;
 wire \u_cpu.ALU.u_wallace._0501_ ;
 wire \u_cpu.ALU.u_wallace._0502_ ;
 wire \u_cpu.ALU.u_wallace._0503_ ;
 wire \u_cpu.ALU.u_wallace._0504_ ;
 wire \u_cpu.ALU.u_wallace._0505_ ;
 wire \u_cpu.ALU.u_wallace._0506_ ;
 wire \u_cpu.ALU.u_wallace._0507_ ;
 wire \u_cpu.ALU.u_wallace._0508_ ;
 wire \u_cpu.ALU.u_wallace._0509_ ;
 wire \u_cpu.ALU.u_wallace._0510_ ;
 wire \u_cpu.ALU.u_wallace._0511_ ;
 wire \u_cpu.ALU.u_wallace._0512_ ;
 wire \u_cpu.ALU.u_wallace._0513_ ;
 wire \u_cpu.ALU.u_wallace._0514_ ;
 wire \u_cpu.ALU.u_wallace._0515_ ;
 wire \u_cpu.ALU.u_wallace._0516_ ;
 wire \u_cpu.ALU.u_wallace._0517_ ;
 wire \u_cpu.ALU.u_wallace._0518_ ;
 wire \u_cpu.ALU.u_wallace._0519_ ;
 wire \u_cpu.ALU.u_wallace._0520_ ;
 wire \u_cpu.ALU.u_wallace._0521_ ;
 wire \u_cpu.ALU.u_wallace._0522_ ;
 wire \u_cpu.ALU.u_wallace._0523_ ;
 wire \u_cpu.ALU.u_wallace._0524_ ;
 wire \u_cpu.ALU.u_wallace._0525_ ;
 wire \u_cpu.ALU.u_wallace._0526_ ;
 wire \u_cpu.ALU.u_wallace._0527_ ;
 wire \u_cpu.ALU.u_wallace._0528_ ;
 wire \u_cpu.ALU.u_wallace._0529_ ;
 wire \u_cpu.ALU.u_wallace._0530_ ;
 wire \u_cpu.ALU.u_wallace._0531_ ;
 wire \u_cpu.ALU.u_wallace._0532_ ;
 wire \u_cpu.ALU.u_wallace._0533_ ;
 wire \u_cpu.ALU.u_wallace._0534_ ;
 wire \u_cpu.ALU.u_wallace._0535_ ;
 wire \u_cpu.ALU.u_wallace._0536_ ;
 wire \u_cpu.ALU.u_wallace._0537_ ;
 wire \u_cpu.ALU.u_wallace._0538_ ;
 wire \u_cpu.ALU.u_wallace._0539_ ;
 wire \u_cpu.ALU.u_wallace._0540_ ;
 wire \u_cpu.ALU.u_wallace._0541_ ;
 wire \u_cpu.ALU.u_wallace._0542_ ;
 wire \u_cpu.ALU.u_wallace._0543_ ;
 wire \u_cpu.ALU.u_wallace._0544_ ;
 wire \u_cpu.ALU.u_wallace._0545_ ;
 wire \u_cpu.ALU.u_wallace._0546_ ;
 wire \u_cpu.ALU.u_wallace._0547_ ;
 wire \u_cpu.ALU.u_wallace._0548_ ;
 wire \u_cpu.ALU.u_wallace._0549_ ;
 wire \u_cpu.ALU.u_wallace._0550_ ;
 wire \u_cpu.ALU.u_wallace._0551_ ;
 wire \u_cpu.ALU.u_wallace._0552_ ;
 wire \u_cpu.ALU.u_wallace._0553_ ;
 wire \u_cpu.ALU.u_wallace._0554_ ;
 wire \u_cpu.ALU.u_wallace._0555_ ;
 wire \u_cpu.ALU.u_wallace._0556_ ;
 wire \u_cpu.ALU.u_wallace._0557_ ;
 wire \u_cpu.ALU.u_wallace._0558_ ;
 wire \u_cpu.ALU.u_wallace._0559_ ;
 wire \u_cpu.ALU.u_wallace._0560_ ;
 wire \u_cpu.ALU.u_wallace._0561_ ;
 wire \u_cpu.ALU.u_wallace._0562_ ;
 wire \u_cpu.ALU.u_wallace._0563_ ;
 wire \u_cpu.ALU.u_wallace._0564_ ;
 wire \u_cpu.ALU.u_wallace._0565_ ;
 wire \u_cpu.ALU.u_wallace._0566_ ;
 wire \u_cpu.ALU.u_wallace._0567_ ;
 wire \u_cpu.ALU.u_wallace._0568_ ;
 wire \u_cpu.ALU.u_wallace._0569_ ;
 wire \u_cpu.ALU.u_wallace._0570_ ;
 wire \u_cpu.ALU.u_wallace._0571_ ;
 wire \u_cpu.ALU.u_wallace._0572_ ;
 wire \u_cpu.ALU.u_wallace._0573_ ;
 wire \u_cpu.ALU.u_wallace._0574_ ;
 wire \u_cpu.ALU.u_wallace._0575_ ;
 wire \u_cpu.ALU.u_wallace._0576_ ;
 wire \u_cpu.ALU.u_wallace._0577_ ;
 wire \u_cpu.ALU.u_wallace._0578_ ;
 wire \u_cpu.ALU.u_wallace._0579_ ;
 wire \u_cpu.ALU.u_wallace._0580_ ;
 wire \u_cpu.ALU.u_wallace._0581_ ;
 wire \u_cpu.ALU.u_wallace._0582_ ;
 wire \u_cpu.ALU.u_wallace._0583_ ;
 wire \u_cpu.ALU.u_wallace._0584_ ;
 wire \u_cpu.ALU.u_wallace._0585_ ;
 wire \u_cpu.ALU.u_wallace._0586_ ;
 wire \u_cpu.ALU.u_wallace._0587_ ;
 wire \u_cpu.ALU.u_wallace._0588_ ;
 wire \u_cpu.ALU.u_wallace._0589_ ;
 wire \u_cpu.ALU.u_wallace._0590_ ;
 wire \u_cpu.ALU.u_wallace._0591_ ;
 wire \u_cpu.ALU.u_wallace._0592_ ;
 wire \u_cpu.ALU.u_wallace._0593_ ;
 wire \u_cpu.ALU.u_wallace._0594_ ;
 wire \u_cpu.ALU.u_wallace._0595_ ;
 wire \u_cpu.ALU.u_wallace._0596_ ;
 wire \u_cpu.ALU.u_wallace._0597_ ;
 wire \u_cpu.ALU.u_wallace._0598_ ;
 wire \u_cpu.ALU.u_wallace._0599_ ;
 wire \u_cpu.ALU.u_wallace._0600_ ;
 wire \u_cpu.ALU.u_wallace._0601_ ;
 wire \u_cpu.ALU.u_wallace._0602_ ;
 wire \u_cpu.ALU.u_wallace._0603_ ;
 wire \u_cpu.ALU.u_wallace._0604_ ;
 wire \u_cpu.ALU.u_wallace._0605_ ;
 wire \u_cpu.ALU.u_wallace._0606_ ;
 wire \u_cpu.ALU.u_wallace._0607_ ;
 wire \u_cpu.ALU.u_wallace._0608_ ;
 wire \u_cpu.ALU.u_wallace._0609_ ;
 wire \u_cpu.ALU.u_wallace._0610_ ;
 wire \u_cpu.ALU.u_wallace._0611_ ;
 wire \u_cpu.ALU.u_wallace._0612_ ;
 wire \u_cpu.ALU.u_wallace._0613_ ;
 wire \u_cpu.ALU.u_wallace._0614_ ;
 wire \u_cpu.ALU.u_wallace._0615_ ;
 wire \u_cpu.ALU.u_wallace._0616_ ;
 wire \u_cpu.ALU.u_wallace._0617_ ;
 wire \u_cpu.ALU.u_wallace._0618_ ;
 wire \u_cpu.ALU.u_wallace._0619_ ;
 wire \u_cpu.ALU.u_wallace._0620_ ;
 wire \u_cpu.ALU.u_wallace._0621_ ;
 wire \u_cpu.ALU.u_wallace._0622_ ;
 wire \u_cpu.ALU.u_wallace._0623_ ;
 wire \u_cpu.ALU.u_wallace._0624_ ;
 wire \u_cpu.ALU.u_wallace._0625_ ;
 wire \u_cpu.ALU.u_wallace._0626_ ;
 wire \u_cpu.ALU.u_wallace._0627_ ;
 wire \u_cpu.ALU.u_wallace._0628_ ;
 wire \u_cpu.ALU.u_wallace._0629_ ;
 wire \u_cpu.ALU.u_wallace._0630_ ;
 wire \u_cpu.ALU.u_wallace._0631_ ;
 wire \u_cpu.ALU.u_wallace._0632_ ;
 wire \u_cpu.ALU.u_wallace._0633_ ;
 wire \u_cpu.ALU.u_wallace._0634_ ;
 wire \u_cpu.ALU.u_wallace._0635_ ;
 wire \u_cpu.ALU.u_wallace._0636_ ;
 wire \u_cpu.ALU.u_wallace._0637_ ;
 wire \u_cpu.ALU.u_wallace._0638_ ;
 wire \u_cpu.ALU.u_wallace._0639_ ;
 wire \u_cpu.ALU.u_wallace._0640_ ;
 wire \u_cpu.ALU.u_wallace._0641_ ;
 wire \u_cpu.ALU.u_wallace._0642_ ;
 wire \u_cpu.ALU.u_wallace._0643_ ;
 wire \u_cpu.ALU.u_wallace._0644_ ;
 wire \u_cpu.ALU.u_wallace._0645_ ;
 wire \u_cpu.ALU.u_wallace._0646_ ;
 wire \u_cpu.ALU.u_wallace._0647_ ;
 wire \u_cpu.ALU.u_wallace._0648_ ;
 wire \u_cpu.ALU.u_wallace._0649_ ;
 wire \u_cpu.ALU.u_wallace._0650_ ;
 wire \u_cpu.ALU.u_wallace._0651_ ;
 wire \u_cpu.ALU.u_wallace._0652_ ;
 wire \u_cpu.ALU.u_wallace._0653_ ;
 wire \u_cpu.ALU.u_wallace._0654_ ;
 wire \u_cpu.ALU.u_wallace._0655_ ;
 wire \u_cpu.ALU.u_wallace._0656_ ;
 wire \u_cpu.ALU.u_wallace._0657_ ;
 wire \u_cpu.ALU.u_wallace._0658_ ;
 wire \u_cpu.ALU.u_wallace._0659_ ;
 wire \u_cpu.ALU.u_wallace._0660_ ;
 wire \u_cpu.ALU.u_wallace._0661_ ;
 wire \u_cpu.ALU.u_wallace._0662_ ;
 wire \u_cpu.ALU.u_wallace._0663_ ;
 wire \u_cpu.ALU.u_wallace._0664_ ;
 wire \u_cpu.ALU.u_wallace._0665_ ;
 wire \u_cpu.ALU.u_wallace._0666_ ;
 wire \u_cpu.ALU.u_wallace._0667_ ;
 wire \u_cpu.ALU.u_wallace._0668_ ;
 wire \u_cpu.ALU.u_wallace._0669_ ;
 wire \u_cpu.ALU.u_wallace._0670_ ;
 wire \u_cpu.ALU.u_wallace._0671_ ;
 wire \u_cpu.ALU.u_wallace._0672_ ;
 wire \u_cpu.ALU.u_wallace._0673_ ;
 wire \u_cpu.ALU.u_wallace._0674_ ;
 wire \u_cpu.ALU.u_wallace._0675_ ;
 wire \u_cpu.ALU.u_wallace._0676_ ;
 wire \u_cpu.ALU.u_wallace._0677_ ;
 wire \u_cpu.ALU.u_wallace._0678_ ;
 wire \u_cpu.ALU.u_wallace._0679_ ;
 wire \u_cpu.ALU.u_wallace._0680_ ;
 wire \u_cpu.ALU.u_wallace._0681_ ;
 wire \u_cpu.ALU.u_wallace._0682_ ;
 wire \u_cpu.ALU.u_wallace._0683_ ;
 wire \u_cpu.ALU.u_wallace._0684_ ;
 wire \u_cpu.ALU.u_wallace._0685_ ;
 wire \u_cpu.ALU.u_wallace._0686_ ;
 wire \u_cpu.ALU.u_wallace._0687_ ;
 wire \u_cpu.ALU.u_wallace._0688_ ;
 wire \u_cpu.ALU.u_wallace._0689_ ;
 wire \u_cpu.ALU.u_wallace._0690_ ;
 wire \u_cpu.ALU.u_wallace._0691_ ;
 wire \u_cpu.ALU.u_wallace._0692_ ;
 wire \u_cpu.ALU.u_wallace._0693_ ;
 wire \u_cpu.ALU.u_wallace._0694_ ;
 wire \u_cpu.ALU.u_wallace._0695_ ;
 wire \u_cpu.ALU.u_wallace._0696_ ;
 wire \u_cpu.ALU.u_wallace._0697_ ;
 wire \u_cpu.ALU.u_wallace._0698_ ;
 wire \u_cpu.ALU.u_wallace._0699_ ;
 wire \u_cpu.ALU.u_wallace._0700_ ;
 wire \u_cpu.ALU.u_wallace._0701_ ;
 wire \u_cpu.ALU.u_wallace._0702_ ;
 wire \u_cpu.ALU.u_wallace._0703_ ;
 wire \u_cpu.ALU.u_wallace._0704_ ;
 wire \u_cpu.ALU.u_wallace._0705_ ;
 wire \u_cpu.ALU.u_wallace._0706_ ;
 wire \u_cpu.ALU.u_wallace._0707_ ;
 wire \u_cpu.ALU.u_wallace._0708_ ;
 wire \u_cpu.ALU.u_wallace._0709_ ;
 wire \u_cpu.ALU.u_wallace._0710_ ;
 wire \u_cpu.ALU.u_wallace._0711_ ;
 wire \u_cpu.ALU.u_wallace._0712_ ;
 wire \u_cpu.ALU.u_wallace._0713_ ;
 wire \u_cpu.ALU.u_wallace._0714_ ;
 wire \u_cpu.ALU.u_wallace._0715_ ;
 wire \u_cpu.ALU.u_wallace._0716_ ;
 wire \u_cpu.ALU.u_wallace._0717_ ;
 wire \u_cpu.ALU.u_wallace._0718_ ;
 wire \u_cpu.ALU.u_wallace._0719_ ;
 wire \u_cpu.ALU.u_wallace._0720_ ;
 wire \u_cpu.ALU.u_wallace._0721_ ;
 wire \u_cpu.ALU.u_wallace._0722_ ;
 wire \u_cpu.ALU.u_wallace._0723_ ;
 wire \u_cpu.ALU.u_wallace._0724_ ;
 wire \u_cpu.ALU.u_wallace._0725_ ;
 wire \u_cpu.ALU.u_wallace._0726_ ;
 wire \u_cpu.ALU.u_wallace._0727_ ;
 wire \u_cpu.ALU.u_wallace._0728_ ;
 wire \u_cpu.ALU.u_wallace._0729_ ;
 wire \u_cpu.ALU.u_wallace._0730_ ;
 wire \u_cpu.ALU.u_wallace._0731_ ;
 wire \u_cpu.ALU.u_wallace._0732_ ;
 wire \u_cpu.ALU.u_wallace._0733_ ;
 wire \u_cpu.ALU.u_wallace._0734_ ;
 wire \u_cpu.ALU.u_wallace._0735_ ;
 wire \u_cpu.ALU.u_wallace._0736_ ;
 wire \u_cpu.ALU.u_wallace._0737_ ;
 wire \u_cpu.ALU.u_wallace._0738_ ;
 wire \u_cpu.ALU.u_wallace._0739_ ;
 wire \u_cpu.ALU.u_wallace._0740_ ;
 wire \u_cpu.ALU.u_wallace._0741_ ;
 wire \u_cpu.ALU.u_wallace._0742_ ;
 wire \u_cpu.ALU.u_wallace._0743_ ;
 wire \u_cpu.ALU.u_wallace._0744_ ;
 wire \u_cpu.ALU.u_wallace._0745_ ;
 wire \u_cpu.ALU.u_wallace._0746_ ;
 wire \u_cpu.ALU.u_wallace._0747_ ;
 wire \u_cpu.ALU.u_wallace._0748_ ;
 wire \u_cpu.ALU.u_wallace._0749_ ;
 wire \u_cpu.ALU.u_wallace._0750_ ;
 wire \u_cpu.ALU.u_wallace._0751_ ;
 wire \u_cpu.ALU.u_wallace._0752_ ;
 wire \u_cpu.ALU.u_wallace._0753_ ;
 wire \u_cpu.ALU.u_wallace._0754_ ;
 wire \u_cpu.ALU.u_wallace._0755_ ;
 wire \u_cpu.ALU.u_wallace._0756_ ;
 wire \u_cpu.ALU.u_wallace._0757_ ;
 wire \u_cpu.ALU.u_wallace._0758_ ;
 wire \u_cpu.ALU.u_wallace._0759_ ;
 wire \u_cpu.ALU.u_wallace._0760_ ;
 wire \u_cpu.ALU.u_wallace._0761_ ;
 wire \u_cpu.ALU.u_wallace._0762_ ;
 wire \u_cpu.ALU.u_wallace._0763_ ;
 wire \u_cpu.ALU.u_wallace._0764_ ;
 wire \u_cpu.ALU.u_wallace._0765_ ;
 wire \u_cpu.ALU.u_wallace._0766_ ;
 wire \u_cpu.ALU.u_wallace._0767_ ;
 wire \u_cpu.ALU.u_wallace._0768_ ;
 wire \u_cpu.ALU.u_wallace._0769_ ;
 wire \u_cpu.ALU.u_wallace._0770_ ;
 wire \u_cpu.ALU.u_wallace._0771_ ;
 wire \u_cpu.ALU.u_wallace._0772_ ;
 wire \u_cpu.ALU.u_wallace._0773_ ;
 wire \u_cpu.ALU.u_wallace._0774_ ;
 wire \u_cpu.ALU.u_wallace._0775_ ;
 wire \u_cpu.ALU.u_wallace._0776_ ;
 wire \u_cpu.ALU.u_wallace._0777_ ;
 wire \u_cpu.ALU.u_wallace._0778_ ;
 wire \u_cpu.ALU.u_wallace._0779_ ;
 wire \u_cpu.ALU.u_wallace._0780_ ;
 wire \u_cpu.ALU.u_wallace._0781_ ;
 wire \u_cpu.ALU.u_wallace._0782_ ;
 wire \u_cpu.ALU.u_wallace._0783_ ;
 wire \u_cpu.ALU.u_wallace._0784_ ;
 wire \u_cpu.ALU.u_wallace._0785_ ;
 wire \u_cpu.ALU.u_wallace._0786_ ;
 wire \u_cpu.ALU.u_wallace._0787_ ;
 wire \u_cpu.ALU.u_wallace._0788_ ;
 wire \u_cpu.ALU.u_wallace._0789_ ;
 wire \u_cpu.ALU.u_wallace._0790_ ;
 wire \u_cpu.ALU.u_wallace._0791_ ;
 wire \u_cpu.ALU.u_wallace._0792_ ;
 wire \u_cpu.ALU.u_wallace._0793_ ;
 wire \u_cpu.ALU.u_wallace._0794_ ;
 wire \u_cpu.ALU.u_wallace._0795_ ;
 wire \u_cpu.ALU.u_wallace._0796_ ;
 wire \u_cpu.ALU.u_wallace._0797_ ;
 wire \u_cpu.ALU.u_wallace._0798_ ;
 wire \u_cpu.ALU.u_wallace._0799_ ;
 wire \u_cpu.ALU.u_wallace._0800_ ;
 wire \u_cpu.ALU.u_wallace._0801_ ;
 wire \u_cpu.ALU.u_wallace._0802_ ;
 wire \u_cpu.ALU.u_wallace._0803_ ;
 wire \u_cpu.ALU.u_wallace._0804_ ;
 wire \u_cpu.ALU.u_wallace._0805_ ;
 wire \u_cpu.ALU.u_wallace._0806_ ;
 wire \u_cpu.ALU.u_wallace._0807_ ;
 wire \u_cpu.ALU.u_wallace._0808_ ;
 wire \u_cpu.ALU.u_wallace._0809_ ;
 wire \u_cpu.ALU.u_wallace._0810_ ;
 wire \u_cpu.ALU.u_wallace._0811_ ;
 wire \u_cpu.ALU.u_wallace._0812_ ;
 wire \u_cpu.ALU.u_wallace._0813_ ;
 wire \u_cpu.ALU.u_wallace._0814_ ;
 wire \u_cpu.ALU.u_wallace._0815_ ;
 wire \u_cpu.ALU.u_wallace._0816_ ;
 wire \u_cpu.ALU.u_wallace._0817_ ;
 wire \u_cpu.ALU.u_wallace._0818_ ;
 wire \u_cpu.ALU.u_wallace._0819_ ;
 wire \u_cpu.ALU.u_wallace._0820_ ;
 wire \u_cpu.ALU.u_wallace._0821_ ;
 wire \u_cpu.ALU.u_wallace._0822_ ;
 wire \u_cpu.ALU.u_wallace._0823_ ;
 wire \u_cpu.ALU.u_wallace._0824_ ;
 wire \u_cpu.ALU.u_wallace._0825_ ;
 wire \u_cpu.ALU.u_wallace._0826_ ;
 wire \u_cpu.ALU.u_wallace._0827_ ;
 wire \u_cpu.ALU.u_wallace._0828_ ;
 wire \u_cpu.ALU.u_wallace._0829_ ;
 wire \u_cpu.ALU.u_wallace._0830_ ;
 wire \u_cpu.ALU.u_wallace._0831_ ;
 wire \u_cpu.ALU.u_wallace._0832_ ;
 wire \u_cpu.ALU.u_wallace._0833_ ;
 wire \u_cpu.ALU.u_wallace._0834_ ;
 wire \u_cpu.ALU.u_wallace._0835_ ;
 wire \u_cpu.ALU.u_wallace._0836_ ;
 wire \u_cpu.ALU.u_wallace._0837_ ;
 wire \u_cpu.ALU.u_wallace._0838_ ;
 wire \u_cpu.ALU.u_wallace._0839_ ;
 wire \u_cpu.ALU.u_wallace._0840_ ;
 wire \u_cpu.ALU.u_wallace._0841_ ;
 wire \u_cpu.ALU.u_wallace._0842_ ;
 wire \u_cpu.ALU.u_wallace._0843_ ;
 wire \u_cpu.ALU.u_wallace._0844_ ;
 wire \u_cpu.ALU.u_wallace._0845_ ;
 wire \u_cpu.ALU.u_wallace._0846_ ;
 wire \u_cpu.ALU.u_wallace._0847_ ;
 wire \u_cpu.ALU.u_wallace._0848_ ;
 wire \u_cpu.ALU.u_wallace._0849_ ;
 wire \u_cpu.ALU.u_wallace._0850_ ;
 wire \u_cpu.ALU.u_wallace._0851_ ;
 wire \u_cpu.ALU.u_wallace._0852_ ;
 wire \u_cpu.ALU.u_wallace._0853_ ;
 wire \u_cpu.ALU.u_wallace._0854_ ;
 wire \u_cpu.ALU.u_wallace._0855_ ;
 wire \u_cpu.ALU.u_wallace._0856_ ;
 wire \u_cpu.ALU.u_wallace._0857_ ;
 wire \u_cpu.ALU.u_wallace._0858_ ;
 wire \u_cpu.ALU.u_wallace._0859_ ;
 wire \u_cpu.ALU.u_wallace._0860_ ;
 wire \u_cpu.ALU.u_wallace._0861_ ;
 wire \u_cpu.ALU.u_wallace._0862_ ;
 wire \u_cpu.ALU.u_wallace._0863_ ;
 wire \u_cpu.ALU.u_wallace._0864_ ;
 wire \u_cpu.ALU.u_wallace._0865_ ;
 wire \u_cpu.ALU.u_wallace._0866_ ;
 wire \u_cpu.ALU.u_wallace._0867_ ;
 wire \u_cpu.ALU.u_wallace._0868_ ;
 wire \u_cpu.ALU.u_wallace._0869_ ;
 wire \u_cpu.ALU.u_wallace._0870_ ;
 wire \u_cpu.ALU.u_wallace._0871_ ;
 wire \u_cpu.ALU.u_wallace._0872_ ;
 wire \u_cpu.ALU.u_wallace._0873_ ;
 wire \u_cpu.ALU.u_wallace._0874_ ;
 wire \u_cpu.ALU.u_wallace._0875_ ;
 wire \u_cpu.ALU.u_wallace._0876_ ;
 wire \u_cpu.ALU.u_wallace._0877_ ;
 wire \u_cpu.ALU.u_wallace._0878_ ;
 wire \u_cpu.ALU.u_wallace._0879_ ;
 wire \u_cpu.ALU.u_wallace._0880_ ;
 wire \u_cpu.ALU.u_wallace._0881_ ;
 wire \u_cpu.ALU.u_wallace._0882_ ;
 wire \u_cpu.ALU.u_wallace._0883_ ;
 wire \u_cpu.ALU.u_wallace._0884_ ;
 wire \u_cpu.ALU.u_wallace._0885_ ;
 wire \u_cpu.ALU.u_wallace._0886_ ;
 wire \u_cpu.ALU.u_wallace._0887_ ;
 wire \u_cpu.ALU.u_wallace._0888_ ;
 wire \u_cpu.ALU.u_wallace._0889_ ;
 wire \u_cpu.ALU.u_wallace._0890_ ;
 wire \u_cpu.ALU.u_wallace._0891_ ;
 wire \u_cpu.ALU.u_wallace._0892_ ;
 wire \u_cpu.ALU.u_wallace._0893_ ;
 wire \u_cpu.ALU.u_wallace._0894_ ;
 wire \u_cpu.ALU.u_wallace._0895_ ;
 wire \u_cpu.ALU.u_wallace._0896_ ;
 wire \u_cpu.ALU.u_wallace._0897_ ;
 wire \u_cpu.ALU.u_wallace._0898_ ;
 wire \u_cpu.ALU.u_wallace._0899_ ;
 wire \u_cpu.ALU.u_wallace._0900_ ;
 wire \u_cpu.ALU.u_wallace._0901_ ;
 wire \u_cpu.ALU.u_wallace._0902_ ;
 wire \u_cpu.ALU.u_wallace._0903_ ;
 wire \u_cpu.ALU.u_wallace._0904_ ;
 wire \u_cpu.ALU.u_wallace._0905_ ;
 wire \u_cpu.ALU.u_wallace._0906_ ;
 wire \u_cpu.ALU.u_wallace._0907_ ;
 wire \u_cpu.ALU.u_wallace._0908_ ;
 wire \u_cpu.ALU.u_wallace._0909_ ;
 wire \u_cpu.ALU.u_wallace._0910_ ;
 wire \u_cpu.ALU.u_wallace._0911_ ;
 wire \u_cpu.ALU.u_wallace._0912_ ;
 wire \u_cpu.ALU.u_wallace._0913_ ;
 wire \u_cpu.ALU.u_wallace._0914_ ;
 wire \u_cpu.ALU.u_wallace._0915_ ;
 wire \u_cpu.ALU.u_wallace._0916_ ;
 wire \u_cpu.ALU.u_wallace._0917_ ;
 wire \u_cpu.ALU.u_wallace._0918_ ;
 wire \u_cpu.ALU.u_wallace._0919_ ;
 wire \u_cpu.ALU.u_wallace._0920_ ;
 wire \u_cpu.ALU.u_wallace._0921_ ;
 wire \u_cpu.ALU.u_wallace._0922_ ;
 wire \u_cpu.ALU.u_wallace._0923_ ;
 wire \u_cpu.ALU.u_wallace._0924_ ;
 wire \u_cpu.ALU.u_wallace._0925_ ;
 wire \u_cpu.ALU.u_wallace._0926_ ;
 wire \u_cpu.ALU.u_wallace._0927_ ;
 wire \u_cpu.ALU.u_wallace._0928_ ;
 wire \u_cpu.ALU.u_wallace._0929_ ;
 wire \u_cpu.ALU.u_wallace._0930_ ;
 wire \u_cpu.ALU.u_wallace._0931_ ;
 wire \u_cpu.ALU.u_wallace._0932_ ;
 wire \u_cpu.ALU.u_wallace._0933_ ;
 wire \u_cpu.ALU.u_wallace._0934_ ;
 wire \u_cpu.ALU.u_wallace._0935_ ;
 wire \u_cpu.ALU.u_wallace._0936_ ;
 wire \u_cpu.ALU.u_wallace._0937_ ;
 wire \u_cpu.ALU.u_wallace._0938_ ;
 wire \u_cpu.ALU.u_wallace._0939_ ;
 wire \u_cpu.ALU.u_wallace._0940_ ;
 wire \u_cpu.ALU.u_wallace._0941_ ;
 wire \u_cpu.ALU.u_wallace._0942_ ;
 wire \u_cpu.ALU.u_wallace._0943_ ;
 wire \u_cpu.ALU.u_wallace._0944_ ;
 wire \u_cpu.ALU.u_wallace._0945_ ;
 wire \u_cpu.ALU.u_wallace._0946_ ;
 wire \u_cpu.ALU.u_wallace._0947_ ;
 wire \u_cpu.ALU.u_wallace._0948_ ;
 wire \u_cpu.ALU.u_wallace._0949_ ;
 wire \u_cpu.ALU.u_wallace._0950_ ;
 wire \u_cpu.ALU.u_wallace._0951_ ;
 wire \u_cpu.ALU.u_wallace._0952_ ;
 wire \u_cpu.ALU.u_wallace._0953_ ;
 wire \u_cpu.ALU.u_wallace._0954_ ;
 wire \u_cpu.ALU.u_wallace._0955_ ;
 wire \u_cpu.ALU.u_wallace._0956_ ;
 wire \u_cpu.ALU.u_wallace._0957_ ;
 wire \u_cpu.ALU.u_wallace._0958_ ;
 wire \u_cpu.ALU.u_wallace._0959_ ;
 wire \u_cpu.ALU.u_wallace._0960_ ;
 wire \u_cpu.ALU.u_wallace._0961_ ;
 wire \u_cpu.ALU.u_wallace._0962_ ;
 wire \u_cpu.ALU.u_wallace._0963_ ;
 wire \u_cpu.ALU.u_wallace._0964_ ;
 wire \u_cpu.ALU.u_wallace._0965_ ;
 wire \u_cpu.ALU.u_wallace._0966_ ;
 wire \u_cpu.ALU.u_wallace._0967_ ;
 wire \u_cpu.ALU.u_wallace._0968_ ;
 wire \u_cpu.ALU.u_wallace._0969_ ;
 wire \u_cpu.ALU.u_wallace._0970_ ;
 wire \u_cpu.ALU.u_wallace._0971_ ;
 wire \u_cpu.ALU.u_wallace._0972_ ;
 wire \u_cpu.ALU.u_wallace._0973_ ;
 wire \u_cpu.ALU.u_wallace._0974_ ;
 wire \u_cpu.ALU.u_wallace._0975_ ;
 wire \u_cpu.ALU.u_wallace._0976_ ;
 wire \u_cpu.ALU.u_wallace._0977_ ;
 wire \u_cpu.ALU.u_wallace._0978_ ;
 wire \u_cpu.ALU.u_wallace._0979_ ;
 wire \u_cpu.ALU.u_wallace._0980_ ;
 wire \u_cpu.ALU.u_wallace._0981_ ;
 wire \u_cpu.ALU.u_wallace._0982_ ;
 wire \u_cpu.ALU.u_wallace._0983_ ;
 wire \u_cpu.ALU.u_wallace._0984_ ;
 wire \u_cpu.ALU.u_wallace._0985_ ;
 wire \u_cpu.ALU.u_wallace._0986_ ;
 wire \u_cpu.ALU.u_wallace._0987_ ;
 wire \u_cpu.ALU.u_wallace._0988_ ;
 wire \u_cpu.ALU.u_wallace._0989_ ;
 wire \u_cpu.ALU.u_wallace._0990_ ;
 wire \u_cpu.ALU.u_wallace._0991_ ;
 wire \u_cpu.ALU.u_wallace._0992_ ;
 wire \u_cpu.ALU.u_wallace._0993_ ;
 wire \u_cpu.ALU.u_wallace._0994_ ;
 wire \u_cpu.ALU.u_wallace._0995_ ;
 wire \u_cpu.ALU.u_wallace._0996_ ;
 wire \u_cpu.ALU.u_wallace._0997_ ;
 wire \u_cpu.ALU.u_wallace._0998_ ;
 wire \u_cpu.ALU.u_wallace._0999_ ;
 wire \u_cpu.ALU.u_wallace._1000_ ;
 wire \u_cpu.ALU.u_wallace._1001_ ;
 wire \u_cpu.ALU.u_wallace._1002_ ;
 wire \u_cpu.ALU.u_wallace._1003_ ;
 wire \u_cpu.ALU.u_wallace._1004_ ;
 wire \u_cpu.ALU.u_wallace._1005_ ;
 wire \u_cpu.ALU.u_wallace._1006_ ;
 wire \u_cpu.ALU.u_wallace._1007_ ;
 wire \u_cpu.ALU.u_wallace._1008_ ;
 wire \u_cpu.ALU.u_wallace._1009_ ;
 wire \u_cpu.ALU.u_wallace._1010_ ;
 wire \u_cpu.ALU.u_wallace._1011_ ;
 wire \u_cpu.ALU.u_wallace._1012_ ;
 wire \u_cpu.ALU.u_wallace._1013_ ;
 wire \u_cpu.ALU.u_wallace._1014_ ;
 wire \u_cpu.ALU.u_wallace._1015_ ;
 wire \u_cpu.ALU.u_wallace._1016_ ;
 wire \u_cpu.ALU.u_wallace._1017_ ;
 wire \u_cpu.ALU.u_wallace._1018_ ;
 wire \u_cpu.ALU.u_wallace._1019_ ;
 wire \u_cpu.ALU.u_wallace._1020_ ;
 wire \u_cpu.ALU.u_wallace._1021_ ;
 wire \u_cpu.ALU.u_wallace._1022_ ;
 wire \u_cpu.ALU.u_wallace._1023_ ;
 wire \u_cpu.ALU.u_wallace._1024_ ;
 wire \u_cpu.ALU.u_wallace._1025_ ;
 wire \u_cpu.ALU.u_wallace._1026_ ;
 wire \u_cpu.ALU.u_wallace._1027_ ;
 wire \u_cpu.ALU.u_wallace._1028_ ;
 wire \u_cpu.ALU.u_wallace._1029_ ;
 wire \u_cpu.ALU.u_wallace._1030_ ;
 wire \u_cpu.ALU.u_wallace._1031_ ;
 wire \u_cpu.ALU.u_wallace._1032_ ;
 wire \u_cpu.ALU.u_wallace._1033_ ;
 wire \u_cpu.ALU.u_wallace._1034_ ;
 wire \u_cpu.ALU.u_wallace._1035_ ;
 wire \u_cpu.ALU.u_wallace._1036_ ;
 wire \u_cpu.ALU.u_wallace._1037_ ;
 wire \u_cpu.ALU.u_wallace._1038_ ;
 wire \u_cpu.ALU.u_wallace._1039_ ;
 wire \u_cpu.ALU.u_wallace._1040_ ;
 wire \u_cpu.ALU.u_wallace._1041_ ;
 wire \u_cpu.ALU.u_wallace._1042_ ;
 wire \u_cpu.ALU.u_wallace._1043_ ;
 wire \u_cpu.ALU.u_wallace._1044_ ;
 wire \u_cpu.ALU.u_wallace._1045_ ;
 wire \u_cpu.ALU.u_wallace._1046_ ;
 wire \u_cpu.ALU.u_wallace._1047_ ;
 wire \u_cpu.ALU.u_wallace._1048_ ;
 wire \u_cpu.ALU.u_wallace._1049_ ;
 wire \u_cpu.ALU.u_wallace._1050_ ;
 wire \u_cpu.ALU.u_wallace._1051_ ;
 wire \u_cpu.ALU.u_wallace._1052_ ;
 wire \u_cpu.ALU.u_wallace._1053_ ;
 wire \u_cpu.ALU.u_wallace._1054_ ;
 wire \u_cpu.ALU.u_wallace._1055_ ;
 wire \u_cpu.ALU.u_wallace._1056_ ;
 wire \u_cpu.ALU.u_wallace._1057_ ;
 wire \u_cpu.ALU.u_wallace._1058_ ;
 wire \u_cpu.ALU.u_wallace._1059_ ;
 wire \u_cpu.ALU.u_wallace._1060_ ;
 wire \u_cpu.ALU.u_wallace._1061_ ;
 wire \u_cpu.ALU.u_wallace._1062_ ;
 wire \u_cpu.ALU.u_wallace._1063_ ;
 wire \u_cpu.ALU.u_wallace._1064_ ;
 wire \u_cpu.ALU.u_wallace._1065_ ;
 wire \u_cpu.ALU.u_wallace._1066_ ;
 wire \u_cpu.ALU.u_wallace._1067_ ;
 wire \u_cpu.ALU.u_wallace._1068_ ;
 wire \u_cpu.ALU.u_wallace._1069_ ;
 wire \u_cpu.ALU.u_wallace._1070_ ;
 wire \u_cpu.ALU.u_wallace._1071_ ;
 wire \u_cpu.ALU.u_wallace._1072_ ;
 wire \u_cpu.ALU.u_wallace._1073_ ;
 wire \u_cpu.ALU.u_wallace._1074_ ;
 wire \u_cpu.ALU.u_wallace._1075_ ;
 wire \u_cpu.ALU.u_wallace._1076_ ;
 wire \u_cpu.ALU.u_wallace._1077_ ;
 wire \u_cpu.ALU.u_wallace._1078_ ;
 wire \u_cpu.ALU.u_wallace._1079_ ;
 wire \u_cpu.ALU.u_wallace._1080_ ;
 wire \u_cpu.ALU.u_wallace._1081_ ;
 wire \u_cpu.ALU.u_wallace._1082_ ;
 wire \u_cpu.ALU.u_wallace._1083_ ;
 wire \u_cpu.ALU.u_wallace._1084_ ;
 wire \u_cpu.ALU.u_wallace._1085_ ;
 wire \u_cpu.ALU.u_wallace._1086_ ;
 wire \u_cpu.ALU.u_wallace._1087_ ;
 wire \u_cpu.ALU.u_wallace._1088_ ;
 wire \u_cpu.ALU.u_wallace._1089_ ;
 wire \u_cpu.ALU.u_wallace._1090_ ;
 wire \u_cpu.ALU.u_wallace._1091_ ;
 wire \u_cpu.ALU.u_wallace._1092_ ;
 wire \u_cpu.ALU.u_wallace._1093_ ;
 wire \u_cpu.ALU.u_wallace._1094_ ;
 wire \u_cpu.ALU.u_wallace._1095_ ;
 wire \u_cpu.ALU.u_wallace._1096_ ;
 wire \u_cpu.ALU.u_wallace._1097_ ;
 wire \u_cpu.ALU.u_wallace._1098_ ;
 wire \u_cpu.ALU.u_wallace._1099_ ;
 wire \u_cpu.ALU.u_wallace._1100_ ;
 wire \u_cpu.ALU.u_wallace._1101_ ;
 wire \u_cpu.ALU.u_wallace._1102_ ;
 wire \u_cpu.ALU.u_wallace._1103_ ;
 wire \u_cpu.ALU.u_wallace._1104_ ;
 wire \u_cpu.ALU.u_wallace._1105_ ;
 wire \u_cpu.ALU.u_wallace._1106_ ;
 wire \u_cpu.ALU.u_wallace._1107_ ;
 wire \u_cpu.ALU.u_wallace._1108_ ;
 wire \u_cpu.ALU.u_wallace._1109_ ;
 wire \u_cpu.ALU.u_wallace._1110_ ;
 wire \u_cpu.ALU.u_wallace._1111_ ;
 wire \u_cpu.ALU.u_wallace._1112_ ;
 wire \u_cpu.ALU.u_wallace._1113_ ;
 wire \u_cpu.ALU.u_wallace._1114_ ;
 wire \u_cpu.ALU.u_wallace._1115_ ;
 wire \u_cpu.ALU.u_wallace._1116_ ;
 wire \u_cpu.ALU.u_wallace._1117_ ;
 wire \u_cpu.ALU.u_wallace._1118_ ;
 wire \u_cpu.ALU.u_wallace._1119_ ;
 wire \u_cpu.ALU.u_wallace._1120_ ;
 wire \u_cpu.ALU.u_wallace._1121_ ;
 wire \u_cpu.ALU.u_wallace._1122_ ;
 wire \u_cpu.ALU.u_wallace._1123_ ;
 wire \u_cpu.ALU.u_wallace._1124_ ;
 wire \u_cpu.ALU.u_wallace._1125_ ;
 wire \u_cpu.ALU.u_wallace._1126_ ;
 wire \u_cpu.ALU.u_wallace._1127_ ;
 wire \u_cpu.ALU.u_wallace._1128_ ;
 wire \u_cpu.ALU.u_wallace._1129_ ;
 wire \u_cpu.ALU.u_wallace._1130_ ;
 wire \u_cpu.ALU.u_wallace._1131_ ;
 wire \u_cpu.ALU.u_wallace._1132_ ;
 wire \u_cpu.ALU.u_wallace._1133_ ;
 wire \u_cpu.ALU.u_wallace._1134_ ;
 wire \u_cpu.ALU.u_wallace._1135_ ;
 wire \u_cpu.ALU.u_wallace._1136_ ;
 wire \u_cpu.ALU.u_wallace._1137_ ;
 wire \u_cpu.ALU.u_wallace._1138_ ;
 wire \u_cpu.ALU.u_wallace._1139_ ;
 wire \u_cpu.ALU.u_wallace._1140_ ;
 wire \u_cpu.ALU.u_wallace._1141_ ;
 wire \u_cpu.ALU.u_wallace._1142_ ;
 wire \u_cpu.ALU.u_wallace._1143_ ;
 wire \u_cpu.ALU.u_wallace._1144_ ;
 wire \u_cpu.ALU.u_wallace._1145_ ;
 wire \u_cpu.ALU.u_wallace._1146_ ;
 wire \u_cpu.ALU.u_wallace._1147_ ;
 wire \u_cpu.ALU.u_wallace._1148_ ;
 wire \u_cpu.ALU.u_wallace._1149_ ;
 wire \u_cpu.ALU.u_wallace._1150_ ;
 wire \u_cpu.ALU.u_wallace._1151_ ;
 wire \u_cpu.ALU.u_wallace._1152_ ;
 wire \u_cpu.ALU.u_wallace._1153_ ;
 wire \u_cpu.ALU.u_wallace._1154_ ;
 wire \u_cpu.ALU.u_wallace._1155_ ;
 wire \u_cpu.ALU.u_wallace._1156_ ;
 wire \u_cpu.ALU.u_wallace._1157_ ;
 wire \u_cpu.ALU.u_wallace._1158_ ;
 wire \u_cpu.ALU.u_wallace._1159_ ;
 wire \u_cpu.ALU.u_wallace._1160_ ;
 wire \u_cpu.ALU.u_wallace._1161_ ;
 wire \u_cpu.ALU.u_wallace._1162_ ;
 wire \u_cpu.ALU.u_wallace._1163_ ;
 wire \u_cpu.ALU.u_wallace._1164_ ;
 wire \u_cpu.ALU.u_wallace._1165_ ;
 wire \u_cpu.ALU.u_wallace._1166_ ;
 wire \u_cpu.ALU.u_wallace._1167_ ;
 wire \u_cpu.ALU.u_wallace._1168_ ;
 wire \u_cpu.ALU.u_wallace._1169_ ;
 wire \u_cpu.ALU.u_wallace._1170_ ;
 wire \u_cpu.ALU.u_wallace._1171_ ;
 wire \u_cpu.ALU.u_wallace._1172_ ;
 wire \u_cpu.ALU.u_wallace._1173_ ;
 wire \u_cpu.ALU.u_wallace._1174_ ;
 wire \u_cpu.ALU.u_wallace._1175_ ;
 wire \u_cpu.ALU.u_wallace._1176_ ;
 wire \u_cpu.ALU.u_wallace._1177_ ;
 wire \u_cpu.ALU.u_wallace._1178_ ;
 wire \u_cpu.ALU.u_wallace._1179_ ;
 wire \u_cpu.ALU.u_wallace._1180_ ;
 wire \u_cpu.ALU.u_wallace._1181_ ;
 wire \u_cpu.ALU.u_wallace._1182_ ;
 wire \u_cpu.ALU.u_wallace._1183_ ;
 wire \u_cpu.ALU.u_wallace._1184_ ;
 wire \u_cpu.ALU.u_wallace._1185_ ;
 wire \u_cpu.ALU.u_wallace._1186_ ;
 wire \u_cpu.ALU.u_wallace._1187_ ;
 wire \u_cpu.ALU.u_wallace._1188_ ;
 wire \u_cpu.ALU.u_wallace._1189_ ;
 wire \u_cpu.ALU.u_wallace._1190_ ;
 wire \u_cpu.ALU.u_wallace._1191_ ;
 wire \u_cpu.ALU.u_wallace._1192_ ;
 wire \u_cpu.ALU.u_wallace._1193_ ;
 wire \u_cpu.ALU.u_wallace._1194_ ;
 wire \u_cpu.ALU.u_wallace._1195_ ;
 wire \u_cpu.ALU.u_wallace._1196_ ;
 wire \u_cpu.ALU.u_wallace._1197_ ;
 wire \u_cpu.ALU.u_wallace._1198_ ;
 wire \u_cpu.ALU.u_wallace._1199_ ;
 wire \u_cpu.ALU.u_wallace._1200_ ;
 wire \u_cpu.ALU.u_wallace._1201_ ;
 wire \u_cpu.ALU.u_wallace._1202_ ;
 wire \u_cpu.ALU.u_wallace._1203_ ;
 wire \u_cpu.ALU.u_wallace._1204_ ;
 wire \u_cpu.ALU.u_wallace._1205_ ;
 wire \u_cpu.ALU.u_wallace._1206_ ;
 wire \u_cpu.ALU.u_wallace._1207_ ;
 wire \u_cpu.ALU.u_wallace._1208_ ;
 wire \u_cpu.ALU.u_wallace._1209_ ;
 wire \u_cpu.ALU.u_wallace._1210_ ;
 wire \u_cpu.ALU.u_wallace._1211_ ;
 wire \u_cpu.ALU.u_wallace._1212_ ;
 wire \u_cpu.ALU.u_wallace._1213_ ;
 wire \u_cpu.ALU.u_wallace._1214_ ;
 wire \u_cpu.ALU.u_wallace._1215_ ;
 wire \u_cpu.ALU.u_wallace._1216_ ;
 wire \u_cpu.ALU.u_wallace._1217_ ;
 wire \u_cpu.ALU.u_wallace._1218_ ;
 wire \u_cpu.ALU.u_wallace._1219_ ;
 wire \u_cpu.ALU.u_wallace._1220_ ;
 wire \u_cpu.ALU.u_wallace._1221_ ;
 wire \u_cpu.ALU.u_wallace._1222_ ;
 wire \u_cpu.ALU.u_wallace._1223_ ;
 wire \u_cpu.ALU.u_wallace._1224_ ;
 wire \u_cpu.ALU.u_wallace._1225_ ;
 wire \u_cpu.ALU.u_wallace._1226_ ;
 wire \u_cpu.ALU.u_wallace._1227_ ;
 wire \u_cpu.ALU.u_wallace._1228_ ;
 wire \u_cpu.ALU.u_wallace._1229_ ;
 wire \u_cpu.ALU.u_wallace._1230_ ;
 wire \u_cpu.ALU.u_wallace._1231_ ;
 wire \u_cpu.ALU.u_wallace._1232_ ;
 wire \u_cpu.ALU.u_wallace._1233_ ;
 wire \u_cpu.ALU.u_wallace._1234_ ;
 wire \u_cpu.ALU.u_wallace._1235_ ;
 wire \u_cpu.ALU.u_wallace._1236_ ;
 wire \u_cpu.ALU.u_wallace._1237_ ;
 wire \u_cpu.ALU.u_wallace._1238_ ;
 wire \u_cpu.ALU.u_wallace._1239_ ;
 wire \u_cpu.ALU.u_wallace._1240_ ;
 wire \u_cpu.ALU.u_wallace._1241_ ;
 wire \u_cpu.ALU.u_wallace._1242_ ;
 wire \u_cpu.ALU.u_wallace._1243_ ;
 wire \u_cpu.ALU.u_wallace._1244_ ;
 wire \u_cpu.ALU.u_wallace._1245_ ;
 wire \u_cpu.ALU.u_wallace._1246_ ;
 wire \u_cpu.ALU.u_wallace._1247_ ;
 wire \u_cpu.ALU.u_wallace._1248_ ;
 wire \u_cpu.ALU.u_wallace._1249_ ;
 wire \u_cpu.ALU.u_wallace._1250_ ;
 wire \u_cpu.ALU.u_wallace._1251_ ;
 wire \u_cpu.ALU.u_wallace._1252_ ;
 wire \u_cpu.ALU.u_wallace._1253_ ;
 wire \u_cpu.ALU.u_wallace._1254_ ;
 wire \u_cpu.ALU.u_wallace._1255_ ;
 wire \u_cpu.ALU.u_wallace._1256_ ;
 wire \u_cpu.ALU.u_wallace._1257_ ;
 wire \u_cpu.ALU.u_wallace._1258_ ;
 wire \u_cpu.ALU.u_wallace._1259_ ;
 wire \u_cpu.ALU.u_wallace._1260_ ;
 wire \u_cpu.ALU.u_wallace._1261_ ;
 wire \u_cpu.ALU.u_wallace._1262_ ;
 wire \u_cpu.ALU.u_wallace._1263_ ;
 wire \u_cpu.ALU.u_wallace._1264_ ;
 wire \u_cpu.ALU.u_wallace._1265_ ;
 wire \u_cpu.ALU.u_wallace._1266_ ;
 wire \u_cpu.ALU.u_wallace._1267_ ;
 wire \u_cpu.ALU.u_wallace._1268_ ;
 wire \u_cpu.ALU.u_wallace._1269_ ;
 wire \u_cpu.ALU.u_wallace._1270_ ;
 wire \u_cpu.ALU.u_wallace._1271_ ;
 wire \u_cpu.ALU.u_wallace._1272_ ;
 wire \u_cpu.ALU.u_wallace._1273_ ;
 wire \u_cpu.ALU.u_wallace._1274_ ;
 wire \u_cpu.ALU.u_wallace._1275_ ;
 wire \u_cpu.ALU.u_wallace._1276_ ;
 wire \u_cpu.ALU.u_wallace._1277_ ;
 wire \u_cpu.ALU.u_wallace._1278_ ;
 wire \u_cpu.ALU.u_wallace._1279_ ;
 wire \u_cpu.ALU.u_wallace._1280_ ;
 wire \u_cpu.ALU.u_wallace._1281_ ;
 wire \u_cpu.ALU.u_wallace._1282_ ;
 wire \u_cpu.ALU.u_wallace._1283_ ;
 wire \u_cpu.ALU.u_wallace._1284_ ;
 wire \u_cpu.ALU.u_wallace._1285_ ;
 wire \u_cpu.ALU.u_wallace._1286_ ;
 wire \u_cpu.ALU.u_wallace._1287_ ;
 wire \u_cpu.ALU.u_wallace._1288_ ;
 wire \u_cpu.ALU.u_wallace._1289_ ;
 wire \u_cpu.ALU.u_wallace._1290_ ;
 wire \u_cpu.ALU.u_wallace._1291_ ;
 wire \u_cpu.ALU.u_wallace._1292_ ;
 wire \u_cpu.ALU.u_wallace._1293_ ;
 wire \u_cpu.ALU.u_wallace._1294_ ;
 wire \u_cpu.ALU.u_wallace._1295_ ;
 wire \u_cpu.ALU.u_wallace._1296_ ;
 wire \u_cpu.ALU.u_wallace._1297_ ;
 wire \u_cpu.ALU.u_wallace._1298_ ;
 wire \u_cpu.ALU.u_wallace._1299_ ;
 wire \u_cpu.ALU.u_wallace._1300_ ;
 wire \u_cpu.ALU.u_wallace._1301_ ;
 wire \u_cpu.ALU.u_wallace._1302_ ;
 wire \u_cpu.ALU.u_wallace._1303_ ;
 wire \u_cpu.ALU.u_wallace._1304_ ;
 wire \u_cpu.ALU.u_wallace._1305_ ;
 wire \u_cpu.ALU.u_wallace._1306_ ;
 wire \u_cpu.ALU.u_wallace._1307_ ;
 wire \u_cpu.ALU.u_wallace._1308_ ;
 wire \u_cpu.ALU.u_wallace._1309_ ;
 wire \u_cpu.ALU.u_wallace._1310_ ;
 wire \u_cpu.ALU.u_wallace._1311_ ;
 wire \u_cpu.ALU.u_wallace._1312_ ;
 wire \u_cpu.ALU.u_wallace._1313_ ;
 wire \u_cpu.ALU.u_wallace._1314_ ;
 wire \u_cpu.ALU.u_wallace._1315_ ;
 wire \u_cpu.ALU.u_wallace._1316_ ;
 wire \u_cpu.ALU.u_wallace._1317_ ;
 wire \u_cpu.ALU.u_wallace._1318_ ;
 wire \u_cpu.ALU.u_wallace._1319_ ;
 wire \u_cpu.ALU.u_wallace._1320_ ;
 wire \u_cpu.ALU.u_wallace._1321_ ;
 wire \u_cpu.ALU.u_wallace._1322_ ;
 wire \u_cpu.ALU.u_wallace._1323_ ;
 wire \u_cpu.ALU.u_wallace._1324_ ;
 wire \u_cpu.ALU.u_wallace._1325_ ;
 wire \u_cpu.ALU.u_wallace._1326_ ;
 wire \u_cpu.ALU.u_wallace._1327_ ;
 wire \u_cpu.ALU.u_wallace._1328_ ;
 wire \u_cpu.ALU.u_wallace._1329_ ;
 wire \u_cpu.ALU.u_wallace._1330_ ;
 wire \u_cpu.ALU.u_wallace._1331_ ;
 wire \u_cpu.ALU.u_wallace._1332_ ;
 wire \u_cpu.ALU.u_wallace._1333_ ;
 wire \u_cpu.ALU.u_wallace._1334_ ;
 wire \u_cpu.ALU.u_wallace._1335_ ;
 wire \u_cpu.ALU.u_wallace._1336_ ;
 wire \u_cpu.ALU.u_wallace._1337_ ;
 wire \u_cpu.ALU.u_wallace._1338_ ;
 wire \u_cpu.ALU.u_wallace._1339_ ;
 wire \u_cpu.ALU.u_wallace._1340_ ;
 wire \u_cpu.ALU.u_wallace._1341_ ;
 wire \u_cpu.ALU.u_wallace._1342_ ;
 wire \u_cpu.ALU.u_wallace._1343_ ;
 wire \u_cpu.ALU.u_wallace._1344_ ;
 wire \u_cpu.ALU.u_wallace._1345_ ;
 wire \u_cpu.ALU.u_wallace._1346_ ;
 wire \u_cpu.ALU.u_wallace._1347_ ;
 wire \u_cpu.ALU.u_wallace._1348_ ;
 wire \u_cpu.ALU.u_wallace._1349_ ;
 wire \u_cpu.ALU.u_wallace._1350_ ;
 wire \u_cpu.ALU.u_wallace._1351_ ;
 wire \u_cpu.ALU.u_wallace._1352_ ;
 wire \u_cpu.ALU.u_wallace._1353_ ;
 wire \u_cpu.ALU.u_wallace._1354_ ;
 wire \u_cpu.ALU.u_wallace._1355_ ;
 wire \u_cpu.ALU.u_wallace._1356_ ;
 wire \u_cpu.ALU.u_wallace._1357_ ;
 wire \u_cpu.ALU.u_wallace._1358_ ;
 wire \u_cpu.ALU.u_wallace._1359_ ;
 wire \u_cpu.ALU.u_wallace._1360_ ;
 wire \u_cpu.ALU.u_wallace._1361_ ;
 wire \u_cpu.ALU.u_wallace._1362_ ;
 wire \u_cpu.ALU.u_wallace._1363_ ;
 wire \u_cpu.ALU.u_wallace._1364_ ;
 wire \u_cpu.ALU.u_wallace._1365_ ;
 wire \u_cpu.ALU.u_wallace._1366_ ;
 wire \u_cpu.ALU.u_wallace._1367_ ;
 wire \u_cpu.ALU.u_wallace._1368_ ;
 wire \u_cpu.ALU.u_wallace._1369_ ;
 wire \u_cpu.ALU.u_wallace._1370_ ;
 wire \u_cpu.ALU.u_wallace._1371_ ;
 wire \u_cpu.ALU.u_wallace._1372_ ;
 wire \u_cpu.ALU.u_wallace._1373_ ;
 wire \u_cpu.ALU.u_wallace._1374_ ;
 wire \u_cpu.ALU.u_wallace._1375_ ;
 wire \u_cpu.ALU.u_wallace._1376_ ;
 wire \u_cpu.ALU.u_wallace._1377_ ;
 wire \u_cpu.ALU.u_wallace._1378_ ;
 wire \u_cpu.ALU.u_wallace._1379_ ;
 wire \u_cpu.ALU.u_wallace._1380_ ;
 wire \u_cpu.ALU.u_wallace._1381_ ;
 wire \u_cpu.ALU.u_wallace._1382_ ;
 wire \u_cpu.ALU.u_wallace._1383_ ;
 wire \u_cpu.ALU.u_wallace._1384_ ;
 wire \u_cpu.ALU.u_wallace._1385_ ;
 wire \u_cpu.ALU.u_wallace._1386_ ;
 wire \u_cpu.ALU.u_wallace._1387_ ;
 wire \u_cpu.ALU.u_wallace._1388_ ;
 wire \u_cpu.ALU.u_wallace._1389_ ;
 wire \u_cpu.ALU.u_wallace._1390_ ;
 wire \u_cpu.ALU.u_wallace._1391_ ;
 wire \u_cpu.ALU.u_wallace._1392_ ;
 wire \u_cpu.ALU.u_wallace._1393_ ;
 wire \u_cpu.ALU.u_wallace._1394_ ;
 wire \u_cpu.ALU.u_wallace._1395_ ;
 wire \u_cpu.ALU.u_wallace._1396_ ;
 wire \u_cpu.ALU.u_wallace._1397_ ;
 wire \u_cpu.ALU.u_wallace._1398_ ;
 wire \u_cpu.ALU.u_wallace._1399_ ;
 wire \u_cpu.ALU.u_wallace._1400_ ;
 wire \u_cpu.ALU.u_wallace._1401_ ;
 wire \u_cpu.ALU.u_wallace._1402_ ;
 wire \u_cpu.ALU.u_wallace._1403_ ;
 wire \u_cpu.ALU.u_wallace._1404_ ;
 wire \u_cpu.ALU.u_wallace._1405_ ;
 wire \u_cpu.ALU.u_wallace._1406_ ;
 wire \u_cpu.ALU.u_wallace._1407_ ;
 wire \u_cpu.ALU.u_wallace._1408_ ;
 wire \u_cpu.ALU.u_wallace._1409_ ;
 wire \u_cpu.ALU.u_wallace._1410_ ;
 wire \u_cpu.ALU.u_wallace._1411_ ;
 wire \u_cpu.ALU.u_wallace._1412_ ;
 wire \u_cpu.ALU.u_wallace._1413_ ;
 wire \u_cpu.ALU.u_wallace._1414_ ;
 wire \u_cpu.ALU.u_wallace._1415_ ;
 wire \u_cpu.ALU.u_wallace._1416_ ;
 wire \u_cpu.ALU.u_wallace._1417_ ;
 wire \u_cpu.ALU.u_wallace._1418_ ;
 wire \u_cpu.ALU.u_wallace._1419_ ;
 wire \u_cpu.ALU.u_wallace._1420_ ;
 wire \u_cpu.ALU.u_wallace._1421_ ;
 wire \u_cpu.ALU.u_wallace._1422_ ;
 wire \u_cpu.ALU.u_wallace._1423_ ;
 wire \u_cpu.ALU.u_wallace._1424_ ;
 wire \u_cpu.ALU.u_wallace._1425_ ;
 wire \u_cpu.ALU.u_wallace._1426_ ;
 wire \u_cpu.ALU.u_wallace._1427_ ;
 wire \u_cpu.ALU.u_wallace._1428_ ;
 wire \u_cpu.ALU.u_wallace._1429_ ;
 wire \u_cpu.ALU.u_wallace._1430_ ;
 wire \u_cpu.ALU.u_wallace._1431_ ;
 wire \u_cpu.ALU.u_wallace._1432_ ;
 wire \u_cpu.ALU.u_wallace._1433_ ;
 wire \u_cpu.ALU.u_wallace._1434_ ;
 wire \u_cpu.ALU.u_wallace._1435_ ;
 wire \u_cpu.ALU.u_wallace._1436_ ;
 wire \u_cpu.ALU.u_wallace._1437_ ;
 wire \u_cpu.ALU.u_wallace._1438_ ;
 wire \u_cpu.ALU.u_wallace._1439_ ;
 wire \u_cpu.ALU.u_wallace._1440_ ;
 wire \u_cpu.ALU.u_wallace._1441_ ;
 wire \u_cpu.ALU.u_wallace._1442_ ;
 wire \u_cpu.ALU.u_wallace._1443_ ;
 wire \u_cpu.ALU.u_wallace._1444_ ;
 wire \u_cpu.ALU.u_wallace._1445_ ;
 wire \u_cpu.ALU.u_wallace._1446_ ;
 wire \u_cpu.ALU.u_wallace._1447_ ;
 wire \u_cpu.ALU.u_wallace._1448_ ;
 wire \u_cpu.ALU.u_wallace._1449_ ;
 wire \u_cpu.ALU.u_wallace._1450_ ;
 wire \u_cpu.ALU.u_wallace._1451_ ;
 wire \u_cpu.ALU.u_wallace._1452_ ;
 wire \u_cpu.ALU.u_wallace._1453_ ;
 wire \u_cpu.ALU.u_wallace._1454_ ;
 wire \u_cpu.ALU.u_wallace._1455_ ;
 wire \u_cpu.ALU.u_wallace._1456_ ;
 wire \u_cpu.ALU.u_wallace._1457_ ;
 wire \u_cpu.ALU.u_wallace._1458_ ;
 wire \u_cpu.ALU.u_wallace._1459_ ;
 wire \u_cpu.ALU.u_wallace._1460_ ;
 wire \u_cpu.ALU.u_wallace._1461_ ;
 wire \u_cpu.ALU.u_wallace._1462_ ;
 wire \u_cpu.ALU.u_wallace._1463_ ;
 wire \u_cpu.ALU.u_wallace._1464_ ;
 wire \u_cpu.ALU.u_wallace._1465_ ;
 wire \u_cpu.ALU.u_wallace._1466_ ;
 wire \u_cpu.ALU.u_wallace._1467_ ;
 wire \u_cpu.ALU.u_wallace._1468_ ;
 wire \u_cpu.ALU.u_wallace._1469_ ;
 wire \u_cpu.ALU.u_wallace._1470_ ;
 wire \u_cpu.ALU.u_wallace._1471_ ;
 wire \u_cpu.ALU.u_wallace._1472_ ;
 wire \u_cpu.ALU.u_wallace._1473_ ;
 wire \u_cpu.ALU.u_wallace._1474_ ;
 wire \u_cpu.ALU.u_wallace._1475_ ;
 wire \u_cpu.ALU.u_wallace._1476_ ;
 wire \u_cpu.ALU.u_wallace._1477_ ;
 wire \u_cpu.ALU.u_wallace._1478_ ;
 wire \u_cpu.ALU.u_wallace._1479_ ;
 wire \u_cpu.ALU.u_wallace._1480_ ;
 wire \u_cpu.ALU.u_wallace._1481_ ;
 wire \u_cpu.ALU.u_wallace._1482_ ;
 wire \u_cpu.ALU.u_wallace._1483_ ;
 wire \u_cpu.ALU.u_wallace._1484_ ;
 wire \u_cpu.ALU.u_wallace._1485_ ;
 wire \u_cpu.ALU.u_wallace._1486_ ;
 wire \u_cpu.ALU.u_wallace._1487_ ;
 wire \u_cpu.ALU.u_wallace._1488_ ;
 wire \u_cpu.ALU.u_wallace._1489_ ;
 wire \u_cpu.ALU.u_wallace._1490_ ;
 wire \u_cpu.ALU.u_wallace._1491_ ;
 wire \u_cpu.ALU.u_wallace._1492_ ;
 wire \u_cpu.ALU.u_wallace._1493_ ;
 wire \u_cpu.ALU.u_wallace._1494_ ;
 wire \u_cpu.ALU.u_wallace._1495_ ;
 wire \u_cpu.ALU.u_wallace._1496_ ;
 wire \u_cpu.ALU.u_wallace._1497_ ;
 wire \u_cpu.ALU.u_wallace._1498_ ;
 wire \u_cpu.ALU.u_wallace._1499_ ;
 wire \u_cpu.ALU.u_wallace._1500_ ;
 wire \u_cpu.ALU.u_wallace._1501_ ;
 wire \u_cpu.ALU.u_wallace._1502_ ;
 wire \u_cpu.ALU.u_wallace._1503_ ;
 wire \u_cpu.ALU.u_wallace._1504_ ;
 wire \u_cpu.ALU.u_wallace._1505_ ;
 wire \u_cpu.ALU.u_wallace._1506_ ;
 wire \u_cpu.ALU.u_wallace._1507_ ;
 wire \u_cpu.ALU.u_wallace._1508_ ;
 wire \u_cpu.ALU.u_wallace._1509_ ;
 wire \u_cpu.ALU.u_wallace._1510_ ;
 wire \u_cpu.ALU.u_wallace._1511_ ;
 wire \u_cpu.ALU.u_wallace._1512_ ;
 wire \u_cpu.ALU.u_wallace._1513_ ;
 wire \u_cpu.ALU.u_wallace._1514_ ;
 wire \u_cpu.ALU.u_wallace._1515_ ;
 wire \u_cpu.ALU.u_wallace._1516_ ;
 wire \u_cpu.ALU.u_wallace._1517_ ;
 wire \u_cpu.ALU.u_wallace._1518_ ;
 wire \u_cpu.ALU.u_wallace._1519_ ;
 wire \u_cpu.ALU.u_wallace._1520_ ;
 wire \u_cpu.ALU.u_wallace._1521_ ;
 wire \u_cpu.ALU.u_wallace._1522_ ;
 wire \u_cpu.ALU.u_wallace._1523_ ;
 wire \u_cpu.ALU.u_wallace._1524_ ;
 wire \u_cpu.ALU.u_wallace._1525_ ;
 wire \u_cpu.ALU.u_wallace._1526_ ;
 wire \u_cpu.ALU.u_wallace._1527_ ;
 wire \u_cpu.ALU.u_wallace._1528_ ;
 wire \u_cpu.ALU.u_wallace._1529_ ;
 wire \u_cpu.ALU.u_wallace._1530_ ;
 wire \u_cpu.ALU.u_wallace._1531_ ;
 wire \u_cpu.ALU.u_wallace._1532_ ;
 wire \u_cpu.ALU.u_wallace._1533_ ;
 wire \u_cpu.ALU.u_wallace._1534_ ;
 wire \u_cpu.ALU.u_wallace._1535_ ;
 wire \u_cpu.ALU.u_wallace._1536_ ;
 wire \u_cpu.ALU.u_wallace._1537_ ;
 wire \u_cpu.ALU.u_wallace._1538_ ;
 wire \u_cpu.ALU.u_wallace._1539_ ;
 wire \u_cpu.ALU.u_wallace._1540_ ;
 wire \u_cpu.ALU.u_wallace._1541_ ;
 wire \u_cpu.ALU.u_wallace._1542_ ;
 wire \u_cpu.ALU.u_wallace._1543_ ;
 wire \u_cpu.ALU.u_wallace._1544_ ;
 wire \u_cpu.ALU.u_wallace._1545_ ;
 wire \u_cpu.ALU.u_wallace._1546_ ;
 wire \u_cpu.ALU.u_wallace._1547_ ;
 wire \u_cpu.ALU.u_wallace._1548_ ;
 wire \u_cpu.ALU.u_wallace._1549_ ;
 wire \u_cpu.ALU.u_wallace._1550_ ;
 wire \u_cpu.ALU.u_wallace._1551_ ;
 wire \u_cpu.ALU.u_wallace._1552_ ;
 wire \u_cpu.ALU.u_wallace._1553_ ;
 wire \u_cpu.ALU.u_wallace._1554_ ;
 wire \u_cpu.ALU.u_wallace._1555_ ;
 wire \u_cpu.ALU.u_wallace._1556_ ;
 wire \u_cpu.ALU.u_wallace._1557_ ;
 wire \u_cpu.ALU.u_wallace._1558_ ;
 wire \u_cpu.ALU.u_wallace._1559_ ;
 wire \u_cpu.ALU.u_wallace._1560_ ;
 wire \u_cpu.ALU.u_wallace._1561_ ;
 wire \u_cpu.ALU.u_wallace._1562_ ;
 wire \u_cpu.ALU.u_wallace._1563_ ;
 wire \u_cpu.ALU.u_wallace._1564_ ;
 wire \u_cpu.ALU.u_wallace._1565_ ;
 wire \u_cpu.ALU.u_wallace._1566_ ;
 wire \u_cpu.ALU.u_wallace._1567_ ;
 wire \u_cpu.ALU.u_wallace._1568_ ;
 wire \u_cpu.ALU.u_wallace._1569_ ;
 wire \u_cpu.ALU.u_wallace._1570_ ;
 wire \u_cpu.ALU.u_wallace._1571_ ;
 wire \u_cpu.ALU.u_wallace._1572_ ;
 wire \u_cpu.ALU.u_wallace._1573_ ;
 wire \u_cpu.ALU.u_wallace._1574_ ;
 wire \u_cpu.ALU.u_wallace._1575_ ;
 wire \u_cpu.ALU.u_wallace._1576_ ;
 wire \u_cpu.ALU.u_wallace._1577_ ;
 wire \u_cpu.ALU.u_wallace._1578_ ;
 wire \u_cpu.ALU.u_wallace._1579_ ;
 wire \u_cpu.ALU.u_wallace._1580_ ;
 wire \u_cpu.ALU.u_wallace._1581_ ;
 wire \u_cpu.ALU.u_wallace._1582_ ;
 wire \u_cpu.ALU.u_wallace._1583_ ;
 wire \u_cpu.ALU.u_wallace._1584_ ;
 wire \u_cpu.ALU.u_wallace._1585_ ;
 wire \u_cpu.ALU.u_wallace._1586_ ;
 wire \u_cpu.ALU.u_wallace._1587_ ;
 wire \u_cpu.ALU.u_wallace._1588_ ;
 wire \u_cpu.ALU.u_wallace._1589_ ;
 wire \u_cpu.ALU.u_wallace._1590_ ;
 wire \u_cpu.ALU.u_wallace._1591_ ;
 wire \u_cpu.ALU.u_wallace._1592_ ;
 wire \u_cpu.ALU.u_wallace._1593_ ;
 wire \u_cpu.ALU.u_wallace._1594_ ;
 wire \u_cpu.ALU.u_wallace._1595_ ;
 wire \u_cpu.ALU.u_wallace._1596_ ;
 wire \u_cpu.ALU.u_wallace._1597_ ;
 wire \u_cpu.ALU.u_wallace._1598_ ;
 wire \u_cpu.ALU.u_wallace._1599_ ;
 wire \u_cpu.ALU.u_wallace._1600_ ;
 wire \u_cpu.ALU.u_wallace._1601_ ;
 wire \u_cpu.ALU.u_wallace._1602_ ;
 wire \u_cpu.ALU.u_wallace._1603_ ;
 wire \u_cpu.ALU.u_wallace._1604_ ;
 wire \u_cpu.ALU.u_wallace._1605_ ;
 wire \u_cpu.ALU.u_wallace._1606_ ;
 wire \u_cpu.ALU.u_wallace._1607_ ;
 wire \u_cpu.ALU.u_wallace._1608_ ;
 wire \u_cpu.ALU.u_wallace._1609_ ;
 wire \u_cpu.ALU.u_wallace._1610_ ;
 wire \u_cpu.ALU.u_wallace._1611_ ;
 wire \u_cpu.ALU.u_wallace._1612_ ;
 wire \u_cpu.ALU.u_wallace._1613_ ;
 wire \u_cpu.ALU.u_wallace._1614_ ;
 wire \u_cpu.ALU.u_wallace._1615_ ;
 wire \u_cpu.ALU.u_wallace._1616_ ;
 wire \u_cpu.ALU.u_wallace._1617_ ;
 wire \u_cpu.ALU.u_wallace._1618_ ;
 wire \u_cpu.ALU.u_wallace._1619_ ;
 wire \u_cpu.ALU.u_wallace._1620_ ;
 wire \u_cpu.ALU.u_wallace._1621_ ;
 wire \u_cpu.ALU.u_wallace._1622_ ;
 wire \u_cpu.ALU.u_wallace._1623_ ;
 wire \u_cpu.ALU.u_wallace._1624_ ;
 wire \u_cpu.ALU.u_wallace._1625_ ;
 wire \u_cpu.ALU.u_wallace._1626_ ;
 wire \u_cpu.ALU.u_wallace._1627_ ;
 wire \u_cpu.ALU.u_wallace._1628_ ;
 wire \u_cpu.ALU.u_wallace._1629_ ;
 wire \u_cpu.ALU.u_wallace._1630_ ;
 wire \u_cpu.ALU.u_wallace._1631_ ;
 wire \u_cpu.ALU.u_wallace._1632_ ;
 wire \u_cpu.ALU.u_wallace._1633_ ;
 wire \u_cpu.ALU.u_wallace._1634_ ;
 wire \u_cpu.ALU.u_wallace._1635_ ;
 wire \u_cpu.ALU.u_wallace._1636_ ;
 wire \u_cpu.ALU.u_wallace._1637_ ;
 wire \u_cpu.ALU.u_wallace._1638_ ;
 wire \u_cpu.ALU.u_wallace._1639_ ;
 wire \u_cpu.ALU.u_wallace._1640_ ;
 wire \u_cpu.ALU.u_wallace._1641_ ;
 wire \u_cpu.ALU.u_wallace._1642_ ;
 wire \u_cpu.ALU.u_wallace._1643_ ;
 wire \u_cpu.ALU.u_wallace._1644_ ;
 wire \u_cpu.ALU.u_wallace._1645_ ;
 wire \u_cpu.ALU.u_wallace._1646_ ;
 wire \u_cpu.ALU.u_wallace._1647_ ;
 wire \u_cpu.ALU.u_wallace._1648_ ;
 wire \u_cpu.ALU.u_wallace._1649_ ;
 wire \u_cpu.ALU.u_wallace._1650_ ;
 wire \u_cpu.ALU.u_wallace._1651_ ;
 wire \u_cpu.ALU.u_wallace._1652_ ;
 wire \u_cpu.ALU.u_wallace._1653_ ;
 wire \u_cpu.ALU.u_wallace._1654_ ;
 wire \u_cpu.ALU.u_wallace._1655_ ;
 wire \u_cpu.ALU.u_wallace._1656_ ;
 wire \u_cpu.ALU.u_wallace._1657_ ;
 wire \u_cpu.ALU.u_wallace._1658_ ;
 wire \u_cpu.ALU.u_wallace._1659_ ;
 wire \u_cpu.ALU.u_wallace._1660_ ;
 wire \u_cpu.ALU.u_wallace._1661_ ;
 wire \u_cpu.ALU.u_wallace._1662_ ;
 wire \u_cpu.ALU.u_wallace._1663_ ;
 wire \u_cpu.ALU.u_wallace._1664_ ;
 wire \u_cpu.ALU.u_wallace._1665_ ;
 wire \u_cpu.ALU.u_wallace._1666_ ;
 wire \u_cpu.ALU.u_wallace._1667_ ;
 wire \u_cpu.ALU.u_wallace._1668_ ;
 wire \u_cpu.ALU.u_wallace._1669_ ;
 wire \u_cpu.ALU.u_wallace._1670_ ;
 wire \u_cpu.ALU.u_wallace._1671_ ;
 wire \u_cpu.ALU.u_wallace._1672_ ;
 wire \u_cpu.ALU.u_wallace._1673_ ;
 wire \u_cpu.ALU.u_wallace._1674_ ;
 wire \u_cpu.ALU.u_wallace._1675_ ;
 wire \u_cpu.ALU.u_wallace._1676_ ;
 wire \u_cpu.ALU.u_wallace._1677_ ;
 wire \u_cpu.ALU.u_wallace._1678_ ;
 wire \u_cpu.ALU.u_wallace._1679_ ;
 wire \u_cpu.ALU.u_wallace._1680_ ;
 wire \u_cpu.ALU.u_wallace._1681_ ;
 wire \u_cpu.ALU.u_wallace._1682_ ;
 wire \u_cpu.ALU.u_wallace._1683_ ;
 wire \u_cpu.ALU.u_wallace._1684_ ;
 wire \u_cpu.ALU.u_wallace._1685_ ;
 wire \u_cpu.ALU.u_wallace._1686_ ;
 wire \u_cpu.ALU.u_wallace._1687_ ;
 wire \u_cpu.ALU.u_wallace._1688_ ;
 wire \u_cpu.ALU.u_wallace._1689_ ;
 wire \u_cpu.ALU.u_wallace._1690_ ;
 wire \u_cpu.ALU.u_wallace._1691_ ;
 wire \u_cpu.ALU.u_wallace._1692_ ;
 wire \u_cpu.ALU.u_wallace._1693_ ;
 wire \u_cpu.ALU.u_wallace._1694_ ;
 wire \u_cpu.ALU.u_wallace._1695_ ;
 wire \u_cpu.ALU.u_wallace._1696_ ;
 wire \u_cpu.ALU.u_wallace._1697_ ;
 wire \u_cpu.ALU.u_wallace._1698_ ;
 wire \u_cpu.ALU.u_wallace._1699_ ;
 wire \u_cpu.ALU.u_wallace._1700_ ;
 wire \u_cpu.ALU.u_wallace._1701_ ;
 wire \u_cpu.ALU.u_wallace._1702_ ;
 wire \u_cpu.ALU.u_wallace._1703_ ;
 wire \u_cpu.ALU.u_wallace._1704_ ;
 wire \u_cpu.ALU.u_wallace._1705_ ;
 wire \u_cpu.ALU.u_wallace._1706_ ;
 wire \u_cpu.ALU.u_wallace._1707_ ;
 wire \u_cpu.ALU.u_wallace._1708_ ;
 wire \u_cpu.ALU.u_wallace._1709_ ;
 wire \u_cpu.ALU.u_wallace._1710_ ;
 wire \u_cpu.ALU.u_wallace._1711_ ;
 wire \u_cpu.ALU.u_wallace._1712_ ;
 wire \u_cpu.ALU.u_wallace._1713_ ;
 wire \u_cpu.ALU.u_wallace._1714_ ;
 wire \u_cpu.ALU.u_wallace._1715_ ;
 wire \u_cpu.ALU.u_wallace._1716_ ;
 wire \u_cpu.ALU.u_wallace._1717_ ;
 wire \u_cpu.ALU.u_wallace._1718_ ;
 wire \u_cpu.ALU.u_wallace._1719_ ;
 wire \u_cpu.ALU.u_wallace._1720_ ;
 wire \u_cpu.ALU.u_wallace._1721_ ;
 wire \u_cpu.ALU.u_wallace._1722_ ;
 wire \u_cpu.ALU.u_wallace._1723_ ;
 wire \u_cpu.ALU.u_wallace._1724_ ;
 wire \u_cpu.ALU.u_wallace._1725_ ;
 wire \u_cpu.ALU.u_wallace._1726_ ;
 wire \u_cpu.ALU.u_wallace._1727_ ;
 wire \u_cpu.ALU.u_wallace._1728_ ;
 wire \u_cpu.ALU.u_wallace._1729_ ;
 wire \u_cpu.ALU.u_wallace._1730_ ;
 wire \u_cpu.ALU.u_wallace._1731_ ;
 wire \u_cpu.ALU.u_wallace._1732_ ;
 wire \u_cpu.ALU.u_wallace._1733_ ;
 wire \u_cpu.ALU.u_wallace._1734_ ;
 wire \u_cpu.ALU.u_wallace._1735_ ;
 wire \u_cpu.ALU.u_wallace._1736_ ;
 wire \u_cpu.ALU.u_wallace._1737_ ;
 wire \u_cpu.ALU.u_wallace._1738_ ;
 wire \u_cpu.ALU.u_wallace._1739_ ;
 wire \u_cpu.ALU.u_wallace._1740_ ;
 wire \u_cpu.ALU.u_wallace._1741_ ;
 wire \u_cpu.ALU.u_wallace._1742_ ;
 wire \u_cpu.ALU.u_wallace._1743_ ;
 wire \u_cpu.ALU.u_wallace._1744_ ;
 wire \u_cpu.ALU.u_wallace._1745_ ;
 wire \u_cpu.ALU.u_wallace._1746_ ;
 wire \u_cpu.ALU.u_wallace._1747_ ;
 wire \u_cpu.ALU.u_wallace._1748_ ;
 wire \u_cpu.ALU.u_wallace._1749_ ;
 wire \u_cpu.ALU.u_wallace._1750_ ;
 wire \u_cpu.ALU.u_wallace._1751_ ;
 wire \u_cpu.ALU.u_wallace._1752_ ;
 wire \u_cpu.ALU.u_wallace._1753_ ;
 wire \u_cpu.ALU.u_wallace._1754_ ;
 wire \u_cpu.ALU.u_wallace._1755_ ;
 wire \u_cpu.ALU.u_wallace._1756_ ;
 wire \u_cpu.ALU.u_wallace._1757_ ;
 wire \u_cpu.ALU.u_wallace._1758_ ;
 wire \u_cpu.ALU.u_wallace._1759_ ;
 wire \u_cpu.ALU.u_wallace._1760_ ;
 wire \u_cpu.ALU.u_wallace._1761_ ;
 wire \u_cpu.ALU.u_wallace._1762_ ;
 wire \u_cpu.ALU.u_wallace._1763_ ;
 wire \u_cpu.ALU.u_wallace._1764_ ;
 wire \u_cpu.ALU.u_wallace._1765_ ;
 wire \u_cpu.ALU.u_wallace._1766_ ;
 wire \u_cpu.ALU.u_wallace._1767_ ;
 wire \u_cpu.ALU.u_wallace._1768_ ;
 wire \u_cpu.ALU.u_wallace._1769_ ;
 wire \u_cpu.ALU.u_wallace._1770_ ;
 wire \u_cpu.ALU.u_wallace._1771_ ;
 wire \u_cpu.ALU.u_wallace._1772_ ;
 wire \u_cpu.ALU.u_wallace._1773_ ;
 wire \u_cpu.ALU.u_wallace._1774_ ;
 wire \u_cpu.ALU.u_wallace._1775_ ;
 wire \u_cpu.ALU.u_wallace._1776_ ;
 wire \u_cpu.ALU.u_wallace._1777_ ;
 wire \u_cpu.ALU.u_wallace._1778_ ;
 wire \u_cpu.ALU.u_wallace._1779_ ;
 wire \u_cpu.ALU.u_wallace._1780_ ;
 wire \u_cpu.ALU.u_wallace._1781_ ;
 wire \u_cpu.ALU.u_wallace._1782_ ;
 wire \u_cpu.ALU.u_wallace._1783_ ;
 wire \u_cpu.ALU.u_wallace._1784_ ;
 wire \u_cpu.ALU.u_wallace._1785_ ;
 wire \u_cpu.ALU.u_wallace._1786_ ;
 wire \u_cpu.ALU.u_wallace._1787_ ;
 wire \u_cpu.ALU.u_wallace._1788_ ;
 wire \u_cpu.ALU.u_wallace._1789_ ;
 wire \u_cpu.ALU.u_wallace._1790_ ;
 wire \u_cpu.ALU.u_wallace._1791_ ;
 wire \u_cpu.ALU.u_wallace._1792_ ;
 wire \u_cpu.ALU.u_wallace._1793_ ;
 wire \u_cpu.ALU.u_wallace._1794_ ;
 wire \u_cpu.ALU.u_wallace._1795_ ;
 wire \u_cpu.ALU.u_wallace._1796_ ;
 wire \u_cpu.ALU.u_wallace._1797_ ;
 wire \u_cpu.ALU.u_wallace._1798_ ;
 wire \u_cpu.ALU.u_wallace._1799_ ;
 wire \u_cpu.ALU.u_wallace._1800_ ;
 wire \u_cpu.ALU.u_wallace._1801_ ;
 wire \u_cpu.ALU.u_wallace._1802_ ;
 wire \u_cpu.ALU.u_wallace._1803_ ;
 wire \u_cpu.ALU.u_wallace._1804_ ;
 wire \u_cpu.ALU.u_wallace._1805_ ;
 wire \u_cpu.ALU.u_wallace._1806_ ;
 wire \u_cpu.ALU.u_wallace._1807_ ;
 wire \u_cpu.ALU.u_wallace._1808_ ;
 wire \u_cpu.ALU.u_wallace._1809_ ;
 wire \u_cpu.ALU.u_wallace._1810_ ;
 wire \u_cpu.ALU.u_wallace._1811_ ;
 wire \u_cpu.ALU.u_wallace._1812_ ;
 wire \u_cpu.ALU.u_wallace._1813_ ;
 wire \u_cpu.ALU.u_wallace._1814_ ;
 wire \u_cpu.ALU.u_wallace._1815_ ;
 wire \u_cpu.ALU.u_wallace._1816_ ;
 wire \u_cpu.ALU.u_wallace._1817_ ;
 wire \u_cpu.ALU.u_wallace._1818_ ;
 wire \u_cpu.ALU.u_wallace._1819_ ;
 wire \u_cpu.ALU.u_wallace._1820_ ;
 wire \u_cpu.ALU.u_wallace._1821_ ;
 wire \u_cpu.ALU.u_wallace._1822_ ;
 wire \u_cpu.ALU.u_wallace._1823_ ;
 wire \u_cpu.ALU.u_wallace._1824_ ;
 wire \u_cpu.ALU.u_wallace._1825_ ;
 wire \u_cpu.ALU.u_wallace._1826_ ;
 wire \u_cpu.ALU.u_wallace._1827_ ;
 wire \u_cpu.ALU.u_wallace._1828_ ;
 wire \u_cpu.ALU.u_wallace._1829_ ;
 wire \u_cpu.ALU.u_wallace._1830_ ;
 wire \u_cpu.ALU.u_wallace._1831_ ;
 wire \u_cpu.ALU.u_wallace._1832_ ;
 wire \u_cpu.ALU.u_wallace._1833_ ;
 wire \u_cpu.ALU.u_wallace._1834_ ;
 wire \u_cpu.ALU.u_wallace._1835_ ;
 wire \u_cpu.ALU.u_wallace._1836_ ;
 wire \u_cpu.ALU.u_wallace._1837_ ;
 wire \u_cpu.ALU.u_wallace._1838_ ;
 wire \u_cpu.ALU.u_wallace._1839_ ;
 wire \u_cpu.ALU.u_wallace._1840_ ;
 wire \u_cpu.ALU.u_wallace._1841_ ;
 wire \u_cpu.ALU.u_wallace._1842_ ;
 wire \u_cpu.ALU.u_wallace._1843_ ;
 wire \u_cpu.ALU.u_wallace._1844_ ;
 wire \u_cpu.ALU.u_wallace._1845_ ;
 wire \u_cpu.ALU.u_wallace._1846_ ;
 wire \u_cpu.ALU.u_wallace._1847_ ;
 wire \u_cpu.ALU.u_wallace._1848_ ;
 wire \u_cpu.ALU.u_wallace._1849_ ;
 wire \u_cpu.ALU.u_wallace._1850_ ;
 wire \u_cpu.ALU.u_wallace._1851_ ;
 wire \u_cpu.ALU.u_wallace._1852_ ;
 wire \u_cpu.ALU.u_wallace._1853_ ;
 wire \u_cpu.ALU.u_wallace._1854_ ;
 wire \u_cpu.ALU.u_wallace._1855_ ;
 wire \u_cpu.ALU.u_wallace._1856_ ;
 wire \u_cpu.ALU.u_wallace._1857_ ;
 wire \u_cpu.ALU.u_wallace._1858_ ;
 wire \u_cpu.ALU.u_wallace._1859_ ;
 wire \u_cpu.ALU.u_wallace._1860_ ;
 wire \u_cpu.ALU.u_wallace._1861_ ;
 wire \u_cpu.ALU.u_wallace._1862_ ;
 wire \u_cpu.ALU.u_wallace._1863_ ;
 wire \u_cpu.ALU.u_wallace._1864_ ;
 wire \u_cpu.ALU.u_wallace._1865_ ;
 wire \u_cpu.ALU.u_wallace._1866_ ;
 wire \u_cpu.ALU.u_wallace._1867_ ;
 wire \u_cpu.ALU.u_wallace._1868_ ;
 wire \u_cpu.ALU.u_wallace._1869_ ;
 wire \u_cpu.ALU.u_wallace._1870_ ;
 wire \u_cpu.ALU.u_wallace._1871_ ;
 wire \u_cpu.ALU.u_wallace._1872_ ;
 wire \u_cpu.ALU.u_wallace._1873_ ;
 wire \u_cpu.ALU.u_wallace._1874_ ;
 wire \u_cpu.ALU.u_wallace._1875_ ;
 wire \u_cpu.ALU.u_wallace._1876_ ;
 wire \u_cpu.ALU.u_wallace._1877_ ;
 wire \u_cpu.ALU.u_wallace._1878_ ;
 wire \u_cpu.ALU.u_wallace._1879_ ;
 wire \u_cpu.ALU.u_wallace._1880_ ;
 wire \u_cpu.ALU.u_wallace._1881_ ;
 wire \u_cpu.ALU.u_wallace._1882_ ;
 wire \u_cpu.ALU.u_wallace._1883_ ;
 wire \u_cpu.ALU.u_wallace._1884_ ;
 wire \u_cpu.ALU.u_wallace._1885_ ;
 wire \u_cpu.ALU.u_wallace._1886_ ;
 wire \u_cpu.ALU.u_wallace._1887_ ;
 wire \u_cpu.ALU.u_wallace._1888_ ;
 wire \u_cpu.ALU.u_wallace._1889_ ;
 wire \u_cpu.ALU.u_wallace._1890_ ;
 wire \u_cpu.ALU.u_wallace._1891_ ;
 wire \u_cpu.ALU.u_wallace._1892_ ;
 wire \u_cpu.ALU.u_wallace._1893_ ;
 wire \u_cpu.ALU.u_wallace._1894_ ;
 wire \u_cpu.ALU.u_wallace._1895_ ;
 wire \u_cpu.ALU.u_wallace._1896_ ;
 wire \u_cpu.ALU.u_wallace._1897_ ;
 wire \u_cpu.ALU.u_wallace._1898_ ;
 wire \u_cpu.ALU.u_wallace._1899_ ;
 wire \u_cpu.ALU.u_wallace._1900_ ;
 wire \u_cpu.ALU.u_wallace._1901_ ;
 wire \u_cpu.ALU.u_wallace._1902_ ;
 wire \u_cpu.ALU.u_wallace._1903_ ;
 wire \u_cpu.ALU.u_wallace._1904_ ;
 wire \u_cpu.ALU.u_wallace._1905_ ;
 wire \u_cpu.ALU.u_wallace._1906_ ;
 wire \u_cpu.ALU.u_wallace._1907_ ;
 wire \u_cpu.ALU.u_wallace._1908_ ;
 wire \u_cpu.ALU.u_wallace._1909_ ;
 wire \u_cpu.ALU.u_wallace._1910_ ;
 wire \u_cpu.ALU.u_wallace._1911_ ;
 wire \u_cpu.ALU.u_wallace._1912_ ;
 wire \u_cpu.ALU.u_wallace._1913_ ;
 wire \u_cpu.ALU.u_wallace._1914_ ;
 wire \u_cpu.ALU.u_wallace._1915_ ;
 wire \u_cpu.ALU.u_wallace._1916_ ;
 wire \u_cpu.ALU.u_wallace._1917_ ;
 wire \u_cpu.ALU.u_wallace._1918_ ;
 wire \u_cpu.ALU.u_wallace._1919_ ;
 wire \u_cpu.ALU.u_wallace._1920_ ;
 wire \u_cpu.ALU.u_wallace._1921_ ;
 wire \u_cpu.ALU.u_wallace._1922_ ;
 wire \u_cpu.ALU.u_wallace._1923_ ;
 wire \u_cpu.ALU.u_wallace._1924_ ;
 wire \u_cpu.ALU.u_wallace._1925_ ;
 wire \u_cpu.ALU.u_wallace._1926_ ;
 wire \u_cpu.ALU.u_wallace._1927_ ;
 wire \u_cpu.ALU.u_wallace._1928_ ;
 wire \u_cpu.ALU.u_wallace._1929_ ;
 wire \u_cpu.ALU.u_wallace._1930_ ;
 wire \u_cpu.ALU.u_wallace._1931_ ;
 wire \u_cpu.ALU.u_wallace._1932_ ;
 wire \u_cpu.ALU.u_wallace._1933_ ;
 wire \u_cpu.ALU.u_wallace._1934_ ;
 wire \u_cpu.ALU.u_wallace._1935_ ;
 wire \u_cpu.ALU.u_wallace._1936_ ;
 wire \u_cpu.ALU.u_wallace._1937_ ;
 wire \u_cpu.ALU.u_wallace._1938_ ;
 wire \u_cpu.ALU.u_wallace._1939_ ;
 wire \u_cpu.ALU.u_wallace._1940_ ;
 wire \u_cpu.ALU.u_wallace._1941_ ;
 wire \u_cpu.ALU.u_wallace._1942_ ;
 wire \u_cpu.ALU.u_wallace._1943_ ;
 wire \u_cpu.ALU.u_wallace._1944_ ;
 wire \u_cpu.ALU.u_wallace._1945_ ;
 wire \u_cpu.ALU.u_wallace._1946_ ;
 wire \u_cpu.ALU.u_wallace._1947_ ;
 wire \u_cpu.ALU.u_wallace._1948_ ;
 wire \u_cpu.ALU.u_wallace._1949_ ;
 wire \u_cpu.ALU.u_wallace._1950_ ;
 wire \u_cpu.ALU.u_wallace._1951_ ;
 wire \u_cpu.ALU.u_wallace._1952_ ;
 wire \u_cpu.ALU.u_wallace._1953_ ;
 wire \u_cpu.ALU.u_wallace._1954_ ;
 wire \u_cpu.ALU.u_wallace._1955_ ;
 wire \u_cpu.ALU.u_wallace._1956_ ;
 wire \u_cpu.ALU.u_wallace._1957_ ;
 wire \u_cpu.ALU.u_wallace._1958_ ;
 wire \u_cpu.ALU.u_wallace._1959_ ;
 wire \u_cpu.ALU.u_wallace._1960_ ;
 wire \u_cpu.ALU.u_wallace._1961_ ;
 wire \u_cpu.ALU.u_wallace._1962_ ;
 wire \u_cpu.ALU.u_wallace._1963_ ;
 wire \u_cpu.ALU.u_wallace._1964_ ;
 wire \u_cpu.ALU.u_wallace._1965_ ;
 wire \u_cpu.ALU.u_wallace._1966_ ;
 wire \u_cpu.ALU.u_wallace._1967_ ;
 wire \u_cpu.ALU.u_wallace._1968_ ;
 wire \u_cpu.ALU.u_wallace._1969_ ;
 wire \u_cpu.ALU.u_wallace._1970_ ;
 wire \u_cpu.ALU.u_wallace._1971_ ;
 wire \u_cpu.ALU.u_wallace._1972_ ;
 wire \u_cpu.ALU.u_wallace._1973_ ;
 wire \u_cpu.ALU.u_wallace._1974_ ;
 wire \u_cpu.ALU.u_wallace._1975_ ;
 wire \u_cpu.ALU.u_wallace._1976_ ;
 wire \u_cpu.ALU.u_wallace._1977_ ;
 wire \u_cpu.ALU.u_wallace._1978_ ;
 wire \u_cpu.ALU.u_wallace._1979_ ;
 wire \u_cpu.ALU.u_wallace._1980_ ;
 wire \u_cpu.ALU.u_wallace._1981_ ;
 wire \u_cpu.ALU.u_wallace._1982_ ;
 wire \u_cpu.ALU.u_wallace._1983_ ;
 wire \u_cpu.ALU.u_wallace._1984_ ;
 wire \u_cpu.ALU.u_wallace._1985_ ;
 wire \u_cpu.ALU.u_wallace._1986_ ;
 wire \u_cpu.ALU.u_wallace._1987_ ;
 wire \u_cpu.ALU.u_wallace._1988_ ;
 wire \u_cpu.ALU.u_wallace._1989_ ;
 wire \u_cpu.ALU.u_wallace._1990_ ;
 wire \u_cpu.ALU.u_wallace._1991_ ;
 wire \u_cpu.ALU.u_wallace._1992_ ;
 wire \u_cpu.ALU.u_wallace._1993_ ;
 wire \u_cpu.ALU.u_wallace._1994_ ;
 wire \u_cpu.ALU.u_wallace._1995_ ;
 wire \u_cpu.ALU.u_wallace._1996_ ;
 wire \u_cpu.ALU.u_wallace._1997_ ;
 wire \u_cpu.ALU.u_wallace._1998_ ;
 wire \u_cpu.ALU.u_wallace._1999_ ;
 wire \u_cpu.ALU.u_wallace._2000_ ;
 wire \u_cpu.ALU.u_wallace._2001_ ;
 wire \u_cpu.ALU.u_wallace._2002_ ;
 wire \u_cpu.ALU.u_wallace._2003_ ;
 wire \u_cpu.ALU.u_wallace._2004_ ;
 wire \u_cpu.ALU.u_wallace._2005_ ;
 wire \u_cpu.ALU.u_wallace._2006_ ;
 wire \u_cpu.ALU.u_wallace._2007_ ;
 wire \u_cpu.ALU.u_wallace._2008_ ;
 wire \u_cpu.ALU.u_wallace._2009_ ;
 wire \u_cpu.ALU.u_wallace._2010_ ;
 wire \u_cpu.ALU.u_wallace._2011_ ;
 wire \u_cpu.ALU.u_wallace._2012_ ;
 wire \u_cpu.ALU.u_wallace._2013_ ;
 wire \u_cpu.ALU.u_wallace._2014_ ;
 wire \u_cpu.ALU.u_wallace._2015_ ;
 wire \u_cpu.ALU.u_wallace._2016_ ;
 wire \u_cpu.ALU.u_wallace._2017_ ;
 wire \u_cpu.ALU.u_wallace._2018_ ;
 wire \u_cpu.ALU.u_wallace._2019_ ;
 wire \u_cpu.ALU.u_wallace._2020_ ;
 wire \u_cpu.ALU.u_wallace._2021_ ;
 wire \u_cpu.ALU.u_wallace._2022_ ;
 wire \u_cpu.ALU.u_wallace._2023_ ;
 wire \u_cpu.ALU.u_wallace._2024_ ;
 wire \u_cpu.ALU.u_wallace._2025_ ;
 wire \u_cpu.ALU.u_wallace._2026_ ;
 wire \u_cpu.ALU.u_wallace._2027_ ;
 wire \u_cpu.ALU.u_wallace._2028_ ;
 wire \u_cpu.ALU.u_wallace._2029_ ;
 wire \u_cpu.ALU.u_wallace._2030_ ;
 wire \u_cpu.ALU.u_wallace._2031_ ;
 wire \u_cpu.ALU.u_wallace._2032_ ;
 wire \u_cpu.ALU.u_wallace._2033_ ;
 wire \u_cpu.ALU.u_wallace._2034_ ;
 wire \u_cpu.ALU.u_wallace._2035_ ;
 wire \u_cpu.ALU.u_wallace._2036_ ;
 wire \u_cpu.ALU.u_wallace._2037_ ;
 wire \u_cpu.ALU.u_wallace._2038_ ;
 wire \u_cpu.ALU.u_wallace._2039_ ;
 wire \u_cpu.ALU.u_wallace._2040_ ;
 wire \u_cpu.ALU.u_wallace._2041_ ;
 wire \u_cpu.ALU.u_wallace._2042_ ;
 wire \u_cpu.ALU.u_wallace._2043_ ;
 wire \u_cpu.ALU.u_wallace._2044_ ;
 wire \u_cpu.ALU.u_wallace._2045_ ;
 wire \u_cpu.ALU.u_wallace._2046_ ;
 wire \u_cpu.ALU.u_wallace._2047_ ;
 wire \u_cpu.ALU.u_wallace._2048_ ;
 wire \u_cpu.ALU.u_wallace._2049_ ;
 wire \u_cpu.ALU.u_wallace._2050_ ;
 wire \u_cpu.ALU.u_wallace._2051_ ;
 wire \u_cpu.ALU.u_wallace._2052_ ;
 wire \u_cpu.ALU.u_wallace._2053_ ;
 wire \u_cpu.ALU.u_wallace._2054_ ;
 wire \u_cpu.ALU.u_wallace._2055_ ;
 wire \u_cpu.ALU.u_wallace._2056_ ;
 wire \u_cpu.ALU.u_wallace._2057_ ;
 wire \u_cpu.ALU.u_wallace._2058_ ;
 wire \u_cpu.ALU.u_wallace._2059_ ;
 wire \u_cpu.ALU.u_wallace._2060_ ;
 wire \u_cpu.ALU.u_wallace._2061_ ;
 wire \u_cpu.ALU.u_wallace._2062_ ;
 wire \u_cpu.ALU.u_wallace._2063_ ;
 wire \u_cpu.ALU.u_wallace._2064_ ;
 wire \u_cpu.ALU.u_wallace._2065_ ;
 wire \u_cpu.ALU.u_wallace._2066_ ;
 wire \u_cpu.ALU.u_wallace._2067_ ;
 wire \u_cpu.ALU.u_wallace._2068_ ;
 wire \u_cpu.ALU.u_wallace._2069_ ;
 wire \u_cpu.ALU.u_wallace._2070_ ;
 wire \u_cpu.ALU.u_wallace._2071_ ;
 wire \u_cpu.ALU.u_wallace._2072_ ;
 wire \u_cpu.ALU.u_wallace._2073_ ;
 wire \u_cpu.ALU.u_wallace._2074_ ;
 wire \u_cpu.ALU.u_wallace._2075_ ;
 wire \u_cpu.ALU.u_wallace._2076_ ;
 wire \u_cpu.ALU.u_wallace._2077_ ;
 wire \u_cpu.ALU.u_wallace._2078_ ;
 wire \u_cpu.ALU.u_wallace._2079_ ;
 wire \u_cpu.ALU.u_wallace._2080_ ;
 wire \u_cpu.ALU.u_wallace._2081_ ;
 wire \u_cpu.ALU.u_wallace._2082_ ;
 wire \u_cpu.ALU.u_wallace._2083_ ;
 wire \u_cpu.ALU.u_wallace._2084_ ;
 wire \u_cpu.ALU.u_wallace._2085_ ;
 wire \u_cpu.ALU.u_wallace._2086_ ;
 wire \u_cpu.ALU.u_wallace._2087_ ;
 wire \u_cpu.ALU.u_wallace._2088_ ;
 wire \u_cpu.ALU.u_wallace._2089_ ;
 wire \u_cpu.ALU.u_wallace._2090_ ;
 wire \u_cpu.ALU.u_wallace._2091_ ;
 wire \u_cpu.ALU.u_wallace._2092_ ;
 wire \u_cpu.ALU.u_wallace._2093_ ;
 wire \u_cpu.ALU.u_wallace._2094_ ;
 wire \u_cpu.ALU.u_wallace._2095_ ;
 wire \u_cpu.ALU.u_wallace._2096_ ;
 wire \u_cpu.ALU.u_wallace._2097_ ;
 wire \u_cpu.ALU.u_wallace._2098_ ;
 wire \u_cpu.ALU.u_wallace._2099_ ;
 wire \u_cpu.ALU.u_wallace._2100_ ;
 wire \u_cpu.ALU.u_wallace._2101_ ;
 wire \u_cpu.ALU.u_wallace._2102_ ;
 wire \u_cpu.ALU.u_wallace._2103_ ;
 wire \u_cpu.ALU.u_wallace._2104_ ;
 wire \u_cpu.ALU.u_wallace._2105_ ;
 wire \u_cpu.ALU.u_wallace._2106_ ;
 wire \u_cpu.ALU.u_wallace._2107_ ;
 wire \u_cpu.ALU.u_wallace._2108_ ;
 wire \u_cpu.ALU.u_wallace._2109_ ;
 wire \u_cpu.ALU.u_wallace._2110_ ;
 wire \u_cpu.ALU.u_wallace._2111_ ;
 wire \u_cpu.ALU.u_wallace._2112_ ;
 wire \u_cpu.ALU.u_wallace._2113_ ;
 wire \u_cpu.ALU.u_wallace._2114_ ;
 wire \u_cpu.ALU.u_wallace._2115_ ;
 wire \u_cpu.ALU.u_wallace._2116_ ;
 wire \u_cpu.ALU.u_wallace._2117_ ;
 wire \u_cpu.ALU.u_wallace._2118_ ;
 wire \u_cpu.ALU.u_wallace._2119_ ;
 wire \u_cpu.ALU.u_wallace._2120_ ;
 wire \u_cpu.ALU.u_wallace._2121_ ;
 wire \u_cpu.ALU.u_wallace._2122_ ;
 wire \u_cpu.ALU.u_wallace._2123_ ;
 wire \u_cpu.ALU.u_wallace._2124_ ;
 wire \u_cpu.ALU.u_wallace._2125_ ;
 wire \u_cpu.ALU.u_wallace._2126_ ;
 wire \u_cpu.ALU.u_wallace._2127_ ;
 wire \u_cpu.ALU.u_wallace._2128_ ;
 wire \u_cpu.ALU.u_wallace._2129_ ;
 wire \u_cpu.ALU.u_wallace._2130_ ;
 wire \u_cpu.ALU.u_wallace._2131_ ;
 wire \u_cpu.ALU.u_wallace._2132_ ;
 wire \u_cpu.ALU.u_wallace._2133_ ;
 wire \u_cpu.ALU.u_wallace._2134_ ;
 wire \u_cpu.ALU.u_wallace._2135_ ;
 wire \u_cpu.ALU.u_wallace._2136_ ;
 wire \u_cpu.ALU.u_wallace._2137_ ;
 wire \u_cpu.ALU.u_wallace._2138_ ;
 wire \u_cpu.ALU.u_wallace._2139_ ;
 wire \u_cpu.ALU.u_wallace._2140_ ;
 wire \u_cpu.ALU.u_wallace._2141_ ;
 wire \u_cpu.ALU.u_wallace._2142_ ;
 wire \u_cpu.ALU.u_wallace._2143_ ;
 wire \u_cpu.ALU.u_wallace._2144_ ;
 wire \u_cpu.ALU.u_wallace._2145_ ;
 wire \u_cpu.ALU.u_wallace._2146_ ;
 wire \u_cpu.ALU.u_wallace._2147_ ;
 wire \u_cpu.ALU.u_wallace._2148_ ;
 wire \u_cpu.ALU.u_wallace._2149_ ;
 wire \u_cpu.ALU.u_wallace._2150_ ;
 wire \u_cpu.ALU.u_wallace._2151_ ;
 wire \u_cpu.ALU.u_wallace._2152_ ;
 wire \u_cpu.ALU.u_wallace._2153_ ;
 wire \u_cpu.ALU.u_wallace._2154_ ;
 wire \u_cpu.ALU.u_wallace._2155_ ;
 wire \u_cpu.ALU.u_wallace._2156_ ;
 wire \u_cpu.ALU.u_wallace._2157_ ;
 wire \u_cpu.ALU.u_wallace._2158_ ;
 wire \u_cpu.ALU.u_wallace._2159_ ;
 wire \u_cpu.ALU.u_wallace._2160_ ;
 wire \u_cpu.ALU.u_wallace._2161_ ;
 wire \u_cpu.ALU.u_wallace._2162_ ;
 wire \u_cpu.ALU.u_wallace._2163_ ;
 wire \u_cpu.ALU.u_wallace._2164_ ;
 wire \u_cpu.ALU.u_wallace._2165_ ;
 wire \u_cpu.ALU.u_wallace._2166_ ;
 wire \u_cpu.ALU.u_wallace._2167_ ;
 wire \u_cpu.ALU.u_wallace._2168_ ;
 wire \u_cpu.ALU.u_wallace._2169_ ;
 wire \u_cpu.ALU.u_wallace._2170_ ;
 wire \u_cpu.ALU.u_wallace._2171_ ;
 wire \u_cpu.ALU.u_wallace._2172_ ;
 wire \u_cpu.ALU.u_wallace._2173_ ;
 wire \u_cpu.ALU.u_wallace._2174_ ;
 wire \u_cpu.ALU.u_wallace._2175_ ;
 wire \u_cpu.ALU.u_wallace._2176_ ;
 wire \u_cpu.ALU.u_wallace._2177_ ;
 wire \u_cpu.ALU.u_wallace._2178_ ;
 wire \u_cpu.ALU.u_wallace._2179_ ;
 wire \u_cpu.ALU.u_wallace._2180_ ;
 wire \u_cpu.ALU.u_wallace._2181_ ;
 wire \u_cpu.ALU.u_wallace._2182_ ;
 wire \u_cpu.ALU.u_wallace._2183_ ;
 wire \u_cpu.ALU.u_wallace._2184_ ;
 wire \u_cpu.ALU.u_wallace._2185_ ;
 wire \u_cpu.ALU.u_wallace._2186_ ;
 wire \u_cpu.ALU.u_wallace._2187_ ;
 wire \u_cpu.ALU.u_wallace._2188_ ;
 wire \u_cpu.ALU.u_wallace._2189_ ;
 wire \u_cpu.ALU.u_wallace._2190_ ;
 wire \u_cpu.ALU.u_wallace._2191_ ;
 wire \u_cpu.ALU.u_wallace._2192_ ;
 wire \u_cpu.ALU.u_wallace._2193_ ;
 wire \u_cpu.ALU.u_wallace._2194_ ;
 wire \u_cpu.ALU.u_wallace._2195_ ;
 wire \u_cpu.ALU.u_wallace._2196_ ;
 wire \u_cpu.ALU.u_wallace._2197_ ;
 wire \u_cpu.ALU.u_wallace._2198_ ;
 wire \u_cpu.ALU.u_wallace._2199_ ;
 wire \u_cpu.ALU.u_wallace._2200_ ;
 wire \u_cpu.ALU.u_wallace._2201_ ;
 wire \u_cpu.ALU.u_wallace._2202_ ;
 wire \u_cpu.ALU.u_wallace._2203_ ;
 wire \u_cpu.ALU.u_wallace._2204_ ;
 wire \u_cpu.ALU.u_wallace._2205_ ;
 wire \u_cpu.ALU.u_wallace._2206_ ;
 wire \u_cpu.ALU.u_wallace._2207_ ;
 wire \u_cpu.ALU.u_wallace._2208_ ;
 wire \u_cpu.ALU.u_wallace._2209_ ;
 wire \u_cpu.ALU.u_wallace._2210_ ;
 wire \u_cpu.ALU.u_wallace._2211_ ;
 wire \u_cpu.ALU.u_wallace._2212_ ;
 wire \u_cpu.ALU.u_wallace._2213_ ;
 wire \u_cpu.ALU.u_wallace._2214_ ;
 wire \u_cpu.ALU.u_wallace._2215_ ;
 wire \u_cpu.ALU.u_wallace._2216_ ;
 wire \u_cpu.ALU.u_wallace._2217_ ;
 wire \u_cpu.ALU.u_wallace._2218_ ;
 wire \u_cpu.ALU.u_wallace._2219_ ;
 wire \u_cpu.ALU.u_wallace._2220_ ;
 wire \u_cpu.ALU.u_wallace._2221_ ;
 wire \u_cpu.ALU.u_wallace._2222_ ;
 wire \u_cpu.ALU.u_wallace._2223_ ;
 wire \u_cpu.ALU.u_wallace._2224_ ;
 wire \u_cpu.ALU.u_wallace._2225_ ;
 wire \u_cpu.ALU.u_wallace._2226_ ;
 wire \u_cpu.ALU.u_wallace._2227_ ;
 wire \u_cpu.ALU.u_wallace._2228_ ;
 wire \u_cpu.ALU.u_wallace._2229_ ;
 wire \u_cpu.ALU.u_wallace._2230_ ;
 wire \u_cpu.ALU.u_wallace._2231_ ;
 wire \u_cpu.ALU.u_wallace._2232_ ;
 wire \u_cpu.ALU.u_wallace._2233_ ;
 wire \u_cpu.ALU.u_wallace._2234_ ;
 wire \u_cpu.ALU.u_wallace._2235_ ;
 wire \u_cpu.ALU.u_wallace._2236_ ;
 wire \u_cpu.ALU.u_wallace._2237_ ;
 wire \u_cpu.ALU.u_wallace._2238_ ;
 wire \u_cpu.ALU.u_wallace._2239_ ;
 wire \u_cpu.ALU.u_wallace._2240_ ;
 wire \u_cpu.ALU.u_wallace._2241_ ;
 wire \u_cpu.ALU.u_wallace._2242_ ;
 wire \u_cpu.ALU.u_wallace._2243_ ;
 wire \u_cpu.ALU.u_wallace._2244_ ;
 wire \u_cpu.ALU.u_wallace._2245_ ;
 wire \u_cpu.ALU.u_wallace._2246_ ;
 wire \u_cpu.ALU.u_wallace._2247_ ;
 wire \u_cpu.ALU.u_wallace._2248_ ;
 wire \u_cpu.ALU.u_wallace._2249_ ;
 wire \u_cpu.ALU.u_wallace._2250_ ;
 wire \u_cpu.ALU.u_wallace._2251_ ;
 wire \u_cpu.ALU.u_wallace._2252_ ;
 wire \u_cpu.ALU.u_wallace._2253_ ;
 wire \u_cpu.ALU.u_wallace._2254_ ;
 wire \u_cpu.ALU.u_wallace._2255_ ;
 wire \u_cpu.ALU.u_wallace._2256_ ;
 wire \u_cpu.ALU.u_wallace._2257_ ;
 wire \u_cpu.ALU.u_wallace._2258_ ;
 wire \u_cpu.ALU.u_wallace._2259_ ;
 wire \u_cpu.ALU.u_wallace._2260_ ;
 wire \u_cpu.ALU.u_wallace._2261_ ;
 wire \u_cpu.ALU.u_wallace._2262_ ;
 wire \u_cpu.ALU.u_wallace._2263_ ;
 wire \u_cpu.ALU.u_wallace._2264_ ;
 wire \u_cpu.ALU.u_wallace._2265_ ;
 wire \u_cpu.ALU.u_wallace._2266_ ;
 wire \u_cpu.ALU.u_wallace._2267_ ;
 wire \u_cpu.ALU.u_wallace._2268_ ;
 wire \u_cpu.ALU.u_wallace._2269_ ;
 wire \u_cpu.ALU.u_wallace._2270_ ;
 wire \u_cpu.ALU.u_wallace._2271_ ;
 wire \u_cpu.ALU.u_wallace._2272_ ;
 wire \u_cpu.ALU.u_wallace._2273_ ;
 wire \u_cpu.ALU.u_wallace._2274_ ;
 wire \u_cpu.ALU.u_wallace._2275_ ;
 wire \u_cpu.ALU.u_wallace._2276_ ;
 wire \u_cpu.ALU.u_wallace._2277_ ;
 wire \u_cpu.ALU.u_wallace._2278_ ;
 wire \u_cpu.ALU.u_wallace._2279_ ;
 wire \u_cpu.ALU.u_wallace._2280_ ;
 wire \u_cpu.ALU.u_wallace._2281_ ;
 wire \u_cpu.ALU.u_wallace._2282_ ;
 wire \u_cpu.ALU.u_wallace._2283_ ;
 wire \u_cpu.ALU.u_wallace._2284_ ;
 wire \u_cpu.ALU.u_wallace._2285_ ;
 wire \u_cpu.ALU.u_wallace._2286_ ;
 wire \u_cpu.ALU.u_wallace._2287_ ;
 wire \u_cpu.ALU.u_wallace._2288_ ;
 wire \u_cpu.ALU.u_wallace._2289_ ;
 wire \u_cpu.ALU.u_wallace._2290_ ;
 wire \u_cpu.ALU.u_wallace._2291_ ;
 wire \u_cpu.ALU.u_wallace._2292_ ;
 wire \u_cpu.ALU.u_wallace._2293_ ;
 wire \u_cpu.ALU.u_wallace._2294_ ;
 wire \u_cpu.ALU.u_wallace._2295_ ;
 wire \u_cpu.ALU.u_wallace._2296_ ;
 wire \u_cpu.ALU.u_wallace._2297_ ;
 wire \u_cpu.ALU.u_wallace._2298_ ;
 wire \u_cpu.ALU.u_wallace._2299_ ;
 wire \u_cpu.ALU.u_wallace._2300_ ;
 wire \u_cpu.ALU.u_wallace._2301_ ;
 wire \u_cpu.ALU.u_wallace._2302_ ;
 wire \u_cpu.ALU.u_wallace._2303_ ;
 wire \u_cpu.ALU.u_wallace._2304_ ;
 wire \u_cpu.ALU.u_wallace._2305_ ;
 wire \u_cpu.ALU.u_wallace._2306_ ;
 wire \u_cpu.ALU.u_wallace._2307_ ;
 wire \u_cpu.ALU.u_wallace._2308_ ;
 wire \u_cpu.ALU.u_wallace._2309_ ;
 wire \u_cpu.ALU.u_wallace._2310_ ;
 wire \u_cpu.ALU.u_wallace._2311_ ;
 wire \u_cpu.ALU.u_wallace._2312_ ;
 wire \u_cpu.ALU.u_wallace._2313_ ;
 wire \u_cpu.ALU.u_wallace._2314_ ;
 wire \u_cpu.ALU.u_wallace._2315_ ;
 wire \u_cpu.ALU.u_wallace._2316_ ;
 wire \u_cpu.ALU.u_wallace._2317_ ;
 wire \u_cpu.ALU.u_wallace._2318_ ;
 wire \u_cpu.ALU.u_wallace._2319_ ;
 wire \u_cpu.ALU.u_wallace._2320_ ;
 wire \u_cpu.ALU.u_wallace._2321_ ;
 wire \u_cpu.ALU.u_wallace._2322_ ;
 wire \u_cpu.ALU.u_wallace._2323_ ;
 wire \u_cpu.ALU.u_wallace._2324_ ;
 wire \u_cpu.ALU.u_wallace._2325_ ;
 wire \u_cpu.ALU.u_wallace._2326_ ;
 wire \u_cpu.ALU.u_wallace._2327_ ;
 wire \u_cpu.ALU.u_wallace._2328_ ;
 wire \u_cpu.ALU.u_wallace._2329_ ;
 wire \u_cpu.ALU.u_wallace._2330_ ;
 wire \u_cpu.ALU.u_wallace._2331_ ;
 wire \u_cpu.ALU.u_wallace._2332_ ;
 wire \u_cpu.ALU.u_wallace._2333_ ;
 wire \u_cpu.ALU.u_wallace._2334_ ;
 wire \u_cpu.ALU.u_wallace._2335_ ;
 wire \u_cpu.ALU.u_wallace._2336_ ;
 wire \u_cpu.ALU.u_wallace._2337_ ;
 wire \u_cpu.ALU.u_wallace._2338_ ;
 wire \u_cpu.ALU.u_wallace._2339_ ;
 wire \u_cpu.ALU.u_wallace._2340_ ;
 wire \u_cpu.ALU.u_wallace._2341_ ;
 wire \u_cpu.ALU.u_wallace._2342_ ;
 wire \u_cpu.ALU.u_wallace._2343_ ;
 wire \u_cpu.ALU.u_wallace._2344_ ;
 wire \u_cpu.ALU.u_wallace._2345_ ;
 wire \u_cpu.ALU.u_wallace._2346_ ;
 wire \u_cpu.ALU.u_wallace._2347_ ;
 wire \u_cpu.ALU.u_wallace._2348_ ;
 wire \u_cpu.ALU.u_wallace._2349_ ;
 wire \u_cpu.ALU.u_wallace._2350_ ;
 wire \u_cpu.ALU.u_wallace._2351_ ;
 wire \u_cpu.ALU.u_wallace._2352_ ;
 wire \u_cpu.ALU.u_wallace._2353_ ;
 wire \u_cpu.ALU.u_wallace._2354_ ;
 wire \u_cpu.ALU.u_wallace._2355_ ;
 wire \u_cpu.ALU.u_wallace._2356_ ;
 wire \u_cpu.ALU.u_wallace._2357_ ;
 wire \u_cpu.ALU.u_wallace._2358_ ;
 wire \u_cpu.ALU.u_wallace._2359_ ;
 wire \u_cpu.ALU.u_wallace._2360_ ;
 wire \u_cpu.ALU.u_wallace._2361_ ;
 wire \u_cpu.ALU.u_wallace._2362_ ;
 wire \u_cpu.ALU.u_wallace._2363_ ;
 wire \u_cpu.ALU.u_wallace._2364_ ;
 wire \u_cpu.ALU.u_wallace._2365_ ;
 wire \u_cpu.ALU.u_wallace._2366_ ;
 wire \u_cpu.ALU.u_wallace._2367_ ;
 wire \u_cpu.ALU.u_wallace._2368_ ;
 wire \u_cpu.ALU.u_wallace._2369_ ;
 wire \u_cpu.ALU.u_wallace._2370_ ;
 wire \u_cpu.ALU.u_wallace._2371_ ;
 wire \u_cpu.ALU.u_wallace._2372_ ;
 wire \u_cpu.ALU.u_wallace._2373_ ;
 wire \u_cpu.ALU.u_wallace._2374_ ;
 wire \u_cpu.ALU.u_wallace._2375_ ;
 wire \u_cpu.ALU.u_wallace._2376_ ;
 wire \u_cpu.ALU.u_wallace._2377_ ;
 wire \u_cpu.ALU.u_wallace._2378_ ;
 wire \u_cpu.ALU.u_wallace._2379_ ;
 wire \u_cpu.ALU.u_wallace._2380_ ;
 wire \u_cpu.ALU.u_wallace._2381_ ;
 wire \u_cpu.ALU.u_wallace._2382_ ;
 wire \u_cpu.ALU.u_wallace._2383_ ;
 wire \u_cpu.ALU.u_wallace._2384_ ;
 wire \u_cpu.ALU.u_wallace._2385_ ;
 wire \u_cpu.ALU.u_wallace._2386_ ;
 wire \u_cpu.ALU.u_wallace._2387_ ;
 wire \u_cpu.ALU.u_wallace._2388_ ;
 wire \u_cpu.ALU.u_wallace._2389_ ;
 wire \u_cpu.ALU.u_wallace._2390_ ;
 wire \u_cpu.ALU.u_wallace._2391_ ;
 wire \u_cpu.ALU.u_wallace._2392_ ;
 wire \u_cpu.ALU.u_wallace._2393_ ;
 wire \u_cpu.ALU.u_wallace._2394_ ;
 wire \u_cpu.ALU.u_wallace._2395_ ;
 wire \u_cpu.ALU.u_wallace._2396_ ;
 wire \u_cpu.ALU.u_wallace._2397_ ;
 wire \u_cpu.ALU.u_wallace._2398_ ;
 wire \u_cpu.ALU.u_wallace._2399_ ;
 wire \u_cpu.ALU.u_wallace._2400_ ;
 wire \u_cpu.ALU.u_wallace._2401_ ;
 wire \u_cpu.ALU.u_wallace._2402_ ;
 wire \u_cpu.ALU.u_wallace._2403_ ;
 wire \u_cpu.ALU.u_wallace._2404_ ;
 wire \u_cpu.ALU.u_wallace._2405_ ;
 wire \u_cpu.ALU.u_wallace._2406_ ;
 wire \u_cpu.ALU.u_wallace._2407_ ;
 wire \u_cpu.ALU.u_wallace._2408_ ;
 wire \u_cpu.ALU.u_wallace._2409_ ;
 wire \u_cpu.ALU.u_wallace._2410_ ;
 wire \u_cpu.ALU.u_wallace._2411_ ;
 wire \u_cpu.ALU.u_wallace._2412_ ;
 wire \u_cpu.ALU.u_wallace._2413_ ;
 wire \u_cpu.ALU.u_wallace._2414_ ;
 wire \u_cpu.ALU.u_wallace._2415_ ;
 wire \u_cpu.ALU.u_wallace._2416_ ;
 wire \u_cpu.ALU.u_wallace._2417_ ;
 wire \u_cpu.ALU.u_wallace._2418_ ;
 wire \u_cpu.ALU.u_wallace._2419_ ;
 wire \u_cpu.ALU.u_wallace._2420_ ;
 wire \u_cpu.ALU.u_wallace._2421_ ;
 wire \u_cpu.ALU.u_wallace._2422_ ;
 wire \u_cpu.ALU.u_wallace._2423_ ;
 wire \u_cpu.ALU.u_wallace._2424_ ;
 wire \u_cpu.ALU.u_wallace._2425_ ;
 wire \u_cpu.ALU.u_wallace._2426_ ;
 wire \u_cpu.ALU.u_wallace._2427_ ;
 wire \u_cpu.ALU.u_wallace._2428_ ;
 wire \u_cpu.ALU.u_wallace._2429_ ;
 wire \u_cpu.ALU.u_wallace._2430_ ;
 wire \u_cpu.ALU.u_wallace._2431_ ;
 wire \u_cpu.ALU.u_wallace._2432_ ;
 wire \u_cpu.ALU.u_wallace._2433_ ;
 wire \u_cpu.ALU.u_wallace._2434_ ;
 wire \u_cpu.ALU.u_wallace._2435_ ;
 wire \u_cpu.ALU.u_wallace._2436_ ;
 wire \u_cpu.ALU.u_wallace._2437_ ;
 wire \u_cpu.ALU.u_wallace._2438_ ;
 wire \u_cpu.ALU.u_wallace._2439_ ;
 wire \u_cpu.ALU.u_wallace._2440_ ;
 wire \u_cpu.ALU.u_wallace._2441_ ;
 wire \u_cpu.ALU.u_wallace._2442_ ;
 wire \u_cpu.ALU.u_wallace._2443_ ;
 wire \u_cpu.ALU.u_wallace._2444_ ;
 wire \u_cpu.ALU.u_wallace._2445_ ;
 wire \u_cpu.ALU.u_wallace._2446_ ;
 wire \u_cpu.ALU.u_wallace._2447_ ;
 wire \u_cpu.ALU.u_wallace._2448_ ;
 wire \u_cpu.ALU.u_wallace._2449_ ;
 wire \u_cpu.ALU.u_wallace._2450_ ;
 wire \u_cpu.ALU.u_wallace._2451_ ;
 wire \u_cpu.ALU.u_wallace._2452_ ;
 wire \u_cpu.ALU.u_wallace._2453_ ;
 wire \u_cpu.ALU.u_wallace._2454_ ;
 wire \u_cpu.ALU.u_wallace._2455_ ;
 wire \u_cpu.ALU.u_wallace._2456_ ;
 wire \u_cpu.ALU.u_wallace._2457_ ;
 wire \u_cpu.ALU.u_wallace._2458_ ;
 wire \u_cpu.ALU.u_wallace._2459_ ;
 wire \u_cpu.ALU.u_wallace._2460_ ;
 wire \u_cpu.ALU.u_wallace._2461_ ;
 wire \u_cpu.ALU.u_wallace._2462_ ;
 wire \u_cpu.ALU.u_wallace._2463_ ;
 wire \u_cpu.ALU.u_wallace._2464_ ;
 wire \u_cpu.ALU.u_wallace._2465_ ;
 wire \u_cpu.ALU.u_wallace._2466_ ;
 wire \u_cpu.ALU.u_wallace._2467_ ;
 wire \u_cpu.ALU.u_wallace._2468_ ;
 wire \u_cpu.ALU.u_wallace._2469_ ;
 wire \u_cpu.ALU.u_wallace._2470_ ;
 wire \u_cpu.ALU.u_wallace._2471_ ;
 wire \u_cpu.ALU.u_wallace._2472_ ;
 wire \u_cpu.ALU.u_wallace._2473_ ;
 wire \u_cpu.ALU.u_wallace._2474_ ;
 wire \u_cpu.ALU.u_wallace._2475_ ;
 wire \u_cpu.ALU.u_wallace._2476_ ;
 wire \u_cpu.ALU.u_wallace._2477_ ;
 wire \u_cpu.ALU.u_wallace._2478_ ;
 wire \u_cpu.ALU.u_wallace._2479_ ;
 wire \u_cpu.ALU.u_wallace._2480_ ;
 wire \u_cpu.ALU.u_wallace._2481_ ;
 wire \u_cpu.ALU.u_wallace._2482_ ;
 wire \u_cpu.ALU.u_wallace._2483_ ;
 wire \u_cpu.ALU.u_wallace._2484_ ;
 wire \u_cpu.ALU.u_wallace._2485_ ;
 wire \u_cpu.ALU.u_wallace._2486_ ;
 wire \u_cpu.ALU.u_wallace._2487_ ;
 wire \u_cpu.ALU.u_wallace._2488_ ;
 wire \u_cpu.ALU.u_wallace._2489_ ;
 wire \u_cpu.ALU.u_wallace._2490_ ;
 wire \u_cpu.ALU.u_wallace._2491_ ;
 wire \u_cpu.ALU.u_wallace._2492_ ;
 wire \u_cpu.ALU.u_wallace._2493_ ;
 wire \u_cpu.ALU.u_wallace._2494_ ;
 wire \u_cpu.ALU.u_wallace._2495_ ;
 wire \u_cpu.ALU.u_wallace._2496_ ;
 wire \u_cpu.ALU.u_wallace._2497_ ;
 wire \u_cpu.ALU.u_wallace._2498_ ;
 wire \u_cpu.ALU.u_wallace._2499_ ;
 wire \u_cpu.ALU.u_wallace._2500_ ;
 wire \u_cpu.ALU.u_wallace._2501_ ;
 wire \u_cpu.ALU.u_wallace._2502_ ;
 wire \u_cpu.ALU.u_wallace._2503_ ;
 wire \u_cpu.ALU.u_wallace._2504_ ;
 wire \u_cpu.ALU.u_wallace._2505_ ;
 wire \u_cpu.ALU.u_wallace._2506_ ;
 wire \u_cpu.ALU.u_wallace._2507_ ;
 wire \u_cpu.ALU.u_wallace._2508_ ;
 wire \u_cpu.ALU.u_wallace._2509_ ;
 wire \u_cpu.ALU.u_wallace._2510_ ;
 wire \u_cpu.ALU.u_wallace._2511_ ;
 wire \u_cpu.ALU.u_wallace._2512_ ;
 wire \u_cpu.ALU.u_wallace._2513_ ;
 wire \u_cpu.ALU.u_wallace._2514_ ;
 wire \u_cpu.ALU.u_wallace._2515_ ;
 wire \u_cpu.ALU.u_wallace._2516_ ;
 wire \u_cpu.ALU.u_wallace._2517_ ;
 wire \u_cpu.ALU.u_wallace._2518_ ;
 wire \u_cpu.ALU.u_wallace._2519_ ;
 wire \u_cpu.ALU.u_wallace._2520_ ;
 wire \u_cpu.ALU.u_wallace._2521_ ;
 wire \u_cpu.ALU.u_wallace._2522_ ;
 wire \u_cpu.ALU.u_wallace._2523_ ;
 wire \u_cpu.ALU.u_wallace._2524_ ;
 wire \u_cpu.ALU.u_wallace._2525_ ;
 wire \u_cpu.ALU.u_wallace._2526_ ;
 wire \u_cpu.ALU.u_wallace._2527_ ;
 wire \u_cpu.ALU.u_wallace._2528_ ;
 wire \u_cpu.ALU.u_wallace._2529_ ;
 wire \u_cpu.ALU.u_wallace._2530_ ;
 wire \u_cpu.ALU.u_wallace._2531_ ;
 wire \u_cpu.ALU.u_wallace._2532_ ;
 wire \u_cpu.ALU.u_wallace._2533_ ;
 wire \u_cpu.ALU.u_wallace._2534_ ;
 wire \u_cpu.ALU.u_wallace._2535_ ;
 wire \u_cpu.ALU.u_wallace._2536_ ;
 wire \u_cpu.ALU.u_wallace._2537_ ;
 wire \u_cpu.ALU.u_wallace._2538_ ;
 wire \u_cpu.ALU.u_wallace._2539_ ;
 wire \u_cpu.ALU.u_wallace._2540_ ;
 wire \u_cpu.ALU.u_wallace._2541_ ;
 wire \u_cpu.ALU.u_wallace._2542_ ;
 wire \u_cpu.ALU.u_wallace._2543_ ;
 wire \u_cpu.ALU.u_wallace._2544_ ;
 wire \u_cpu.ALU.u_wallace._2545_ ;
 wire \u_cpu.ALU.u_wallace._2546_ ;
 wire \u_cpu.ALU.u_wallace._2547_ ;
 wire \u_cpu.ALU.u_wallace._2548_ ;
 wire \u_cpu.ALU.u_wallace._2549_ ;
 wire \u_cpu.ALU.u_wallace._2550_ ;
 wire \u_cpu.ALU.u_wallace._2551_ ;
 wire \u_cpu.ALU.u_wallace._2552_ ;
 wire \u_cpu.ALU.u_wallace._2553_ ;
 wire \u_cpu.ALU.u_wallace._2554_ ;
 wire \u_cpu.ALU.u_wallace._2555_ ;
 wire \u_cpu.ALU.u_wallace._2556_ ;
 wire \u_cpu.ALU.u_wallace._2557_ ;
 wire \u_cpu.ALU.u_wallace._2558_ ;
 wire \u_cpu.ALU.u_wallace._2559_ ;
 wire \u_cpu.ALU.u_wallace._2560_ ;
 wire \u_cpu.ALU.u_wallace._2561_ ;
 wire \u_cpu.ALU.u_wallace._2562_ ;
 wire \u_cpu.ALU.u_wallace._2563_ ;
 wire \u_cpu.ALU.u_wallace._2564_ ;
 wire \u_cpu.ALU.u_wallace._2565_ ;
 wire \u_cpu.ALU.u_wallace._2566_ ;
 wire \u_cpu.ALU.u_wallace._2567_ ;
 wire \u_cpu.ALU.u_wallace._2568_ ;
 wire \u_cpu.ALU.u_wallace._2569_ ;
 wire \u_cpu.ALU.u_wallace._2570_ ;
 wire \u_cpu.ALU.u_wallace._2571_ ;
 wire \u_cpu.ALU.u_wallace._2572_ ;
 wire \u_cpu.ALU.u_wallace._2573_ ;
 wire \u_cpu.ALU.u_wallace._2574_ ;
 wire \u_cpu.ALU.u_wallace._2575_ ;
 wire \u_cpu.ALU.u_wallace._2576_ ;
 wire \u_cpu.ALU.u_wallace._2577_ ;
 wire \u_cpu.ALU.u_wallace._2578_ ;
 wire \u_cpu.ALU.u_wallace._2579_ ;
 wire \u_cpu.ALU.u_wallace._2580_ ;
 wire \u_cpu.ALU.u_wallace._2581_ ;
 wire \u_cpu.ALU.u_wallace._2582_ ;
 wire \u_cpu.ALU.u_wallace._2583_ ;
 wire \u_cpu.ALU.u_wallace._2584_ ;
 wire \u_cpu.ALU.u_wallace._2585_ ;
 wire \u_cpu.ALU.u_wallace._2586_ ;
 wire \u_cpu.ALU.u_wallace._2587_ ;
 wire \u_cpu.ALU.u_wallace._2588_ ;
 wire \u_cpu.ALU.u_wallace._2589_ ;
 wire \u_cpu.ALU.u_wallace._2590_ ;
 wire \u_cpu.ALU.u_wallace._2591_ ;
 wire \u_cpu.ALU.u_wallace._2592_ ;
 wire \u_cpu.ALU.u_wallace._2593_ ;
 wire \u_cpu.ALU.u_wallace._2594_ ;
 wire \u_cpu.ALU.u_wallace._2595_ ;
 wire \u_cpu.ALU.u_wallace._2596_ ;
 wire \u_cpu.ALU.u_wallace._2597_ ;
 wire \u_cpu.ALU.u_wallace._2598_ ;
 wire \u_cpu.ALU.u_wallace._2599_ ;
 wire \u_cpu.ALU.u_wallace._2600_ ;
 wire \u_cpu.ALU.u_wallace._2601_ ;
 wire \u_cpu.ALU.u_wallace._2602_ ;
 wire \u_cpu.ALU.u_wallace._2603_ ;
 wire \u_cpu.ALU.u_wallace._2604_ ;
 wire \u_cpu.ALU.u_wallace._2605_ ;
 wire \u_cpu.ALU.u_wallace._2606_ ;
 wire \u_cpu.ALU.u_wallace._2607_ ;
 wire \u_cpu.ALU.u_wallace._2608_ ;
 wire \u_cpu.ALU.u_wallace._2609_ ;
 wire \u_cpu.ALU.u_wallace._2610_ ;
 wire \u_cpu.ALU.u_wallace._2611_ ;
 wire \u_cpu.ALU.u_wallace._2612_ ;
 wire \u_cpu.ALU.u_wallace._2613_ ;
 wire \u_cpu.ALU.u_wallace._2614_ ;
 wire \u_cpu.ALU.u_wallace._2615_ ;
 wire \u_cpu.ALU.u_wallace._2616_ ;
 wire \u_cpu.ALU.u_wallace._2617_ ;
 wire \u_cpu.ALU.u_wallace._2618_ ;
 wire \u_cpu.ALU.u_wallace._2619_ ;
 wire \u_cpu.ALU.u_wallace._2620_ ;
 wire \u_cpu.ALU.u_wallace._2621_ ;
 wire \u_cpu.ALU.u_wallace._2622_ ;
 wire \u_cpu.ALU.u_wallace._2623_ ;
 wire \u_cpu.ALU.u_wallace._2624_ ;
 wire \u_cpu.ALU.u_wallace._2625_ ;
 wire \u_cpu.ALU.u_wallace._2626_ ;
 wire \u_cpu.ALU.u_wallace._2627_ ;
 wire \u_cpu.ALU.u_wallace._2628_ ;
 wire \u_cpu.ALU.u_wallace._2629_ ;
 wire \u_cpu.ALU.u_wallace._2630_ ;
 wire \u_cpu.ALU.u_wallace._2631_ ;
 wire \u_cpu.ALU.u_wallace._2632_ ;
 wire \u_cpu.ALU.u_wallace._2633_ ;
 wire \u_cpu.ALU.u_wallace._2634_ ;
 wire \u_cpu.ALU.u_wallace._2635_ ;
 wire \u_cpu.ALU.u_wallace._2636_ ;
 wire \u_cpu.ALU.u_wallace._2637_ ;
 wire \u_cpu.ALU.u_wallace._2638_ ;
 wire \u_cpu.ALU.u_wallace._2639_ ;
 wire \u_cpu.ALU.u_wallace._2640_ ;
 wire \u_cpu.ALU.u_wallace._2641_ ;
 wire \u_cpu.ALU.u_wallace._2642_ ;
 wire \u_cpu.ALU.u_wallace._2643_ ;
 wire \u_cpu.ALU.u_wallace._2644_ ;
 wire \u_cpu.ALU.u_wallace._2645_ ;
 wire \u_cpu.ALU.u_wallace._2646_ ;
 wire \u_cpu.ALU.u_wallace._2647_ ;
 wire \u_cpu.ALU.u_wallace._2648_ ;
 wire \u_cpu.ALU.u_wallace._2649_ ;
 wire \u_cpu.ALU.u_wallace._2650_ ;
 wire \u_cpu.ALU.u_wallace._2651_ ;
 wire \u_cpu.ALU.u_wallace._2652_ ;
 wire \u_cpu.ALU.u_wallace._2653_ ;
 wire \u_cpu.ALU.u_wallace._2654_ ;
 wire \u_cpu.ALU.u_wallace._2655_ ;
 wire \u_cpu.ALU.u_wallace._2656_ ;
 wire \u_cpu.ALU.u_wallace._2657_ ;
 wire \u_cpu.ALU.u_wallace._2658_ ;
 wire \u_cpu.ALU.u_wallace._2659_ ;
 wire \u_cpu.ALU.u_wallace._2660_ ;
 wire \u_cpu.ALU.u_wallace._2661_ ;
 wire \u_cpu.ALU.u_wallace._2662_ ;
 wire \u_cpu.ALU.u_wallace._2663_ ;
 wire \u_cpu.ALU.u_wallace._2664_ ;
 wire \u_cpu.ALU.u_wallace._2665_ ;
 wire \u_cpu.ALU.u_wallace._2666_ ;
 wire \u_cpu.ALU.u_wallace._2667_ ;
 wire \u_cpu.ALU.u_wallace._2668_ ;
 wire \u_cpu.ALU.u_wallace._2669_ ;
 wire \u_cpu.ALU.u_wallace._2670_ ;
 wire \u_cpu.ALU.u_wallace._2671_ ;
 wire \u_cpu.ALU.u_wallace._2672_ ;
 wire \u_cpu.ALU.u_wallace._2673_ ;
 wire \u_cpu.ALU.u_wallace._2674_ ;
 wire \u_cpu.ALU.u_wallace._2675_ ;
 wire \u_cpu.ALU.u_wallace._2676_ ;
 wire \u_cpu.ALU.u_wallace._2677_ ;
 wire \u_cpu.ALU.u_wallace._2678_ ;
 wire \u_cpu.ALU.u_wallace._2679_ ;
 wire \u_cpu.ALU.u_wallace._2680_ ;
 wire \u_cpu.ALU.u_wallace._2681_ ;
 wire \u_cpu.ALU.u_wallace._2682_ ;
 wire \u_cpu.ALU.u_wallace._2683_ ;
 wire \u_cpu.ALU.u_wallace._2684_ ;
 wire \u_cpu.ALU.u_wallace._2685_ ;
 wire \u_cpu.ALU.u_wallace._2686_ ;
 wire \u_cpu.ALU.u_wallace._2687_ ;
 wire \u_cpu.ALU.u_wallace._2688_ ;
 wire \u_cpu.ALU.u_wallace._2689_ ;
 wire \u_cpu.ALU.u_wallace._2690_ ;
 wire \u_cpu.ALU.u_wallace._2691_ ;
 wire \u_cpu.ALU.u_wallace._2692_ ;
 wire \u_cpu.ALU.u_wallace._2693_ ;
 wire \u_cpu.ALU.u_wallace._2694_ ;
 wire \u_cpu.ALU.u_wallace._2695_ ;
 wire \u_cpu.ALU.u_wallace._2696_ ;
 wire \u_cpu.ALU.u_wallace._2697_ ;
 wire \u_cpu.ALU.u_wallace._2698_ ;
 wire \u_cpu.ALU.u_wallace._2699_ ;
 wire \u_cpu.ALU.u_wallace._2700_ ;
 wire \u_cpu.ALU.u_wallace._2701_ ;
 wire \u_cpu.ALU.u_wallace._2702_ ;
 wire \u_cpu.ALU.u_wallace._2703_ ;
 wire \u_cpu.ALU.u_wallace._2704_ ;
 wire \u_cpu.ALU.u_wallace._2705_ ;
 wire \u_cpu.ALU.u_wallace._2706_ ;
 wire \u_cpu.ALU.u_wallace._2707_ ;
 wire \u_cpu.ALU.u_wallace._2708_ ;
 wire \u_cpu.ALU.u_wallace._2709_ ;
 wire \u_cpu.ALU.u_wallace._2710_ ;
 wire \u_cpu.ALU.u_wallace._2711_ ;
 wire \u_cpu.ALU.u_wallace._2712_ ;
 wire \u_cpu.ALU.u_wallace._2713_ ;
 wire \u_cpu.ALU.u_wallace._2714_ ;
 wire \u_cpu.ALU.u_wallace._2715_ ;
 wire \u_cpu.ALU.u_wallace._2716_ ;
 wire \u_cpu.ALU.u_wallace._2717_ ;
 wire \u_cpu.ALU.u_wallace._2718_ ;
 wire \u_cpu.ALU.u_wallace._2719_ ;
 wire \u_cpu.ALU.u_wallace._2720_ ;
 wire \u_cpu.ALU.u_wallace._2721_ ;
 wire \u_cpu.ALU.u_wallace._2722_ ;
 wire \u_cpu.ALU.u_wallace._2723_ ;
 wire \u_cpu.ALU.u_wallace._2724_ ;
 wire \u_cpu.ALU.u_wallace._2725_ ;
 wire \u_cpu.ALU.u_wallace._2726_ ;
 wire \u_cpu.ALU.u_wallace._2727_ ;
 wire \u_cpu.ALU.u_wallace._2728_ ;
 wire \u_cpu.ALU.u_wallace._2729_ ;
 wire \u_cpu.ALU.u_wallace._2730_ ;
 wire \u_cpu.ALU.u_wallace._2731_ ;
 wire \u_cpu.ALU.u_wallace._2732_ ;
 wire \u_cpu.ALU.u_wallace._2733_ ;
 wire \u_cpu.ALU.u_wallace._2734_ ;
 wire \u_cpu.ALU.u_wallace._2735_ ;
 wire \u_cpu.ALU.u_wallace._2736_ ;
 wire \u_cpu.ALU.u_wallace._2737_ ;
 wire \u_cpu.ALU.u_wallace._2738_ ;
 wire \u_cpu.ALU.u_wallace._2739_ ;
 wire \u_cpu.ALU.u_wallace._2740_ ;
 wire \u_cpu.ALU.u_wallace._2741_ ;
 wire \u_cpu.ALU.u_wallace._2742_ ;
 wire \u_cpu.ALU.u_wallace._2743_ ;
 wire \u_cpu.ALU.u_wallace._2744_ ;
 wire \u_cpu.ALU.u_wallace._2745_ ;
 wire \u_cpu.ALU.u_wallace._2746_ ;
 wire \u_cpu.ALU.u_wallace._2747_ ;
 wire \u_cpu.ALU.u_wallace._2748_ ;
 wire \u_cpu.ALU.u_wallace._2749_ ;
 wire \u_cpu.ALU.u_wallace._2750_ ;
 wire \u_cpu.ALU.u_wallace._2751_ ;
 wire \u_cpu.ALU.u_wallace._2752_ ;
 wire \u_cpu.ALU.u_wallace._2753_ ;
 wire \u_cpu.ALU.u_wallace._2754_ ;
 wire \u_cpu.ALU.u_wallace._2755_ ;
 wire \u_cpu.ALU.u_wallace._2756_ ;
 wire \u_cpu.ALU.u_wallace._2757_ ;
 wire \u_cpu.ALU.u_wallace._2758_ ;
 wire \u_cpu.ALU.u_wallace._2759_ ;
 wire \u_cpu.ALU.u_wallace._2760_ ;
 wire \u_cpu.ALU.u_wallace._2761_ ;
 wire \u_cpu.ALU.u_wallace._2762_ ;
 wire \u_cpu.ALU.u_wallace._2763_ ;
 wire \u_cpu.ALU.u_wallace._2764_ ;
 wire \u_cpu.ALU.u_wallace._2765_ ;
 wire \u_cpu.ALU.u_wallace._2766_ ;
 wire \u_cpu.ALU.u_wallace._2767_ ;
 wire \u_cpu.ALU.u_wallace._2768_ ;
 wire \u_cpu.ALU.u_wallace._2769_ ;
 wire \u_cpu.ALU.u_wallace._2770_ ;
 wire \u_cpu.ALU.u_wallace._2771_ ;
 wire \u_cpu.ALU.u_wallace._2772_ ;
 wire \u_cpu.ALU.u_wallace._2773_ ;
 wire \u_cpu.ALU.u_wallace._2774_ ;
 wire \u_cpu.ALU.u_wallace._2775_ ;
 wire \u_cpu.ALU.u_wallace._2776_ ;
 wire \u_cpu.ALU.u_wallace._2777_ ;
 wire \u_cpu.ALU.u_wallace._2778_ ;
 wire \u_cpu.ALU.u_wallace._2779_ ;
 wire \u_cpu.ALU.u_wallace._2780_ ;
 wire \u_cpu.ALU.u_wallace._2781_ ;
 wire \u_cpu.ALU.u_wallace._2782_ ;
 wire \u_cpu.ALU.u_wallace._2783_ ;
 wire \u_cpu.ALU.u_wallace._2784_ ;
 wire \u_cpu.ALU.u_wallace._2785_ ;
 wire \u_cpu.ALU.u_wallace._2786_ ;
 wire \u_cpu.ALU.u_wallace._2787_ ;
 wire \u_cpu.ALU.u_wallace._2788_ ;
 wire \u_cpu.ALU.u_wallace._2789_ ;
 wire \u_cpu.ALU.u_wallace._2790_ ;
 wire \u_cpu.ALU.u_wallace._2791_ ;
 wire \u_cpu.ALU.u_wallace._2792_ ;
 wire \u_cpu.ALU.u_wallace._2793_ ;
 wire \u_cpu.ALU.u_wallace._2794_ ;
 wire \u_cpu.ALU.u_wallace._2795_ ;
 wire \u_cpu.ALU.u_wallace._2796_ ;
 wire \u_cpu.ALU.u_wallace._2797_ ;
 wire \u_cpu.ALU.u_wallace._2798_ ;
 wire \u_cpu.ALU.u_wallace._2799_ ;
 wire \u_cpu.ALU.u_wallace._2800_ ;
 wire \u_cpu.ALU.u_wallace._2801_ ;
 wire \u_cpu.ALU.u_wallace._2802_ ;
 wire \u_cpu.ALU.u_wallace._2803_ ;
 wire \u_cpu.ALU.u_wallace._2804_ ;
 wire \u_cpu.ALU.u_wallace._2805_ ;
 wire \u_cpu.ALU.u_wallace._2806_ ;
 wire \u_cpu.ALU.u_wallace._2807_ ;
 wire \u_cpu.ALU.u_wallace._2808_ ;
 wire \u_cpu.ALU.u_wallace._2809_ ;
 wire \u_cpu.ALU.u_wallace._2810_ ;
 wire \u_cpu.ALU.u_wallace._2811_ ;
 wire \u_cpu.ALU.u_wallace._2812_ ;
 wire \u_cpu.ALU.u_wallace._2813_ ;
 wire \u_cpu.ALU.u_wallace._2814_ ;
 wire \u_cpu.ALU.u_wallace._2815_ ;
 wire \u_cpu.ALU.u_wallace._2816_ ;
 wire \u_cpu.ALU.u_wallace._2817_ ;
 wire \u_cpu.ALU.u_wallace._2818_ ;
 wire \u_cpu.ALU.u_wallace._2819_ ;
 wire \u_cpu.ALU.u_wallace._2820_ ;
 wire \u_cpu.ALU.u_wallace._2821_ ;
 wire \u_cpu.ALU.u_wallace._2822_ ;
 wire \u_cpu.ALU.u_wallace._2823_ ;
 wire \u_cpu.ALU.u_wallace._2824_ ;
 wire \u_cpu.ALU.u_wallace._2825_ ;
 wire \u_cpu.ALU.u_wallace._2826_ ;
 wire \u_cpu.ALU.u_wallace._2827_ ;
 wire \u_cpu.ALU.u_wallace._2828_ ;
 wire \u_cpu.ALU.u_wallace._2829_ ;
 wire \u_cpu.ALU.u_wallace._2830_ ;
 wire \u_cpu.ALU.u_wallace._2831_ ;
 wire \u_cpu.ALU.u_wallace._2832_ ;
 wire \u_cpu.ALU.u_wallace._2833_ ;
 wire \u_cpu.ALU.u_wallace._2834_ ;
 wire \u_cpu.ALU.u_wallace._2835_ ;
 wire \u_cpu.ALU.u_wallace._2836_ ;
 wire \u_cpu.ALU.u_wallace._2837_ ;
 wire \u_cpu.ALU.u_wallace._2838_ ;
 wire \u_cpu.ALU.u_wallace._2839_ ;
 wire \u_cpu.ALU.u_wallace._2840_ ;
 wire \u_cpu.ALU.u_wallace._2841_ ;
 wire \u_cpu.ALU.u_wallace._2842_ ;
 wire \u_cpu.ALU.u_wallace._2843_ ;
 wire \u_cpu.ALU.u_wallace._2844_ ;
 wire \u_cpu.ALU.u_wallace._2845_ ;
 wire \u_cpu.ALU.u_wallace._2846_ ;
 wire \u_cpu.ALU.u_wallace._2847_ ;
 wire \u_cpu.ALU.u_wallace._2848_ ;
 wire \u_cpu.ALU.u_wallace._2849_ ;
 wire \u_cpu.ALU.u_wallace._2850_ ;
 wire \u_cpu.ALU.u_wallace._2851_ ;
 wire \u_cpu.ALU.u_wallace._2852_ ;
 wire \u_cpu.ALU.u_wallace._2853_ ;
 wire \u_cpu.ALU.u_wallace._2854_ ;
 wire \u_cpu.ALU.u_wallace._2855_ ;
 wire \u_cpu.ALU.u_wallace._2856_ ;
 wire \u_cpu.ALU.u_wallace._2857_ ;
 wire \u_cpu.ALU.u_wallace._2858_ ;
 wire \u_cpu.ALU.u_wallace._2859_ ;
 wire \u_cpu.ALU.u_wallace._2860_ ;
 wire \u_cpu.ALU.u_wallace._2861_ ;
 wire \u_cpu.ALU.u_wallace._2862_ ;
 wire \u_cpu.ALU.u_wallace._2863_ ;
 wire \u_cpu.ALU.u_wallace._2864_ ;
 wire \u_cpu.ALU.u_wallace._2865_ ;
 wire \u_cpu.ALU.u_wallace._2866_ ;
 wire \u_cpu.ALU.u_wallace._2867_ ;
 wire \u_cpu.ALU.u_wallace._2868_ ;
 wire \u_cpu.ALU.u_wallace._2869_ ;
 wire \u_cpu.ALU.u_wallace._2870_ ;
 wire \u_cpu.ALU.u_wallace._2871_ ;
 wire \u_cpu.ALU.u_wallace._2872_ ;
 wire \u_cpu.ALU.u_wallace._2873_ ;
 wire \u_cpu.ALU.u_wallace._2874_ ;
 wire \u_cpu.ALU.u_wallace._2875_ ;
 wire \u_cpu.ALU.u_wallace._2876_ ;
 wire \u_cpu.ALU.u_wallace._2877_ ;
 wire \u_cpu.ALU.u_wallace._2878_ ;
 wire \u_cpu.ALU.u_wallace._2879_ ;
 wire \u_cpu.ALU.u_wallace._2880_ ;
 wire \u_cpu.ALU.u_wallace._2881_ ;
 wire \u_cpu.ALU.u_wallace._2882_ ;
 wire \u_cpu.ALU.u_wallace._2883_ ;
 wire \u_cpu.ALU.u_wallace._2884_ ;
 wire \u_cpu.ALU.u_wallace._2885_ ;
 wire \u_cpu.ALU.u_wallace._2886_ ;
 wire \u_cpu.ALU.u_wallace._2887_ ;
 wire \u_cpu.ALU.u_wallace._2888_ ;
 wire \u_cpu.ALU.u_wallace._2889_ ;
 wire \u_cpu.ALU.u_wallace._2890_ ;
 wire \u_cpu.ALU.u_wallace._2891_ ;
 wire \u_cpu.ALU.u_wallace._2892_ ;
 wire \u_cpu.ALU.u_wallace._2893_ ;
 wire \u_cpu.ALU.u_wallace._2894_ ;
 wire \u_cpu.ALU.u_wallace._2895_ ;
 wire \u_cpu.ALU.u_wallace._2896_ ;
 wire \u_cpu.ALU.u_wallace._2897_ ;
 wire \u_cpu.ALU.u_wallace._2898_ ;
 wire \u_cpu.ALU.u_wallace._2899_ ;
 wire \u_cpu.ALU.u_wallace._2900_ ;
 wire \u_cpu.ALU.u_wallace._2901_ ;
 wire \u_cpu.ALU.u_wallace._2902_ ;
 wire \u_cpu.ALU.u_wallace._2903_ ;
 wire \u_cpu.ALU.u_wallace._2904_ ;
 wire \u_cpu.ALU.u_wallace._2905_ ;
 wire \u_cpu.ALU.u_wallace._2906_ ;
 wire \u_cpu.ALU.u_wallace._2907_ ;
 wire \u_cpu.ALU.u_wallace._2908_ ;
 wire \u_cpu.ALU.u_wallace._2909_ ;
 wire \u_cpu.ALU.u_wallace._2910_ ;
 wire \u_cpu.ALU.u_wallace._2911_ ;
 wire \u_cpu.ALU.u_wallace._2912_ ;
 wire \u_cpu.ALU.u_wallace._2913_ ;
 wire \u_cpu.ALU.u_wallace._2914_ ;
 wire \u_cpu.ALU.u_wallace._2915_ ;
 wire \u_cpu.ALU.u_wallace._2916_ ;
 wire \u_cpu.ALU.u_wallace._2917_ ;
 wire \u_cpu.ALU.u_wallace._2918_ ;
 wire \u_cpu.ALU.u_wallace._2919_ ;
 wire \u_cpu.ALU.u_wallace._2920_ ;
 wire \u_cpu.ALU.u_wallace._2921_ ;
 wire \u_cpu.ALU.u_wallace._2922_ ;
 wire \u_cpu.ALU.u_wallace._2923_ ;
 wire \u_cpu.ALU.u_wallace._2924_ ;
 wire \u_cpu.ALU.u_wallace._2925_ ;
 wire \u_cpu.ALU.u_wallace._2926_ ;
 wire \u_cpu.ALU.u_wallace._2927_ ;
 wire \u_cpu.ALU.u_wallace._2928_ ;
 wire \u_cpu.ALU.u_wallace._2929_ ;
 wire \u_cpu.ALU.u_wallace._2930_ ;
 wire \u_cpu.ALU.u_wallace._2931_ ;
 wire \u_cpu.ALU.u_wallace._2932_ ;
 wire \u_cpu.ALU.u_wallace._2933_ ;
 wire \u_cpu.ALU.u_wallace._2934_ ;
 wire \u_cpu.ALU.u_wallace._2935_ ;
 wire \u_cpu.ALU.u_wallace._2936_ ;
 wire \u_cpu.ALU.u_wallace._2937_ ;
 wire \u_cpu.ALU.u_wallace._2938_ ;
 wire \u_cpu.ALU.u_wallace._2939_ ;
 wire \u_cpu.ALU.u_wallace._2940_ ;
 wire \u_cpu.ALU.u_wallace._2941_ ;
 wire \u_cpu.ALU.u_wallace._2942_ ;
 wire \u_cpu.ALU.u_wallace._2943_ ;
 wire \u_cpu.ALU.u_wallace._2944_ ;
 wire \u_cpu.ALU.u_wallace._2945_ ;
 wire \u_cpu.ALU.u_wallace._2946_ ;
 wire \u_cpu.ALU.u_wallace._2947_ ;
 wire \u_cpu.ALU.u_wallace._2948_ ;
 wire \u_cpu.ALU.u_wallace._2949_ ;
 wire \u_cpu.ALU.u_wallace._2950_ ;
 wire \u_cpu.ALU.u_wallace._2951_ ;
 wire \u_cpu.ALU.u_wallace._2952_ ;
 wire \u_cpu.ALU.u_wallace._2953_ ;
 wire \u_cpu.ALU.u_wallace._2954_ ;
 wire \u_cpu.ALU.u_wallace._2955_ ;
 wire \u_cpu.ALU.u_wallace._2956_ ;
 wire \u_cpu.ALU.u_wallace._2957_ ;
 wire \u_cpu.ALU.u_wallace._2958_ ;
 wire \u_cpu.ALU.u_wallace._2959_ ;
 wire \u_cpu.ALU.u_wallace._2960_ ;
 wire \u_cpu.ALU.u_wallace._2961_ ;
 wire \u_cpu.ALU.u_wallace._2962_ ;
 wire \u_cpu.ALU.u_wallace._2963_ ;
 wire \u_cpu.ALU.u_wallace._2964_ ;
 wire \u_cpu.ALU.u_wallace._2965_ ;
 wire \u_cpu.ALU.u_wallace._2966_ ;
 wire \u_cpu.ALU.u_wallace._2967_ ;
 wire \u_cpu.ALU.u_wallace._2968_ ;
 wire \u_cpu.ALU.u_wallace._2969_ ;
 wire \u_cpu.ALU.u_wallace._2970_ ;
 wire \u_cpu.ALU.u_wallace._2971_ ;
 wire \u_cpu.ALU.u_wallace._2972_ ;
 wire \u_cpu.ALU.u_wallace._2973_ ;
 wire \u_cpu.ALU.u_wallace._2974_ ;
 wire \u_cpu.ALU.u_wallace._2975_ ;
 wire \u_cpu.ALU.u_wallace._2976_ ;
 wire \u_cpu.ALU.u_wallace._2977_ ;
 wire \u_cpu.ALU.u_wallace._2978_ ;
 wire \u_cpu.ALU.u_wallace._2979_ ;
 wire \u_cpu.ALU.u_wallace._2980_ ;
 wire \u_cpu.ALU.u_wallace._2981_ ;
 wire \u_cpu.ALU.u_wallace._2982_ ;
 wire \u_cpu.ALU.u_wallace._2983_ ;
 wire \u_cpu.ALU.u_wallace._2984_ ;
 wire \u_cpu.ALU.u_wallace._2985_ ;
 wire \u_cpu.ALU.u_wallace._2986_ ;
 wire \u_cpu.ALU.u_wallace._2987_ ;
 wire \u_cpu.ALU.u_wallace._2988_ ;
 wire \u_cpu.ALU.u_wallace._2989_ ;
 wire \u_cpu.ALU.u_wallace._2990_ ;
 wire \u_cpu.ALU.u_wallace._2991_ ;
 wire \u_cpu.ALU.u_wallace._2992_ ;
 wire \u_cpu.ALU.u_wallace._2993_ ;
 wire \u_cpu.ALU.u_wallace._2994_ ;
 wire \u_cpu.ALU.u_wallace._2995_ ;
 wire \u_cpu.ALU.u_wallace._2996_ ;
 wire \u_cpu.ALU.u_wallace._2997_ ;
 wire \u_cpu.ALU.u_wallace._2998_ ;
 wire \u_cpu.ALU.u_wallace._2999_ ;
 wire \u_cpu.ALU.u_wallace._3000_ ;
 wire \u_cpu.ALU.u_wallace._3001_ ;
 wire \u_cpu.ALU.u_wallace._3002_ ;
 wire \u_cpu.ALU.u_wallace._3003_ ;
 wire \u_cpu.ALU.u_wallace._3004_ ;
 wire \u_cpu.ALU.u_wallace._3005_ ;
 wire \u_cpu.ALU.u_wallace._3006_ ;
 wire \u_cpu.ALU.u_wallace._3007_ ;
 wire \u_cpu.ALU.u_wallace._3008_ ;
 wire \u_cpu.ALU.u_wallace._3009_ ;
 wire \u_cpu.ALU.u_wallace._3010_ ;
 wire \u_cpu.ALU.u_wallace._3011_ ;
 wire \u_cpu.ALU.u_wallace._3012_ ;
 wire \u_cpu.ALU.u_wallace._3013_ ;
 wire \u_cpu.ALU.u_wallace._3014_ ;
 wire \u_cpu.ALU.u_wallace._3015_ ;
 wire \u_cpu.ALU.u_wallace._3016_ ;
 wire \u_cpu.ALU.u_wallace._3017_ ;
 wire \u_cpu.ALU.u_wallace._3018_ ;
 wire \u_cpu.ALU.u_wallace._3019_ ;
 wire \u_cpu.ALU.u_wallace._3020_ ;
 wire \u_cpu.ALU.u_wallace._3021_ ;
 wire \u_cpu.ALU.u_wallace._3022_ ;
 wire \u_cpu.ALU.u_wallace._3023_ ;
 wire \u_cpu.ALU.u_wallace._3024_ ;
 wire \u_cpu.ALU.u_wallace._3025_ ;
 wire \u_cpu.ALU.u_wallace._3026_ ;
 wire \u_cpu.ALU.u_wallace._3027_ ;
 wire \u_cpu.ALU.u_wallace._3028_ ;
 wire \u_cpu.ALU.u_wallace._3029_ ;
 wire \u_cpu.ALU.u_wallace._3030_ ;
 wire \u_cpu.ALU.u_wallace._3031_ ;
 wire \u_cpu.ALU.u_wallace._3032_ ;
 wire \u_cpu.ALU.u_wallace._3033_ ;
 wire \u_cpu.ALU.u_wallace._3034_ ;
 wire \u_cpu.ALU.u_wallace._3035_ ;
 wire \u_cpu.ALU.u_wallace._3036_ ;
 wire \u_cpu.ALU.u_wallace._3037_ ;
 wire \u_cpu.ALU.u_wallace._3038_ ;
 wire \u_cpu.ALU.u_wallace._3039_ ;
 wire \u_cpu.ALU.u_wallace._3040_ ;
 wire \u_cpu.ALU.u_wallace._3041_ ;
 wire \u_cpu.ALU.u_wallace._3042_ ;
 wire \u_cpu.ALU.u_wallace._3043_ ;
 wire \u_cpu.ALU.u_wallace._3044_ ;
 wire \u_cpu.ALU.u_wallace._3045_ ;
 wire \u_cpu.ALU.u_wallace._3046_ ;
 wire \u_cpu.ALU.u_wallace._3047_ ;
 wire \u_cpu.ALU.u_wallace._3048_ ;
 wire \u_cpu.ALU.u_wallace._3049_ ;
 wire \u_cpu.ALU.u_wallace._3050_ ;
 wire \u_cpu.ALU.u_wallace._3051_ ;
 wire \u_cpu.ALU.u_wallace._3052_ ;
 wire \u_cpu.ALU.u_wallace._3053_ ;
 wire \u_cpu.ALU.u_wallace._3054_ ;
 wire \u_cpu.ALU.u_wallace._3055_ ;
 wire \u_cpu.ALU.u_wallace._3056_ ;
 wire \u_cpu.ALU.u_wallace._3057_ ;
 wire \u_cpu.ALU.u_wallace._3058_ ;
 wire \u_cpu.ALU.u_wallace._3059_ ;
 wire \u_cpu.ALU.u_wallace._3060_ ;
 wire \u_cpu.ALU.u_wallace._3061_ ;
 wire \u_cpu.ALU.u_wallace._3062_ ;
 wire \u_cpu.ALU.u_wallace._3063_ ;
 wire \u_cpu.ALU.u_wallace._3064_ ;
 wire \u_cpu.ALU.u_wallace._3065_ ;
 wire \u_cpu.ALU.u_wallace._3066_ ;
 wire \u_cpu.ALU.u_wallace._3067_ ;
 wire \u_cpu.ALU.u_wallace._3068_ ;
 wire \u_cpu.ALU.u_wallace._3069_ ;
 wire \u_cpu.ALU.u_wallace._3070_ ;
 wire \u_cpu.ALU.u_wallace._3071_ ;
 wire \u_cpu.ALU.u_wallace._3072_ ;
 wire \u_cpu.ALU.u_wallace._3073_ ;
 wire \u_cpu.ALU.u_wallace._3074_ ;
 wire \u_cpu.ALU.u_wallace._3075_ ;
 wire \u_cpu.ALU.u_wallace._3076_ ;
 wire \u_cpu.ALU.u_wallace._3077_ ;
 wire \u_cpu.ALU.u_wallace._3078_ ;
 wire \u_cpu.ALU.u_wallace._3079_ ;
 wire \u_cpu.ALU.u_wallace._3080_ ;
 wire \u_cpu.ALU.u_wallace._3081_ ;
 wire \u_cpu.ALU.u_wallace._3082_ ;
 wire \u_cpu.ALU.u_wallace._3083_ ;
 wire \u_cpu.ALU.u_wallace._3084_ ;
 wire \u_cpu.ALU.u_wallace._3085_ ;
 wire \u_cpu.ALU.u_wallace._3086_ ;
 wire \u_cpu.ALU.u_wallace._3087_ ;
 wire \u_cpu.ALU.u_wallace._3088_ ;
 wire \u_cpu.ALU.u_wallace._3089_ ;
 wire \u_cpu.ALU.u_wallace._3090_ ;
 wire \u_cpu.ALU.u_wallace._3091_ ;
 wire \u_cpu.ALU.u_wallace._3092_ ;
 wire \u_cpu.ALU.u_wallace._3093_ ;
 wire \u_cpu.ALU.u_wallace._3094_ ;
 wire \u_cpu.ALU.u_wallace._3095_ ;
 wire \u_cpu.ALU.u_wallace._3096_ ;
 wire \u_cpu.ALU.u_wallace._3097_ ;
 wire \u_cpu.ALU.u_wallace._3098_ ;
 wire \u_cpu.ALU.u_wallace._3099_ ;
 wire \u_cpu.ALU.u_wallace._3100_ ;
 wire \u_cpu.ALU.u_wallace._3101_ ;
 wire \u_cpu.ALU.u_wallace._3102_ ;
 wire \u_cpu.ALU.u_wallace._3103_ ;
 wire \u_cpu.ALU.u_wallace._3104_ ;
 wire \u_cpu.ALU.u_wallace._3105_ ;
 wire \u_cpu.ALU.u_wallace._3106_ ;
 wire \u_cpu.ALU.u_wallace._3107_ ;
 wire \u_cpu.ALU.u_wallace._3108_ ;
 wire \u_cpu.ALU.u_wallace._3109_ ;
 wire \u_cpu.ALU.u_wallace._3110_ ;
 wire \u_cpu.ALU.u_wallace._3111_ ;
 wire \u_cpu.ALU.u_wallace._3112_ ;
 wire \u_cpu.ALU.u_wallace._3113_ ;
 wire \u_cpu.ALU.u_wallace._3114_ ;
 wire \u_cpu.ALU.u_wallace._3115_ ;
 wire \u_cpu.ALU.u_wallace._3116_ ;
 wire \u_cpu.ALU.u_wallace._3117_ ;
 wire \u_cpu.ALU.u_wallace._3118_ ;
 wire \u_cpu.ALU.u_wallace._3119_ ;
 wire \u_cpu.ALU.u_wallace._3120_ ;
 wire \u_cpu.ALU.u_wallace._3121_ ;
 wire \u_cpu.ALU.u_wallace._3122_ ;
 wire \u_cpu.ALU.u_wallace._3123_ ;
 wire \u_cpu.ALU.u_wallace._3124_ ;
 wire \u_cpu.ALU.u_wallace._3125_ ;
 wire \u_cpu.ALU.u_wallace._3126_ ;
 wire \u_cpu.ALU.u_wallace._3127_ ;
 wire \u_cpu.ALU.u_wallace._3128_ ;
 wire \u_cpu.ALU.u_wallace._3129_ ;
 wire \u_cpu.ALU.u_wallace._3130_ ;
 wire \u_cpu.ALU.u_wallace._3131_ ;
 wire \u_cpu.ALU.u_wallace._3132_ ;
 wire \u_cpu.ALU.u_wallace._3133_ ;
 wire \u_cpu.ALU.u_wallace._3134_ ;
 wire \u_cpu.ALU.u_wallace._3135_ ;
 wire \u_cpu.ALU.u_wallace._3136_ ;
 wire \u_cpu.ALU.u_wallace._3137_ ;
 wire \u_cpu.ALU.u_wallace._3138_ ;
 wire \u_cpu.ALU.u_wallace._3139_ ;
 wire \u_cpu.ALU.u_wallace._3140_ ;
 wire \u_cpu.ALU.u_wallace._3141_ ;
 wire \u_cpu.ALU.u_wallace._3142_ ;
 wire \u_cpu.ALU.u_wallace._3143_ ;
 wire \u_cpu.ALU.u_wallace._3144_ ;
 wire \u_cpu.ALU.u_wallace._3145_ ;
 wire \u_cpu.ALU.u_wallace._3146_ ;
 wire \u_cpu.ALU.u_wallace._3147_ ;
 wire \u_cpu.ALU.u_wallace._3148_ ;
 wire \u_cpu.ALU.u_wallace._3149_ ;
 wire \u_cpu.ALU.u_wallace._3150_ ;
 wire \u_cpu.ALU.u_wallace._3151_ ;
 wire \u_cpu.ALU.u_wallace._3152_ ;
 wire \u_cpu.ALU.u_wallace._3153_ ;
 wire \u_cpu.ALU.u_wallace._3154_ ;
 wire \u_cpu.ALU.u_wallace._3155_ ;
 wire \u_cpu.ALU.u_wallace._3156_ ;
 wire \u_cpu.ALU.u_wallace._3157_ ;
 wire \u_cpu.ALU.u_wallace._3158_ ;
 wire \u_cpu.ALU.u_wallace._3159_ ;
 wire \u_cpu.ALU.u_wallace._3160_ ;
 wire \u_cpu.ALU.u_wallace._3161_ ;
 wire \u_cpu.ALU.u_wallace._3162_ ;
 wire \u_cpu.ALU.u_wallace._3163_ ;
 wire \u_cpu.ALU.u_wallace._3164_ ;
 wire \u_cpu.ALU.u_wallace._3165_ ;
 wire \u_cpu.ALU.u_wallace._3166_ ;
 wire \u_cpu.ALU.u_wallace._3167_ ;
 wire \u_cpu.ALU.u_wallace._3168_ ;
 wire \u_cpu.ALU.u_wallace._3169_ ;
 wire \u_cpu.ALU.u_wallace._3170_ ;
 wire \u_cpu.ALU.u_wallace._3171_ ;
 wire \u_cpu.ALU.u_wallace._3172_ ;
 wire \u_cpu.ALU.u_wallace._3173_ ;
 wire \u_cpu.ALU.u_wallace._3174_ ;
 wire \u_cpu.ALU.u_wallace._3175_ ;
 wire \u_cpu.ALU.u_wallace._3176_ ;
 wire \u_cpu.ALU.u_wallace._3177_ ;
 wire \u_cpu.ALU.u_wallace._3178_ ;
 wire \u_cpu.ALU.u_wallace._3179_ ;
 wire \u_cpu.ALU.u_wallace._3180_ ;
 wire \u_cpu.ALU.u_wallace._3181_ ;
 wire \u_cpu.ALU.u_wallace._3182_ ;
 wire \u_cpu.ALU.u_wallace._3183_ ;
 wire \u_cpu.ALU.u_wallace._3184_ ;
 wire \u_cpu.ALU.u_wallace._3185_ ;
 wire \u_cpu.ALU.u_wallace._3186_ ;
 wire \u_cpu.ALU.u_wallace._3187_ ;
 wire \u_cpu.ALU.u_wallace._3188_ ;
 wire \u_cpu.ALU.u_wallace._3189_ ;
 wire \u_cpu.ALU.u_wallace._3190_ ;
 wire \u_cpu.ALU.u_wallace._3191_ ;
 wire \u_cpu.ALU.u_wallace._3192_ ;
 wire \u_cpu.ALU.u_wallace._3193_ ;
 wire \u_cpu.ALU.u_wallace._3194_ ;
 wire \u_cpu.ALU.u_wallace._3195_ ;
 wire \u_cpu.ALU.u_wallace._3196_ ;
 wire \u_cpu.ALU.u_wallace._3197_ ;
 wire \u_cpu.ALU.u_wallace._3198_ ;
 wire \u_cpu.ALU.u_wallace._3199_ ;
 wire \u_cpu.ALU.u_wallace._3200_ ;
 wire \u_cpu.ALU.u_wallace._3201_ ;
 wire \u_cpu.ALU.u_wallace._3202_ ;
 wire \u_cpu.ALU.u_wallace._3203_ ;
 wire \u_cpu.ALU.u_wallace._3204_ ;
 wire \u_cpu.ALU.u_wallace._3205_ ;
 wire \u_cpu.ALU.u_wallace._3206_ ;
 wire \u_cpu.ALU.u_wallace._3207_ ;
 wire \u_cpu.ALU.u_wallace._3208_ ;
 wire \u_cpu.ALU.u_wallace._3209_ ;
 wire \u_cpu.ALU.u_wallace._3210_ ;
 wire \u_cpu.ALU.u_wallace._3211_ ;
 wire \u_cpu.ALU.u_wallace._3212_ ;
 wire \u_cpu.ALU.u_wallace._3213_ ;
 wire \u_cpu.ALU.u_wallace._3214_ ;
 wire \u_cpu.ALU.u_wallace._3215_ ;
 wire \u_cpu.ALU.u_wallace._3216_ ;
 wire \u_cpu.ALU.u_wallace._3217_ ;
 wire \u_cpu.ALU.u_wallace._3218_ ;
 wire \u_cpu.ALU.u_wallace._3219_ ;
 wire \u_cpu.ALU.u_wallace._3220_ ;
 wire \u_cpu.ALU.u_wallace._3221_ ;
 wire \u_cpu.ALU.u_wallace._3222_ ;
 wire \u_cpu.ALU.u_wallace._3223_ ;
 wire \u_cpu.ALU.u_wallace._3224_ ;
 wire \u_cpu.ALU.u_wallace._3225_ ;
 wire \u_cpu.ALU.u_wallace._3226_ ;
 wire \u_cpu.ALU.u_wallace._3227_ ;
 wire \u_cpu.ALU.u_wallace._3228_ ;
 wire \u_cpu.ALU.u_wallace._3229_ ;
 wire \u_cpu.ALU.u_wallace._3230_ ;
 wire \u_cpu.ALU.u_wallace._3231_ ;
 wire \u_cpu.ALU.u_wallace._3232_ ;
 wire \u_cpu.ALU.u_wallace._3233_ ;
 wire \u_cpu.ALU.u_wallace._3234_ ;
 wire \u_cpu.ALU.u_wallace._3235_ ;
 wire \u_cpu.ALU.u_wallace._3236_ ;
 wire \u_cpu.ALU.u_wallace._3237_ ;
 wire \u_cpu.ALU.u_wallace._3238_ ;
 wire \u_cpu.ALU.u_wallace._3239_ ;
 wire \u_cpu.ALU.u_wallace._3240_ ;
 wire \u_cpu.ALU.u_wallace._3241_ ;
 wire \u_cpu.ALU.u_wallace._3242_ ;
 wire \u_cpu.ALU.u_wallace._3243_ ;
 wire \u_cpu.ALU.u_wallace._3244_ ;
 wire \u_cpu.ALU.u_wallace._3245_ ;
 wire \u_cpu.ALU.u_wallace._3246_ ;
 wire \u_cpu.ALU.u_wallace._3247_ ;
 wire \u_cpu.ALU.u_wallace._3248_ ;
 wire \u_cpu.ALU.u_wallace._3249_ ;
 wire \u_cpu.ALU.u_wallace._3250_ ;
 wire \u_cpu.ALU.u_wallace._3251_ ;
 wire \u_cpu.ALU.u_wallace._3252_ ;
 wire \u_cpu.ALU.u_wallace._3253_ ;
 wire \u_cpu.ALU.u_wallace._3254_ ;
 wire \u_cpu.ALU.u_wallace._3255_ ;
 wire \u_cpu.ALU.u_wallace._3256_ ;
 wire \u_cpu.ALU.u_wallace._3257_ ;
 wire \u_cpu.ALU.u_wallace._3258_ ;
 wire \u_cpu.ALU.u_wallace._3259_ ;
 wire \u_cpu.ALU.u_wallace._3260_ ;
 wire \u_cpu.ALU.u_wallace._3261_ ;
 wire \u_cpu.ALU.u_wallace._3262_ ;
 wire \u_cpu.ALU.u_wallace._3263_ ;
 wire \u_cpu.ALU.u_wallace._3264_ ;
 wire \u_cpu.ALU.u_wallace._3265_ ;
 wire \u_cpu.ALU.u_wallace._3266_ ;
 wire \u_cpu.ALU.u_wallace._3267_ ;
 wire \u_cpu.ALU.u_wallace._3268_ ;
 wire \u_cpu.ALU.u_wallace._3269_ ;
 wire \u_cpu.ALU.u_wallace._3270_ ;
 wire \u_cpu.ALU.u_wallace._3271_ ;
 wire \u_cpu.ALU.u_wallace._3272_ ;
 wire \u_cpu.ALU.u_wallace._3273_ ;
 wire \u_cpu.ALU.u_wallace._3274_ ;
 wire \u_cpu.ALU.u_wallace._3275_ ;
 wire \u_cpu.ALU.u_wallace._3276_ ;
 wire \u_cpu.ALU.u_wallace._3277_ ;
 wire \u_cpu.ALU.u_wallace._3278_ ;
 wire \u_cpu.ALU.u_wallace._3279_ ;
 wire \u_cpu.ALU.u_wallace._3280_ ;
 wire \u_cpu.ALU.u_wallace._3281_ ;
 wire \u_cpu.ALU.u_wallace._3282_ ;
 wire \u_cpu.ALU.u_wallace._3283_ ;
 wire \u_cpu.ALU.u_wallace._3284_ ;
 wire \u_cpu.ALU.u_wallace._3285_ ;
 wire \u_cpu.ALU.u_wallace._3286_ ;
 wire \u_cpu.ALU.u_wallace._3287_ ;
 wire \u_cpu.ALU.u_wallace._3288_ ;
 wire \u_cpu.ALU.u_wallace._3289_ ;
 wire \u_cpu.ALU.u_wallace._3290_ ;
 wire \u_cpu.ALU.u_wallace._3291_ ;
 wire \u_cpu.ALU.u_wallace._3292_ ;
 wire \u_cpu.ALU.u_wallace._3293_ ;
 wire \u_cpu.ALU.u_wallace._3294_ ;
 wire \u_cpu.ALU.u_wallace._3295_ ;
 wire \u_cpu.ALU.u_wallace._3296_ ;
 wire \u_cpu.ALU.u_wallace._3297_ ;
 wire \u_cpu.ALU.u_wallace._3298_ ;
 wire \u_cpu.ALU.u_wallace._3299_ ;
 wire \u_cpu.ALU.u_wallace._3300_ ;
 wire \u_cpu.ALU.u_wallace._3301_ ;
 wire \u_cpu.ALU.u_wallace._3302_ ;
 wire \u_cpu.ALU.u_wallace._3303_ ;
 wire \u_cpu.ALU.u_wallace._3304_ ;
 wire \u_cpu.ALU.u_wallace._3305_ ;
 wire \u_cpu.ALU.u_wallace._3306_ ;
 wire \u_cpu.ALU.u_wallace._3307_ ;
 wire \u_cpu.ALU.u_wallace._3308_ ;
 wire \u_cpu.ALU.u_wallace._3309_ ;
 wire \u_cpu.ALU.u_wallace._3310_ ;
 wire \u_cpu.ALU.u_wallace._3311_ ;
 wire \u_cpu.ALU.u_wallace._3312_ ;
 wire \u_cpu.ALU.u_wallace._3313_ ;
 wire \u_cpu.ALU.u_wallace._3314_ ;
 wire \u_cpu.ALU.u_wallace._3315_ ;
 wire \u_cpu.ALU.u_wallace._3316_ ;
 wire \u_cpu.ALU.u_wallace._3317_ ;
 wire \u_cpu.ALU.u_wallace._3318_ ;
 wire \u_cpu.ALU.u_wallace._3319_ ;
 wire \u_cpu.ALU.u_wallace._3320_ ;
 wire \u_cpu.ALU.u_wallace._3321_ ;
 wire \u_cpu.ALU.u_wallace._3322_ ;
 wire \u_cpu.ALU.u_wallace._3323_ ;
 wire \u_cpu.ALU.u_wallace._3324_ ;
 wire \u_cpu.ALU.u_wallace._3325_ ;
 wire \u_cpu.ALU.u_wallace._3326_ ;
 wire \u_cpu.ALU.u_wallace._3327_ ;
 wire \u_cpu.ALU.u_wallace._3328_ ;
 wire \u_cpu.ALU.u_wallace._3329_ ;
 wire \u_cpu.ALU.u_wallace._3330_ ;
 wire \u_cpu.ALU.u_wallace._3331_ ;
 wire \u_cpu.ALU.u_wallace._3332_ ;
 wire \u_cpu.ALU.u_wallace._3333_ ;
 wire \u_cpu.ALU.u_wallace._3334_ ;
 wire \u_cpu.ALU.u_wallace._3335_ ;
 wire \u_cpu.ALU.u_wallace._3336_ ;
 wire \u_cpu.ALU.u_wallace._3337_ ;
 wire \u_cpu.ALU.u_wallace._3338_ ;
 wire \u_cpu.ALU.u_wallace._3339_ ;
 wire \u_cpu.ALU.u_wallace._3340_ ;
 wire \u_cpu.ALU.u_wallace._3341_ ;
 wire \u_cpu.ALU.u_wallace._3342_ ;
 wire \u_cpu.ALU.u_wallace._3343_ ;
 wire \u_cpu.ALU.u_wallace._3344_ ;
 wire \u_cpu.ALU.u_wallace._3345_ ;
 wire \u_cpu.ALU.u_wallace._3346_ ;
 wire \u_cpu.ALU.u_wallace._3347_ ;
 wire \u_cpu.ALU.u_wallace._3348_ ;
 wire \u_cpu.ALU.u_wallace._3349_ ;
 wire \u_cpu.ALU.u_wallace._3350_ ;
 wire \u_cpu.ALU.u_wallace._3351_ ;
 wire \u_cpu.ALU.u_wallace._3352_ ;
 wire \u_cpu.ALU.u_wallace._3353_ ;
 wire \u_cpu.ALU.u_wallace._3354_ ;
 wire \u_cpu.ALU.u_wallace._3355_ ;
 wire \u_cpu.ALU.u_wallace._3356_ ;
 wire \u_cpu.ALU.u_wallace._3357_ ;
 wire \u_cpu.ALU.u_wallace._3358_ ;
 wire \u_cpu.ALU.u_wallace._3359_ ;
 wire \u_cpu.ALU.u_wallace._3360_ ;
 wire \u_cpu.ALU.u_wallace._3361_ ;
 wire \u_cpu.ALU.u_wallace._3362_ ;
 wire \u_cpu.ALU.u_wallace._3363_ ;
 wire \u_cpu.ALU.u_wallace._3364_ ;
 wire \u_cpu.ALU.u_wallace._3365_ ;
 wire \u_cpu.ALU.u_wallace._3366_ ;
 wire \u_cpu.ALU.u_wallace._3367_ ;
 wire \u_cpu.ALU.u_wallace._3368_ ;
 wire \u_cpu.ALU.u_wallace._3369_ ;
 wire \u_cpu.ALU.u_wallace._3370_ ;
 wire \u_cpu.ALU.u_wallace._3371_ ;
 wire \u_cpu.ALU.u_wallace._3372_ ;
 wire \u_cpu.ALU.u_wallace._3373_ ;
 wire \u_cpu.ALU.u_wallace._3374_ ;
 wire \u_cpu.ALU.u_wallace._3375_ ;
 wire \u_cpu.ALU.u_wallace._3376_ ;
 wire \u_cpu.ALU.u_wallace._3377_ ;
 wire \u_cpu.ALU.u_wallace._3378_ ;
 wire \u_cpu.ALU.u_wallace._3379_ ;
 wire \u_cpu.ALU.u_wallace._3380_ ;
 wire \u_cpu.ALU.u_wallace._3381_ ;
 wire \u_cpu.ALU.u_wallace._3382_ ;
 wire \u_cpu.ALU.u_wallace._3383_ ;
 wire \u_cpu.ALU.u_wallace._3384_ ;
 wire \u_cpu.ALU.u_wallace._3385_ ;
 wire \u_cpu.ALU.u_wallace._3386_ ;
 wire \u_cpu.ALU.u_wallace._3387_ ;
 wire \u_cpu.ALU.u_wallace._3388_ ;
 wire \u_cpu.ALU.u_wallace._3389_ ;
 wire \u_cpu.ALU.u_wallace._3390_ ;
 wire \u_cpu.ALU.u_wallace._3391_ ;
 wire \u_cpu.ALU.u_wallace._3392_ ;
 wire \u_cpu.ALU.u_wallace._3393_ ;
 wire \u_cpu.ALU.u_wallace._3394_ ;
 wire \u_cpu.ALU.u_wallace._3395_ ;
 wire \u_cpu.ALU.u_wallace._3396_ ;
 wire \u_cpu.ALU.u_wallace._3397_ ;
 wire \u_cpu.ALU.u_wallace._3398_ ;
 wire \u_cpu.ALU.u_wallace._3399_ ;
 wire \u_cpu.ALU.u_wallace._3400_ ;
 wire \u_cpu.ALU.u_wallace._3401_ ;
 wire \u_cpu.ALU.u_wallace._3402_ ;
 wire \u_cpu.ALU.u_wallace._3403_ ;
 wire \u_cpu.ALU.u_wallace._3404_ ;
 wire \u_cpu.ALU.u_wallace._3405_ ;
 wire \u_cpu.ALU.u_wallace._3406_ ;
 wire \u_cpu.ALU.u_wallace._3407_ ;
 wire \u_cpu.ALU.u_wallace._3408_ ;
 wire \u_cpu.ALU.u_wallace._3409_ ;
 wire \u_cpu.ALU.u_wallace._3410_ ;
 wire \u_cpu.ALU.u_wallace._3411_ ;
 wire \u_cpu.ALU.u_wallace._3412_ ;
 wire \u_cpu.ALU.u_wallace._3413_ ;
 wire \u_cpu.ALU.u_wallace._3414_ ;
 wire \u_cpu.ALU.u_wallace._3415_ ;
 wire \u_cpu.ALU.u_wallace._3416_ ;
 wire \u_cpu.ALU.u_wallace._3417_ ;
 wire \u_cpu.ALU.u_wallace._3418_ ;
 wire \u_cpu.ALU.u_wallace._3419_ ;
 wire \u_cpu.ALU.u_wallace._3420_ ;
 wire \u_cpu.ALU.u_wallace._3421_ ;
 wire \u_cpu.ALU.u_wallace._3422_ ;
 wire \u_cpu.ALU.u_wallace._3423_ ;
 wire \u_cpu.ALU.u_wallace._3424_ ;
 wire \u_cpu.ALU.u_wallace._3425_ ;
 wire \u_cpu.ALU.u_wallace._3426_ ;
 wire \u_cpu.ALU.u_wallace._3427_ ;
 wire \u_cpu.ALU.u_wallace._3428_ ;
 wire \u_cpu.ALU.u_wallace._3429_ ;
 wire \u_cpu.ALU.u_wallace._3430_ ;
 wire \u_cpu.ALU.u_wallace._3431_ ;
 wire \u_cpu.ALU.u_wallace._3432_ ;
 wire \u_cpu.ALU.u_wallace._3433_ ;
 wire \u_cpu.ALU.u_wallace._3434_ ;
 wire \u_cpu.ALU.u_wallace._3435_ ;
 wire \u_cpu.ALU.u_wallace._3436_ ;
 wire \u_cpu.ALU.u_wallace._3437_ ;
 wire \u_cpu.ALU.u_wallace._3438_ ;
 wire \u_cpu.ALU.u_wallace._3439_ ;
 wire \u_cpu.ALU.u_wallace._3440_ ;
 wire \u_cpu.ALU.u_wallace._3441_ ;
 wire \u_cpu.ALU.u_wallace._3442_ ;
 wire \u_cpu.ALU.u_wallace._3443_ ;
 wire \u_cpu.ALU.u_wallace._3444_ ;
 wire \u_cpu.ALU.u_wallace._3445_ ;
 wire \u_cpu.ALU.u_wallace._3446_ ;
 wire \u_cpu.ALU.u_wallace._3447_ ;
 wire \u_cpu.ALU.u_wallace._3448_ ;
 wire \u_cpu.ALU.u_wallace._3449_ ;
 wire \u_cpu.ALU.u_wallace._3450_ ;
 wire \u_cpu.ALU.u_wallace._3451_ ;
 wire \u_cpu.ALU.u_wallace._3452_ ;
 wire \u_cpu.ALU.u_wallace._3453_ ;
 wire \u_cpu.ALU.u_wallace._3454_ ;
 wire \u_cpu.ALU.u_wallace._3455_ ;
 wire \u_cpu.ALU.u_wallace._3456_ ;
 wire \u_cpu.ALU.u_wallace._3457_ ;
 wire \u_cpu.ALU.u_wallace._3458_ ;
 wire \u_cpu.ALU.u_wallace._3459_ ;
 wire \u_cpu.ALU.u_wallace._3460_ ;
 wire \u_cpu.ALU.u_wallace._3461_ ;
 wire \u_cpu.ALU.u_wallace._3462_ ;
 wire \u_cpu.ALU.u_wallace._3463_ ;
 wire \u_cpu.ALU.u_wallace._3464_ ;
 wire \u_cpu.ALU.u_wallace._3465_ ;
 wire \u_cpu.ALU.u_wallace._3466_ ;
 wire \u_cpu.ALU.u_wallace._3467_ ;
 wire \u_cpu.ALU.u_wallace._3468_ ;
 wire \u_cpu.ALU.u_wallace._3469_ ;
 wire \u_cpu.ALU.u_wallace._3470_ ;
 wire \u_cpu.ALU.u_wallace._3471_ ;
 wire \u_cpu.ALU.u_wallace._3472_ ;
 wire \u_cpu.ALU.u_wallace._3473_ ;
 wire \u_cpu.ALU.u_wallace._3474_ ;
 wire \u_cpu.ALU.u_wallace._3475_ ;
 wire \u_cpu.ALU.u_wallace._3476_ ;
 wire \u_cpu.ALU.u_wallace._3477_ ;
 wire \u_cpu.ALU.u_wallace._3478_ ;
 wire \u_cpu.ALU.u_wallace._3479_ ;
 wire \u_cpu.ALU.u_wallace._3480_ ;
 wire \u_cpu.ALU.u_wallace._3481_ ;
 wire \u_cpu.ALU.u_wallace._3482_ ;
 wire \u_cpu.ALU.u_wallace._3483_ ;
 wire \u_cpu.ALU.u_wallace._3484_ ;
 wire \u_cpu.ALU.u_wallace._3485_ ;
 wire \u_cpu.ALU.u_wallace._3486_ ;
 wire \u_cpu.ALU.u_wallace._3487_ ;
 wire \u_cpu.ALU.u_wallace._3488_ ;
 wire \u_cpu.ALU.u_wallace._3489_ ;
 wire \u_cpu.ALU.u_wallace._3490_ ;
 wire \u_cpu.ALU.u_wallace._3491_ ;
 wire \u_cpu.ALU.u_wallace._3492_ ;
 wire \u_cpu.ALU.u_wallace._3493_ ;
 wire \u_cpu.ALU.u_wallace._3494_ ;
 wire \u_cpu.ALU.u_wallace._3495_ ;
 wire \u_cpu.ALU.u_wallace._3496_ ;
 wire \u_cpu.ALU.u_wallace._3497_ ;
 wire \u_cpu.ALU.u_wallace._3498_ ;
 wire \u_cpu.ALU.u_wallace._3499_ ;
 wire \u_cpu.ALU.u_wallace._3500_ ;
 wire \u_cpu.ALU.u_wallace._3501_ ;
 wire \u_cpu.ALU.u_wallace._3502_ ;
 wire \u_cpu.ALU.u_wallace._3503_ ;
 wire \u_cpu.ALU.u_wallace._3504_ ;
 wire \u_cpu.ALU.u_wallace._3505_ ;
 wire \u_cpu.ALU.u_wallace._3506_ ;
 wire \u_cpu.ALU.u_wallace._3507_ ;
 wire \u_cpu.ALU.u_wallace._3508_ ;
 wire \u_cpu.ALU.u_wallace._3509_ ;
 wire \u_cpu.ALU.u_wallace._3510_ ;
 wire \u_cpu.ALU.u_wallace._3511_ ;
 wire \u_cpu.ALU.u_wallace._3512_ ;
 wire \u_cpu.ALU.u_wallace._3513_ ;
 wire \u_cpu.ALU.u_wallace._3514_ ;
 wire \u_cpu.ALU.u_wallace._3515_ ;
 wire \u_cpu.ALU.u_wallace._3516_ ;
 wire \u_cpu.ALU.u_wallace._3517_ ;
 wire \u_cpu.ALU.u_wallace._3518_ ;
 wire \u_cpu.ALU.u_wallace._3519_ ;
 wire \u_cpu.ALU.u_wallace._3520_ ;
 wire \u_cpu.ALU.u_wallace._3521_ ;
 wire \u_cpu.ALU.u_wallace._3522_ ;
 wire \u_cpu.ALU.u_wallace._3523_ ;
 wire \u_cpu.ALU.u_wallace._3524_ ;
 wire \u_cpu.ALU.u_wallace._3525_ ;
 wire \u_cpu.ALU.u_wallace._3526_ ;
 wire \u_cpu.ALU.u_wallace._3527_ ;
 wire \u_cpu.ALU.u_wallace._3528_ ;
 wire \u_cpu.ALU.u_wallace._3529_ ;
 wire \u_cpu.ALU.u_wallace._3530_ ;
 wire \u_cpu.ALU.u_wallace._3531_ ;
 wire \u_cpu.ALU.u_wallace._3532_ ;
 wire \u_cpu.ALU.u_wallace._3533_ ;
 wire \u_cpu.ALU.u_wallace._3534_ ;
 wire \u_cpu.ALU.u_wallace._3535_ ;
 wire \u_cpu.ALU.u_wallace._3536_ ;
 wire \u_cpu.ALU.u_wallace._3537_ ;
 wire \u_cpu.ALU.u_wallace._3538_ ;
 wire \u_cpu.ALU.u_wallace._3539_ ;
 wire \u_cpu.ALU.u_wallace._3540_ ;
 wire \u_cpu.ALU.u_wallace._3541_ ;
 wire \u_cpu.ALU.u_wallace._3542_ ;
 wire \u_cpu.ALU.u_wallace._3543_ ;
 wire \u_cpu.ALU.u_wallace._3544_ ;
 wire \u_cpu.ALU.u_wallace._3545_ ;
 wire \u_cpu.ALU.u_wallace._3546_ ;
 wire \u_cpu.ALU.u_wallace._3547_ ;
 wire \u_cpu.ALU.u_wallace._3548_ ;
 wire \u_cpu.ALU.u_wallace._3549_ ;
 wire \u_cpu.ALU.u_wallace._3550_ ;
 wire \u_cpu.ALU.u_wallace._3551_ ;
 wire \u_cpu.ALU.u_wallace._3552_ ;
 wire \u_cpu.ALU.u_wallace._3553_ ;
 wire \u_cpu.ALU.u_wallace._3554_ ;
 wire \u_cpu.ALU.u_wallace._3555_ ;
 wire \u_cpu.ALU.u_wallace._3556_ ;
 wire \u_cpu.ALU.u_wallace._3557_ ;
 wire \u_cpu.ALU.u_wallace._3558_ ;
 wire \u_cpu.ALU.u_wallace._3559_ ;
 wire \u_cpu.ALU.u_wallace._3560_ ;
 wire \u_cpu.ALU.u_wallace._3561_ ;
 wire \u_cpu.ALU.u_wallace._3562_ ;
 wire \u_cpu.ALU.u_wallace._3563_ ;
 wire \u_cpu.ALU.u_wallace._3564_ ;
 wire \u_cpu.ALU.u_wallace._3565_ ;
 wire \u_cpu.ALU.u_wallace._3566_ ;
 wire \u_cpu.ALU.u_wallace._3567_ ;
 wire \u_cpu.ALU.u_wallace._3568_ ;
 wire \u_cpu.ALU.u_wallace._3569_ ;
 wire \u_cpu.ALU.u_wallace._3570_ ;
 wire \u_cpu.ALU.u_wallace._3571_ ;
 wire \u_cpu.ALU.u_wallace._3572_ ;
 wire \u_cpu.ALU.u_wallace._3573_ ;
 wire \u_cpu.ALU.u_wallace._3574_ ;
 wire \u_cpu.ALU.u_wallace._3575_ ;
 wire \u_cpu.ALU.u_wallace._3576_ ;
 wire \u_cpu.ALU.u_wallace._3577_ ;
 wire \u_cpu.ALU.u_wallace._3578_ ;
 wire \u_cpu.ALU.u_wallace._3579_ ;
 wire \u_cpu.ALU.u_wallace._3580_ ;
 wire \u_cpu.ALU.u_wallace._3581_ ;
 wire \u_cpu.ALU.u_wallace._3582_ ;
 wire \u_cpu.ALU.u_wallace._3583_ ;
 wire \u_cpu.ALU.u_wallace._3584_ ;
 wire \u_cpu.ALU.u_wallace._3585_ ;
 wire \u_cpu.ALU.u_wallace._3586_ ;
 wire \u_cpu.ALU.u_wallace._3587_ ;
 wire \u_cpu.ALU.u_wallace._3588_ ;
 wire \u_cpu.ALU.u_wallace._3589_ ;
 wire \u_cpu.ALU.u_wallace._3590_ ;
 wire \u_cpu.ALU.u_wallace._3591_ ;
 wire \u_cpu.ALU.u_wallace._3592_ ;
 wire \u_cpu.ALU.u_wallace._3593_ ;
 wire \u_cpu.ALU.u_wallace._3594_ ;
 wire \u_cpu.ALU.u_wallace._3595_ ;
 wire \u_cpu.ALU.u_wallace._3596_ ;
 wire \u_cpu.ALU.u_wallace._3597_ ;
 wire \u_cpu.ALU.u_wallace._3598_ ;
 wire \u_cpu.ALU.u_wallace._3599_ ;
 wire \u_cpu.ALU.u_wallace._3600_ ;
 wire \u_cpu.ALU.u_wallace._3601_ ;
 wire \u_cpu.ALU.u_wallace._3602_ ;
 wire \u_cpu.ALU.u_wallace._3603_ ;
 wire \u_cpu.ALU.u_wallace._3604_ ;
 wire \u_cpu.ALU.u_wallace._3605_ ;
 wire \u_cpu.ALU.u_wallace._3606_ ;
 wire \u_cpu.ALU.u_wallace._3607_ ;
 wire \u_cpu.ALU.u_wallace._3608_ ;
 wire \u_cpu.ALU.u_wallace._3609_ ;
 wire \u_cpu.ALU.u_wallace._3610_ ;
 wire \u_cpu.ALU.u_wallace._3611_ ;
 wire \u_cpu.ALU.u_wallace._3612_ ;
 wire \u_cpu.ALU.u_wallace._3613_ ;
 wire \u_cpu.ALU.u_wallace._3614_ ;
 wire \u_cpu.ALU.u_wallace._3615_ ;
 wire \u_cpu.ALU.u_wallace._3616_ ;
 wire \u_cpu.ALU.u_wallace._3617_ ;
 wire \u_cpu.ALU.u_wallace._3618_ ;
 wire \u_cpu.ALU.u_wallace._3619_ ;
 wire \u_cpu.ALU.u_wallace._3620_ ;
 wire \u_cpu.ALU.u_wallace._3621_ ;
 wire \u_cpu.ALU.u_wallace._3622_ ;
 wire \u_cpu.ALU.u_wallace._3623_ ;
 wire \u_cpu.ALU.u_wallace._3624_ ;
 wire \u_cpu.ALU.u_wallace._3625_ ;
 wire \u_cpu.ALU.u_wallace._3626_ ;
 wire \u_cpu.ALU.u_wallace._3627_ ;
 wire \u_cpu.ALU.u_wallace._3628_ ;
 wire \u_cpu.ALU.u_wallace._3629_ ;
 wire \u_cpu.ALU.u_wallace._3630_ ;
 wire \u_cpu.ALU.u_wallace._3631_ ;
 wire \u_cpu.ALU.u_wallace._3632_ ;
 wire \u_cpu.ALU.u_wallace._3633_ ;
 wire \u_cpu.ALU.u_wallace._3634_ ;
 wire \u_cpu.ALU.u_wallace._3635_ ;
 wire \u_cpu.ALU.u_wallace._3636_ ;
 wire \u_cpu.ALU.u_wallace._3637_ ;
 wire \u_cpu.ALU.u_wallace._3638_ ;
 wire \u_cpu.ALU.u_wallace._3639_ ;
 wire \u_cpu.ALU.u_wallace._3640_ ;
 wire \u_cpu.ALU.u_wallace._3641_ ;
 wire \u_cpu.ALU.u_wallace._3642_ ;
 wire \u_cpu.ALU.u_wallace._3643_ ;
 wire \u_cpu.ALU.u_wallace._3644_ ;
 wire \u_cpu.ALU.u_wallace._3645_ ;
 wire \u_cpu.ALU.u_wallace._3646_ ;
 wire \u_cpu.ALU.u_wallace._3647_ ;
 wire \u_cpu.ALU.u_wallace._3648_ ;
 wire \u_cpu.ALU.u_wallace._3649_ ;
 wire \u_cpu.ALU.u_wallace._3650_ ;
 wire \u_cpu.ALU.u_wallace._3651_ ;
 wire \u_cpu.ALU.u_wallace._3652_ ;
 wire \u_cpu.ALU.u_wallace._3653_ ;
 wire \u_cpu.ALU.u_wallace._3654_ ;
 wire \u_cpu.ALU.u_wallace._3655_ ;
 wire \u_cpu.ALU.u_wallace._3656_ ;
 wire \u_cpu.ALU.u_wallace._3657_ ;
 wire \u_cpu.ALU.u_wallace._3658_ ;
 wire \u_cpu.ALU.u_wallace._3659_ ;
 wire \u_cpu.ALU.u_wallace._3660_ ;
 wire \u_cpu.ALU.u_wallace._3661_ ;
 wire \u_cpu.ALU.u_wallace._3662_ ;
 wire \u_cpu.ALU.u_wallace._3663_ ;
 wire \u_cpu.ALU.u_wallace._3664_ ;
 wire \u_cpu.ALU.u_wallace._3665_ ;
 wire \u_cpu.ALU.u_wallace._3666_ ;
 wire \u_cpu.ALU.u_wallace._3667_ ;
 wire \u_cpu.ALU.u_wallace._3668_ ;
 wire \u_cpu.ALU.u_wallace._3669_ ;
 wire \u_cpu.ALU.u_wallace._3670_ ;
 wire \u_cpu.ALU.u_wallace._3671_ ;
 wire \u_cpu.ALU.u_wallace._3672_ ;
 wire \u_cpu.ALU.u_wallace._3673_ ;
 wire \u_cpu.ALU.u_wallace._3674_ ;
 wire \u_cpu.ALU.u_wallace._3675_ ;
 wire \u_cpu.ALU.u_wallace._3676_ ;
 wire \u_cpu.ALU.u_wallace._3677_ ;
 wire \u_cpu.ALU.u_wallace._3678_ ;
 wire \u_cpu.ALU.u_wallace._3679_ ;
 wire \u_cpu.ALU.u_wallace._3680_ ;
 wire \u_cpu.ALU.u_wallace._3681_ ;
 wire \u_cpu.ALU.u_wallace._3682_ ;
 wire \u_cpu.ALU.u_wallace._3683_ ;
 wire \u_cpu.ALU.u_wallace._3684_ ;
 wire \u_cpu.ALU.u_wallace._3685_ ;
 wire \u_cpu.ALU.u_wallace._3686_ ;
 wire \u_cpu.ALU.u_wallace._3687_ ;
 wire \u_cpu.ALU.u_wallace._3688_ ;
 wire \u_cpu.ALU.u_wallace._3689_ ;
 wire \u_cpu.ALU.u_wallace._3690_ ;
 wire \u_cpu.ALU.u_wallace._3691_ ;
 wire \u_cpu.ALU.u_wallace._3692_ ;
 wire \u_cpu.ALU.u_wallace._3693_ ;
 wire \u_cpu.ALU.u_wallace._3694_ ;
 wire \u_cpu.ALU.u_wallace._3695_ ;
 wire \u_cpu.ALU.u_wallace._3696_ ;
 wire \u_cpu.ALU.u_wallace._3697_ ;
 wire \u_cpu.ALU.u_wallace._3698_ ;
 wire \u_cpu.ALU.u_wallace._3699_ ;
 wire \u_cpu.ALU.u_wallace._3700_ ;
 wire \u_cpu.ALU.u_wallace._3701_ ;
 wire \u_cpu.ALU.u_wallace._3702_ ;
 wire \u_cpu.ALU.u_wallace._3703_ ;
 wire \u_cpu.ALU.u_wallace._3704_ ;
 wire \u_cpu.ALU.u_wallace._3705_ ;
 wire \u_cpu.ALU.u_wallace._3706_ ;
 wire \u_cpu.ALU.u_wallace._3707_ ;
 wire \u_cpu.ALU.u_wallace._3708_ ;
 wire \u_cpu.ALU.u_wallace._3709_ ;
 wire \u_cpu.ALU.u_wallace._3710_ ;
 wire \u_cpu.ALU.u_wallace._3711_ ;
 wire \u_cpu.ALU.u_wallace._3712_ ;
 wire \u_cpu.ALU.u_wallace._3713_ ;
 wire \u_cpu.ALU.u_wallace._3714_ ;
 wire \u_cpu.ALU.u_wallace._3715_ ;
 wire \u_cpu.ALU.u_wallace._3716_ ;
 wire \u_cpu.ALU.u_wallace._3717_ ;
 wire \u_cpu.ALU.u_wallace._3718_ ;
 wire \u_cpu.ALU.u_wallace._3719_ ;
 wire \u_cpu.ALU.u_wallace._3720_ ;
 wire \u_cpu.ALU.u_wallace._3721_ ;
 wire \u_cpu.ALU.u_wallace._3722_ ;
 wire \u_cpu.ALU.u_wallace._3723_ ;
 wire \u_cpu.ALU.u_wallace._3724_ ;
 wire \u_cpu.ALU.u_wallace._3725_ ;
 wire \u_cpu.ALU.u_wallace._3726_ ;
 wire \u_cpu.ALU.u_wallace._3727_ ;
 wire \u_cpu.ALU.u_wallace._3728_ ;
 wire \u_cpu.ALU.u_wallace._3729_ ;
 wire \u_cpu.ALU.u_wallace._3730_ ;
 wire \u_cpu.ALU.u_wallace._3731_ ;
 wire \u_cpu.ALU.u_wallace._3732_ ;
 wire \u_cpu.ALU.u_wallace._3733_ ;
 wire \u_cpu.ALU.u_wallace._3734_ ;
 wire \u_cpu.ALU.u_wallace._3735_ ;
 wire \u_cpu.ALU.u_wallace._3736_ ;
 wire \u_cpu.ALU.u_wallace._3737_ ;
 wire \u_cpu.ALU.u_wallace._3738_ ;
 wire \u_cpu.ALU.u_wallace._3739_ ;
 wire \u_cpu.ALU.u_wallace._3740_ ;
 wire \u_cpu.ALU.u_wallace._3741_ ;
 wire \u_cpu.ALU.u_wallace._3742_ ;
 wire \u_cpu.ALU.u_wallace._3743_ ;
 wire \u_cpu.ALU.u_wallace._3744_ ;
 wire \u_cpu.ALU.u_wallace._3745_ ;
 wire \u_cpu.ALU.u_wallace._3746_ ;
 wire \u_cpu.ALU.u_wallace._3747_ ;
 wire \u_cpu.ALU.u_wallace._3748_ ;
 wire \u_cpu.ALU.u_wallace._3749_ ;
 wire \u_cpu.ALU.u_wallace._3750_ ;
 wire \u_cpu.ALU.u_wallace._3751_ ;
 wire \u_cpu.ALU.u_wallace._3752_ ;
 wire \u_cpu.ALU.u_wallace._3753_ ;
 wire \u_cpu.ALU.u_wallace._3754_ ;
 wire \u_cpu.ALU.u_wallace._3755_ ;
 wire \u_cpu.ALU.u_wallace._3756_ ;
 wire \u_cpu.ALU.u_wallace._3757_ ;
 wire \u_cpu.ALU.u_wallace._3758_ ;
 wire \u_cpu.ALU.u_wallace._3759_ ;
 wire \u_cpu.ALU.u_wallace._3760_ ;
 wire \u_cpu.ALU.u_wallace._3761_ ;
 wire \u_cpu.ALU.u_wallace._3762_ ;
 wire \u_cpu.ALU.u_wallace._3763_ ;
 wire \u_cpu.ALU.u_wallace._3764_ ;
 wire \u_cpu.ALU.u_wallace._3765_ ;
 wire \u_cpu.ALU.u_wallace._3766_ ;
 wire \u_cpu.ALU.u_wallace._3767_ ;
 wire \u_cpu.ALU.u_wallace._3768_ ;
 wire \u_cpu.ALU.u_wallace._3769_ ;
 wire \u_cpu.ALU.u_wallace._3770_ ;
 wire \u_cpu.ALU.u_wallace._3771_ ;
 wire \u_cpu.ALU.u_wallace._3772_ ;
 wire \u_cpu.ALU.u_wallace._3773_ ;
 wire \u_cpu.ALU.u_wallace._3774_ ;
 wire \u_cpu.ALU.u_wallace._3775_ ;
 wire \u_cpu.ALU.u_wallace._3776_ ;
 wire \u_cpu.ALU.u_wallace._3777_ ;
 wire \u_cpu.ALU.u_wallace._3778_ ;
 wire \u_cpu.ALU.u_wallace._3779_ ;
 wire \u_cpu.ALU.u_wallace._3780_ ;
 wire \u_cpu.ALU.u_wallace._3781_ ;
 wire \u_cpu.ALU.u_wallace._3782_ ;
 wire \u_cpu.ALU.u_wallace._3783_ ;
 wire \u_cpu.ALU.u_wallace._3784_ ;
 wire \u_cpu.ALU.u_wallace._3785_ ;
 wire \u_cpu.ALU.u_wallace._3786_ ;
 wire \u_cpu.ALU.u_wallace._3787_ ;
 wire \u_cpu.ALU.u_wallace._3788_ ;
 wire \u_cpu.ALU.u_wallace._3789_ ;
 wire \u_cpu.ALU.u_wallace._3790_ ;
 wire \u_cpu.ALU.u_wallace._3791_ ;
 wire \u_cpu.ALU.u_wallace._3792_ ;
 wire \u_cpu.ALU.u_wallace._3793_ ;
 wire \u_cpu.ALU.u_wallace._3794_ ;
 wire \u_cpu.ALU.u_wallace._3795_ ;
 wire \u_cpu.ALU.u_wallace._3796_ ;
 wire \u_cpu.ALU.u_wallace._3797_ ;
 wire \u_cpu.ALU.u_wallace._3798_ ;
 wire \u_cpu.ALU.u_wallace._3799_ ;
 wire \u_cpu.ALU.u_wallace._3800_ ;
 wire \u_cpu.ALU.u_wallace._3801_ ;
 wire \u_cpu.ALU.u_wallace._3802_ ;
 wire \u_cpu.ALU.u_wallace._3803_ ;
 wire \u_cpu.ALU.u_wallace._3804_ ;
 wire \u_cpu.ALU.u_wallace._3805_ ;
 wire \u_cpu.ALU.u_wallace._3806_ ;
 wire \u_cpu.ALU.u_wallace._3807_ ;
 wire \u_cpu.ALU.u_wallace._3808_ ;
 wire \u_cpu.ALU.u_wallace._3809_ ;
 wire \u_cpu.ALU.u_wallace._3810_ ;
 wire \u_cpu.ALU.u_wallace._3811_ ;
 wire \u_cpu.ALU.u_wallace._3812_ ;
 wire \u_cpu.ALU.u_wallace._3813_ ;
 wire \u_cpu.ALU.u_wallace._3814_ ;
 wire \u_cpu.ALU.u_wallace._3815_ ;
 wire \u_cpu.ALU.u_wallace._3816_ ;
 wire \u_cpu.ALU.u_wallace._3817_ ;
 wire \u_cpu.ALU.u_wallace._3818_ ;
 wire \u_cpu.ALU.u_wallace._3819_ ;
 wire \u_cpu.ALU.u_wallace._3820_ ;
 wire \u_cpu.ALU.u_wallace._3821_ ;
 wire \u_cpu.ALU.u_wallace._3822_ ;
 wire \u_cpu.ALU.u_wallace._3823_ ;
 wire \u_cpu.ALU.u_wallace._3824_ ;
 wire \u_cpu.ALU.u_wallace._3825_ ;
 wire \u_cpu.ALU.u_wallace._3826_ ;
 wire \u_cpu.ALU.u_wallace._3827_ ;
 wire \u_cpu.ALU.u_wallace._3828_ ;
 wire \u_cpu.ALU.u_wallace._3829_ ;
 wire \u_cpu.ALU.u_wallace._3830_ ;
 wire \u_cpu.ALU.u_wallace._3831_ ;
 wire \u_cpu.ALU.u_wallace._3832_ ;
 wire \u_cpu.ALU.u_wallace._3833_ ;
 wire \u_cpu.ALU.u_wallace._3834_ ;
 wire \u_cpu.ALU.u_wallace._3835_ ;
 wire \u_cpu.ALU.u_wallace._3836_ ;
 wire \u_cpu.ALU.u_wallace._3837_ ;
 wire \u_cpu.ALU.u_wallace._3838_ ;
 wire \u_cpu.ALU.u_wallace._3839_ ;
 wire \u_cpu.ALU.u_wallace._3840_ ;
 wire \u_cpu.ALU.u_wallace._3841_ ;
 wire \u_cpu.ALU.u_wallace._3842_ ;
 wire \u_cpu.ALU.u_wallace._3843_ ;
 wire \u_cpu.ALU.u_wallace._3844_ ;
 wire \u_cpu.ALU.u_wallace._3845_ ;
 wire \u_cpu.ALU.u_wallace._3846_ ;
 wire \u_cpu.ALU.u_wallace._3847_ ;
 wire \u_cpu.ALU.u_wallace._3848_ ;
 wire \u_cpu.ALU.u_wallace._3849_ ;
 wire \u_cpu.ALU.u_wallace._3850_ ;
 wire \u_cpu.ALU.u_wallace._3851_ ;
 wire \u_cpu.ALU.u_wallace._3852_ ;
 wire \u_cpu.ALU.u_wallace._3853_ ;
 wire \u_cpu.ALU.u_wallace._3854_ ;
 wire \u_cpu.ALU.u_wallace._3855_ ;
 wire \u_cpu.ALU.u_wallace._3856_ ;
 wire \u_cpu.ALU.u_wallace._3857_ ;
 wire \u_cpu.ALU.u_wallace._3858_ ;
 wire \u_cpu.ALU.u_wallace._3859_ ;
 wire \u_cpu.ALU.u_wallace._3860_ ;
 wire \u_cpu.ALU.u_wallace._3861_ ;
 wire \u_cpu.ALU.u_wallace._3862_ ;
 wire \u_cpu.ALU.u_wallace._3863_ ;
 wire \u_cpu.ALU.u_wallace._3864_ ;
 wire \u_cpu.ALU.u_wallace._3865_ ;
 wire \u_cpu.ALU.u_wallace._3866_ ;
 wire \u_cpu.ALU.u_wallace._3867_ ;
 wire \u_cpu.ALU.u_wallace._3868_ ;
 wire \u_cpu.ALU.u_wallace._3869_ ;
 wire \u_cpu.ALU.u_wallace._3870_ ;
 wire \u_cpu.ALU.u_wallace._3871_ ;
 wire \u_cpu.ALU.u_wallace._3872_ ;
 wire \u_cpu.ALU.u_wallace._3873_ ;
 wire \u_cpu.ALU.u_wallace._3874_ ;
 wire \u_cpu.ALU.u_wallace._3875_ ;
 wire \u_cpu.ALU.u_wallace._3876_ ;
 wire \u_cpu.ALU.u_wallace._3877_ ;
 wire \u_cpu.ALU.u_wallace._3878_ ;
 wire \u_cpu.ALU.u_wallace._3879_ ;
 wire \u_cpu.ALU.u_wallace._3880_ ;
 wire \u_cpu.ALU.u_wallace._3881_ ;
 wire \u_cpu.ALU.u_wallace._3882_ ;
 wire \u_cpu.ALU.u_wallace._3883_ ;
 wire \u_cpu.ALU.u_wallace._3884_ ;
 wire \u_cpu.ALU.u_wallace._3885_ ;
 wire \u_cpu.ALU.u_wallace._3886_ ;
 wire \u_cpu.ALU.u_wallace._3887_ ;
 wire \u_cpu.ALU.u_wallace._3888_ ;
 wire \u_cpu.ALU.u_wallace._3889_ ;
 wire \u_cpu.ALU.u_wallace._3890_ ;
 wire \u_cpu.ALU.u_wallace._3891_ ;
 wire \u_cpu.ALU.u_wallace._3892_ ;
 wire \u_cpu.ALU.u_wallace._3893_ ;
 wire \u_cpu.ALU.u_wallace._3894_ ;
 wire \u_cpu.ALU.u_wallace._3895_ ;
 wire \u_cpu.ALU.u_wallace._3896_ ;
 wire \u_cpu.ALU.u_wallace._3897_ ;
 wire \u_cpu.ALU.u_wallace._3898_ ;
 wire \u_cpu.ALU.u_wallace._3899_ ;
 wire \u_cpu.ALU.u_wallace._3900_ ;
 wire \u_cpu.ALU.u_wallace._3901_ ;
 wire \u_cpu.ALU.u_wallace._3902_ ;
 wire \u_cpu.ALU.u_wallace._3903_ ;
 wire \u_cpu.ALU.u_wallace._3904_ ;
 wire \u_cpu.ALU.u_wallace._3905_ ;
 wire \u_cpu.ALU.u_wallace._3906_ ;
 wire \u_cpu.ALU.u_wallace._3907_ ;
 wire \u_cpu.ALU.u_wallace._3908_ ;
 wire \u_cpu.ALU.u_wallace._3909_ ;
 wire \u_cpu.ALU.u_wallace._3910_ ;
 wire \u_cpu.ALU.u_wallace._3911_ ;
 wire \u_cpu.ALU.u_wallace._3912_ ;
 wire \u_cpu.ALU.u_wallace._3913_ ;
 wire \u_cpu.ALU.u_wallace._3914_ ;
 wire \u_cpu.ALU.u_wallace._3915_ ;
 wire \u_cpu.ALU.u_wallace._3916_ ;
 wire \u_cpu.ALU.u_wallace._3917_ ;
 wire \u_cpu.ALU.u_wallace._3918_ ;
 wire \u_cpu.ALU.u_wallace._3919_ ;
 wire \u_cpu.ALU.u_wallace._3920_ ;
 wire \u_cpu.ALU.u_wallace._3921_ ;
 wire \u_cpu.ALU.u_wallace._3922_ ;
 wire \u_cpu.ALU.u_wallace._3923_ ;
 wire \u_cpu.ALU.u_wallace._3924_ ;
 wire \u_cpu.ALU.u_wallace._3925_ ;
 wire \u_cpu.ALU.u_wallace._3926_ ;
 wire \u_cpu.ALU.u_wallace._3927_ ;
 wire \u_cpu.ALU.u_wallace._3928_ ;
 wire \u_cpu.ALU.u_wallace._3929_ ;
 wire \u_cpu.ALU.u_wallace._3930_ ;
 wire \u_cpu.ALU.u_wallace._3931_ ;
 wire \u_cpu.ALU.u_wallace._3932_ ;
 wire \u_cpu.ALU.u_wallace._3933_ ;
 wire \u_cpu.ALU.u_wallace._3934_ ;
 wire \u_cpu.ALU.u_wallace._3935_ ;
 wire \u_cpu.ALU.u_wallace._3936_ ;
 wire \u_cpu.ALU.u_wallace._3937_ ;
 wire \u_cpu.ALU.u_wallace._3938_ ;
 wire \u_cpu.ALU.u_wallace._3939_ ;
 wire \u_cpu.ALU.u_wallace._3940_ ;
 wire \u_cpu.ALU.u_wallace._3941_ ;
 wire \u_cpu.ALU.u_wallace._3942_ ;
 wire \u_cpu.ALU.u_wallace._3943_ ;
 wire \u_cpu.ALU.u_wallace._3944_ ;
 wire \u_cpu.ALU.u_wallace._3945_ ;
 wire \u_cpu.ALU.u_wallace._3946_ ;
 wire \u_cpu.ALU.u_wallace._3947_ ;
 wire \u_cpu.ALU.u_wallace._3948_ ;
 wire \u_cpu.ALU.u_wallace._3949_ ;
 wire \u_cpu.ALU.u_wallace._3950_ ;
 wire \u_cpu.ALU.u_wallace._3951_ ;
 wire \u_cpu.ALU.u_wallace._3952_ ;
 wire \u_cpu.ALU.u_wallace._3953_ ;
 wire \u_cpu.ALU.u_wallace._3954_ ;
 wire \u_cpu.ALU.u_wallace._3955_ ;
 wire \u_cpu.ALU.u_wallace._3956_ ;
 wire \u_cpu.ALU.u_wallace._3957_ ;
 wire \u_cpu.ALU.u_wallace._3958_ ;
 wire \u_cpu.ALU.u_wallace._3959_ ;
 wire \u_cpu.ALU.u_wallace._3960_ ;
 wire \u_cpu.ALU.u_wallace._3961_ ;
 wire \u_cpu.ALU.u_wallace._3962_ ;
 wire \u_cpu.ALU.u_wallace._3963_ ;
 wire \u_cpu.ALU.u_wallace._3964_ ;
 wire \u_cpu.ALU.u_wallace._3965_ ;
 wire \u_cpu.ALU.u_wallace._3966_ ;
 wire \u_cpu.ALU.u_wallace._3967_ ;
 wire \u_cpu.ALU.u_wallace._3968_ ;
 wire \u_cpu.ALU.u_wallace._3969_ ;
 wire \u_cpu.ALU.u_wallace._3970_ ;
 wire \u_cpu.ALU.u_wallace._3971_ ;
 wire \u_cpu.ALU.u_wallace._3972_ ;
 wire \u_cpu.ALU.u_wallace._3973_ ;
 wire \u_cpu.ALU.u_wallace._3974_ ;
 wire \u_cpu.ALU.u_wallace._3975_ ;
 wire \u_cpu.ALU.u_wallace._3976_ ;
 wire \u_cpu.ALU.u_wallace._3977_ ;
 wire \u_cpu.ALU.u_wallace._3978_ ;
 wire \u_cpu.ALU.u_wallace._3979_ ;
 wire \u_cpu.ALU.u_wallace._3980_ ;
 wire \u_cpu.ALU.u_wallace._3981_ ;
 wire \u_cpu.ALU.u_wallace._3982_ ;
 wire \u_cpu.ALU.u_wallace._3983_ ;
 wire \u_cpu.ALU.u_wallace._3984_ ;
 wire \u_cpu.ALU.u_wallace._3985_ ;
 wire \u_cpu.ALU.u_wallace._3986_ ;
 wire \u_cpu.ALU.u_wallace._3987_ ;
 wire \u_cpu.ALU.u_wallace._3988_ ;
 wire \u_cpu.ALU.u_wallace._3989_ ;
 wire \u_cpu.ALU.u_wallace._3990_ ;
 wire \u_cpu.ALU.u_wallace._3991_ ;
 wire \u_cpu.ALU.u_wallace._3992_ ;
 wire \u_cpu.ALU.u_wallace._3993_ ;
 wire \u_cpu.ALU.u_wallace._3994_ ;
 wire \u_cpu.ALU.u_wallace._3995_ ;
 wire \u_cpu.ALU.u_wallace._3996_ ;
 wire \u_cpu.ALU.u_wallace._3997_ ;
 wire \u_cpu.ALU.u_wallace._3998_ ;
 wire \u_cpu.ALU.u_wallace._3999_ ;
 wire \u_cpu.ALU.u_wallace._4000_ ;
 wire \u_cpu.ALU.u_wallace._4001_ ;
 wire \u_cpu.ALU.u_wallace._4002_ ;
 wire \u_cpu.ALU.u_wallace._4003_ ;
 wire \u_cpu.ALU.u_wallace._4004_ ;
 wire \u_cpu.ALU.u_wallace._4005_ ;
 wire \u_cpu.ALU.u_wallace._4006_ ;
 wire \u_cpu.ALU.u_wallace._4007_ ;
 wire \u_cpu.ALU.u_wallace._4008_ ;
 wire \u_cpu.ALU.u_wallace._4009_ ;
 wire \u_cpu.ALU.u_wallace._4010_ ;
 wire \u_cpu.ALU.u_wallace._4011_ ;
 wire \u_cpu.ALU.u_wallace._4012_ ;
 wire \u_cpu.ALU.u_wallace._4013_ ;
 wire \u_cpu.ALU.u_wallace._4014_ ;
 wire \u_cpu.ALU.u_wallace._4015_ ;
 wire \u_cpu.ALU.u_wallace._4016_ ;
 wire \u_cpu.ALU.u_wallace._4017_ ;
 wire \u_cpu.ALU.u_wallace._4018_ ;
 wire \u_cpu.ALU.u_wallace._4019_ ;
 wire \u_cpu.ALU.u_wallace._4020_ ;
 wire \u_cpu.ALU.u_wallace._4021_ ;
 wire \u_cpu.ALU.u_wallace._4022_ ;
 wire \u_cpu.ALU.u_wallace._4023_ ;
 wire \u_cpu.ALU.u_wallace._4024_ ;
 wire \u_cpu.ALU.u_wallace._4025_ ;
 wire \u_cpu.ALU.u_wallace._4026_ ;
 wire \u_cpu.ALU.u_wallace._4027_ ;
 wire \u_cpu.ALU.u_wallace._4028_ ;
 wire \u_cpu.ALU.u_wallace._4029_ ;
 wire \u_cpu.ALU.u_wallace._4030_ ;
 wire \u_cpu.ALU.u_wallace._4031_ ;
 wire \u_cpu.ALU.u_wallace._4032_ ;
 wire \u_cpu.ALU.u_wallace._4033_ ;
 wire \u_cpu.ALU.u_wallace._4034_ ;
 wire \u_cpu.ALU.u_wallace._4035_ ;
 wire \u_cpu.ALU.u_wallace._4036_ ;
 wire \u_cpu.ALU.u_wallace._4037_ ;
 wire \u_cpu.ALU.u_wallace._4038_ ;
 wire \u_cpu.ALU.u_wallace._4039_ ;
 wire \u_cpu.ALU.u_wallace._4040_ ;
 wire \u_cpu.ALU.u_wallace._4041_ ;
 wire \u_cpu.ALU.u_wallace._4042_ ;
 wire \u_cpu.ALU.u_wallace._4043_ ;
 wire \u_cpu.ALU.u_wallace._4044_ ;
 wire \u_cpu.ALU.u_wallace._4045_ ;
 wire \u_cpu.ALU.u_wallace._4046_ ;
 wire \u_cpu.ALU.u_wallace._4047_ ;
 wire \u_cpu.ALU.u_wallace._4048_ ;
 wire \u_cpu.ALU.u_wallace._4049_ ;
 wire \u_cpu.ALU.u_wallace._4050_ ;
 wire \u_cpu.ALU.u_wallace._4051_ ;
 wire \u_cpu.ALU.u_wallace._4052_ ;
 wire \u_cpu.ALU.u_wallace._4053_ ;
 wire \u_cpu.ALU.u_wallace._4054_ ;
 wire \u_cpu.ALU.u_wallace._4055_ ;
 wire \u_cpu.ALU.u_wallace._4056_ ;
 wire \u_cpu.ALU.u_wallace._4057_ ;
 wire \u_cpu.ALU.u_wallace._4058_ ;
 wire \u_cpu.ALU.u_wallace._4059_ ;
 wire \u_cpu.ALU.u_wallace._4060_ ;
 wire \u_cpu.ALU.u_wallace._4061_ ;
 wire \u_cpu.ALU.u_wallace._4062_ ;
 wire \u_cpu.ALU.u_wallace._4063_ ;
 wire \u_cpu.ALU.u_wallace._4064_ ;
 wire \u_cpu.ALU.u_wallace._4065_ ;
 wire \u_cpu.ALU.u_wallace._4066_ ;
 wire \u_cpu.ALU.u_wallace._4067_ ;
 wire \u_cpu.ALU.u_wallace._4068_ ;
 wire \u_cpu.ALU.u_wallace._4069_ ;
 wire \u_cpu.ALU.u_wallace._4070_ ;
 wire \u_cpu.ALU.u_wallace._4071_ ;
 wire \u_cpu.ALU.u_wallace._4072_ ;
 wire \u_cpu.ALU.u_wallace._4073_ ;
 wire \u_cpu.ALU.u_wallace._4074_ ;
 wire \u_cpu.ALU.u_wallace._4075_ ;
 wire \u_cpu.ALU.u_wallace._4076_ ;
 wire \u_cpu.ALU.u_wallace._4077_ ;
 wire \u_cpu.ALU.u_wallace._4078_ ;
 wire \u_cpu.ALU.u_wallace._4079_ ;
 wire \u_cpu.ALU.u_wallace._4080_ ;
 wire \u_cpu.ALU.u_wallace._4081_ ;
 wire \u_cpu.ALU.u_wallace._4082_ ;
 wire \u_cpu.ALU.u_wallace._4083_ ;
 wire \u_cpu.ALU.u_wallace._4084_ ;
 wire \u_cpu.ALU.u_wallace._4085_ ;
 wire \u_cpu.ALU.u_wallace._4086_ ;
 wire \u_cpu.ALU.u_wallace._4087_ ;
 wire \u_cpu.ALU.u_wallace._4088_ ;
 wire \u_cpu.ALU.u_wallace._4089_ ;
 wire \u_cpu.ALU.u_wallace._4090_ ;
 wire \u_cpu.ALU.u_wallace._4091_ ;
 wire \u_cpu.ALU.u_wallace._4092_ ;
 wire \u_cpu.ALU.u_wallace._4093_ ;
 wire \u_cpu.ALU.u_wallace._4094_ ;
 wire \u_cpu.ALU.u_wallace._4095_ ;
 wire \u_cpu.ALU.u_wallace._4096_ ;
 wire \u_cpu.ALU.u_wallace._4097_ ;
 wire \u_cpu.ALU.u_wallace._4098_ ;
 wire \u_cpu.ALU.u_wallace._4099_ ;
 wire \u_cpu.ALU.u_wallace._4100_ ;
 wire \u_cpu.ALU.u_wallace._4101_ ;
 wire \u_cpu.ALU.u_wallace._4102_ ;
 wire \u_cpu.ALU.u_wallace._4103_ ;
 wire \u_cpu.ALU.u_wallace._4104_ ;
 wire \u_cpu.ALU.u_wallace._4105_ ;
 wire \u_cpu.ALU.u_wallace._4106_ ;
 wire \u_cpu.ALU.u_wallace._4107_ ;
 wire \u_cpu.ALU.u_wallace._4108_ ;
 wire \u_cpu.ALU.u_wallace._4109_ ;
 wire \u_cpu.ALU.u_wallace._4110_ ;
 wire \u_cpu.ALU.u_wallace._4111_ ;
 wire \u_cpu.ALU.u_wallace._4112_ ;
 wire \u_cpu.ALU.u_wallace._4113_ ;
 wire \u_cpu.ALU.u_wallace._4114_ ;
 wire \u_cpu.ALU.u_wallace._4115_ ;
 wire \u_cpu.ALU.u_wallace._4116_ ;
 wire \u_cpu.ALU.u_wallace._4117_ ;
 wire \u_cpu.ALU.u_wallace._4118_ ;
 wire \u_cpu.ALU.u_wallace._4119_ ;
 wire \u_cpu.ALU.u_wallace._4120_ ;
 wire \u_cpu.ALU.u_wallace._4121_ ;
 wire \u_cpu.ALU.u_wallace._4122_ ;
 wire \u_cpu.ALU.u_wallace._4123_ ;
 wire \u_cpu.ALU.u_wallace._4124_ ;
 wire \u_cpu.ALU.u_wallace._4125_ ;
 wire \u_cpu.ALU.u_wallace._4126_ ;
 wire \u_cpu.ALU.u_wallace._4127_ ;
 wire \u_cpu.ALU.u_wallace._4128_ ;
 wire \u_cpu.ALU.u_wallace._4129_ ;
 wire \u_cpu.ALU.u_wallace._4130_ ;
 wire \u_cpu.ALU.u_wallace._4131_ ;
 wire \u_cpu.ALU.u_wallace._4132_ ;
 wire \u_cpu.ALU.u_wallace._4133_ ;
 wire \u_cpu.ALU.u_wallace._4134_ ;
 wire \u_cpu.ALU.u_wallace._4135_ ;
 wire \u_cpu.ALU.u_wallace._4136_ ;
 wire \u_cpu.ALU.u_wallace._4137_ ;
 wire \u_cpu.ALU.u_wallace._4138_ ;
 wire \u_cpu.ALU.u_wallace._4139_ ;
 wire \u_cpu.ALU.u_wallace._4140_ ;
 wire \u_cpu.ALU.u_wallace._4141_ ;
 wire \u_cpu.ALU.u_wallace._4142_ ;
 wire \u_cpu.ALU.u_wallace._4143_ ;
 wire \u_cpu.ALU.u_wallace._4144_ ;
 wire \u_cpu.ALU.u_wallace._4145_ ;
 wire \u_cpu.ALU.u_wallace._4146_ ;
 wire \u_cpu.ALU.u_wallace._4147_ ;
 wire \u_cpu.ALU.u_wallace._4148_ ;
 wire \u_cpu.ALU.u_wallace._4149_ ;
 wire \u_cpu.ALU.u_wallace._4150_ ;
 wire \u_cpu.ALU.u_wallace._4151_ ;
 wire \u_cpu.ALU.u_wallace._4152_ ;
 wire \u_cpu.ALU.u_wallace._4153_ ;
 wire \u_cpu.ALU.u_wallace._4154_ ;
 wire \u_cpu.ALU.u_wallace._4155_ ;
 wire \u_cpu.ALU.u_wallace._4156_ ;
 wire \u_cpu.ALU.u_wallace._4157_ ;
 wire \u_cpu.ALU.u_wallace._4158_ ;
 wire \u_cpu.ALU.u_wallace._4159_ ;
 wire \u_cpu.ALU.u_wallace._4160_ ;
 wire \u_cpu.ALU.u_wallace._4161_ ;
 wire \u_cpu.ALU.u_wallace._4162_ ;
 wire \u_cpu.ALU.u_wallace._4163_ ;
 wire \u_cpu.ALU.u_wallace._4164_ ;
 wire \u_cpu.ALU.u_wallace._4165_ ;
 wire \u_cpu.ALU.u_wallace._4166_ ;
 wire \u_cpu.ALU.u_wallace._4167_ ;
 wire \u_cpu.ALU.u_wallace._4168_ ;
 wire \u_cpu.ALU.u_wallace._4169_ ;
 wire \u_cpu.ALU.u_wallace._4170_ ;
 wire \u_cpu.ALU.u_wallace._4171_ ;
 wire \u_cpu.ALU.u_wallace._4172_ ;
 wire \u_cpu.ALU.u_wallace._4173_ ;
 wire \u_cpu.ALU.u_wallace._4174_ ;
 wire \u_cpu.ALU.u_wallace._4175_ ;
 wire \u_cpu.ALU.u_wallace._4176_ ;
 wire \u_cpu.ALU.u_wallace._4177_ ;
 wire \u_cpu.ALU.u_wallace._4178_ ;
 wire \u_cpu.ALU.u_wallace._4179_ ;
 wire \u_cpu.ALU.u_wallace._4180_ ;
 wire \u_cpu.ALU.u_wallace._4181_ ;
 wire \u_cpu.ALU.u_wallace._4182_ ;
 wire \u_cpu.ALU.u_wallace._4183_ ;
 wire \u_cpu.ALU.u_wallace._4184_ ;
 wire \u_cpu.ALU.u_wallace._4185_ ;
 wire \u_cpu.ALU.u_wallace._4186_ ;
 wire \u_cpu.ALU.u_wallace._4187_ ;
 wire \u_cpu.ALU.u_wallace._4188_ ;
 wire \u_cpu.ALU.u_wallace._4189_ ;
 wire \u_cpu.ALU.u_wallace._4190_ ;
 wire \u_cpu.ALU.u_wallace._4191_ ;
 wire \u_cpu.ALU.u_wallace._4192_ ;
 wire \u_cpu.ALU.u_wallace._4193_ ;
 wire \u_cpu.ALU.u_wallace._4194_ ;
 wire \u_cpu.ALU.u_wallace._4195_ ;
 wire \u_cpu.ALU.u_wallace._4196_ ;
 wire \u_cpu.ALU.u_wallace._4197_ ;
 wire \u_cpu.ALU.u_wallace._4198_ ;
 wire \u_cpu.ALU.u_wallace._4199_ ;
 wire \u_cpu.ALU.u_wallace._4200_ ;
 wire \u_cpu.ALU.u_wallace._4201_ ;
 wire \u_cpu.ALU.u_wallace._4202_ ;
 wire \u_cpu.ALU.u_wallace._4203_ ;
 wire \u_cpu.ALU.u_wallace._4204_ ;
 wire \u_cpu.ALU.u_wallace._4205_ ;
 wire \u_cpu.ALU.u_wallace._4206_ ;
 wire \u_cpu.ALU.u_wallace._4207_ ;
 wire \u_cpu.ALU.u_wallace._4208_ ;
 wire \u_cpu.ALU.u_wallace._4209_ ;
 wire \u_cpu.ALU.u_wallace._4210_ ;
 wire \u_cpu.ALU.u_wallace._4211_ ;
 wire \u_cpu.ALU.u_wallace._4212_ ;
 wire \u_cpu.ALU.u_wallace._4213_ ;
 wire \u_cpu.ALU.u_wallace._4214_ ;
 wire \u_cpu.ALU.u_wallace._4215_ ;
 wire \u_cpu.ALU.u_wallace._4216_ ;
 wire \u_cpu.ALU.u_wallace._4217_ ;
 wire \u_cpu.ALU.u_wallace._4218_ ;
 wire \u_cpu.ALU.u_wallace._4219_ ;
 wire \u_cpu.ALU.u_wallace._4220_ ;
 wire \u_cpu.ALU.u_wallace._4221_ ;
 wire \u_cpu.ALU.u_wallace._4222_ ;
 wire \u_cpu.ALU.u_wallace._4223_ ;
 wire \u_cpu.ALU.u_wallace._4224_ ;
 wire \u_cpu.ALU.u_wallace._4225_ ;
 wire \u_cpu.ALU.u_wallace._4226_ ;
 wire \u_cpu.ALU.u_wallace._4227_ ;
 wire \u_cpu.ALU.u_wallace._4228_ ;
 wire \u_cpu.ALU.u_wallace._4229_ ;
 wire \u_cpu.ALU.u_wallace._4230_ ;
 wire \u_cpu.ALU.u_wallace._4231_ ;
 wire \u_cpu.ALU.u_wallace._4232_ ;
 wire \u_cpu.ALU.u_wallace._4233_ ;
 wire \u_cpu.ALU.u_wallace._4234_ ;
 wire \u_cpu.ALU.u_wallace._4235_ ;
 wire \u_cpu.ALU.u_wallace._4236_ ;
 wire \u_cpu.ALU.u_wallace._4237_ ;
 wire \u_cpu.ALU.u_wallace._4238_ ;
 wire \u_cpu.ALU.u_wallace._4239_ ;
 wire \u_cpu.ALU.u_wallace._4240_ ;
 wire \u_cpu.ALU.u_wallace._4241_ ;
 wire \u_cpu.ALU.u_wallace._4242_ ;
 wire \u_cpu.ALU.u_wallace._4243_ ;
 wire \u_cpu.ALU.u_wallace._4244_ ;
 wire \u_cpu.ALU.u_wallace._4245_ ;
 wire \u_cpu.ALU.u_wallace._4246_ ;
 wire \u_cpu.ALU.u_wallace._4247_ ;
 wire \u_cpu.ALU.u_wallace._4248_ ;
 wire \u_cpu.ALU.u_wallace._4249_ ;
 wire \u_cpu.ALU.u_wallace._4250_ ;
 wire \u_cpu.ALU.u_wallace._4251_ ;
 wire \u_cpu.ALU.u_wallace._4252_ ;
 wire \u_cpu.ALU.u_wallace._4253_ ;
 wire \u_cpu.ALU.u_wallace._4254_ ;
 wire \u_cpu.ALU.u_wallace._4255_ ;
 wire \u_cpu.ALU.u_wallace._4256_ ;
 wire \u_cpu.ALU.u_wallace._4257_ ;
 wire \u_cpu.ALU.u_wallace._4258_ ;
 wire \u_cpu.ALU.u_wallace._4259_ ;
 wire \u_cpu.ALU.u_wallace._4260_ ;
 wire \u_cpu.ALU.u_wallace._4261_ ;
 wire \u_cpu.ALU.u_wallace._4262_ ;
 wire \u_cpu.ALU.u_wallace._4263_ ;
 wire \u_cpu.ALU.u_wallace._4264_ ;
 wire \u_cpu.ALU.u_wallace._4265_ ;
 wire \u_cpu.ALU.u_wallace._4266_ ;
 wire \u_cpu.ALU.u_wallace._4267_ ;
 wire \u_cpu.ALU.u_wallace._4268_ ;
 wire \u_cpu.ALU.u_wallace._4269_ ;
 wire \u_cpu.ALU.u_wallace._4270_ ;
 wire \u_cpu.ALU.u_wallace._4271_ ;
 wire \u_cpu.ALU.u_wallace._4272_ ;
 wire \u_cpu.ALU.u_wallace._4273_ ;
 wire \u_cpu.ALU.u_wallace._4274_ ;
 wire \u_cpu.ALU.u_wallace._4275_ ;
 wire \u_cpu.ALU.u_wallace._4276_ ;
 wire \u_cpu.ALU.u_wallace._4277_ ;
 wire \u_cpu.ALU.u_wallace._4278_ ;
 wire \u_cpu.ALU.u_wallace._4279_ ;
 wire \u_cpu.ALU.u_wallace._4280_ ;
 wire \u_cpu.ALU.u_wallace._4281_ ;
 wire \u_cpu.ALU.u_wallace._4282_ ;
 wire \u_cpu.ALU.u_wallace._4283_ ;
 wire \u_cpu.ALU.u_wallace._4284_ ;
 wire \u_cpu.ALU.u_wallace._4285_ ;
 wire \u_cpu.ALU.u_wallace._4286_ ;
 wire \u_cpu.ALU.u_wallace._4287_ ;
 wire \u_cpu.ALU.u_wallace._4288_ ;
 wire \u_cpu.ALU.u_wallace._4289_ ;
 wire \u_cpu.ALU.u_wallace._4290_ ;
 wire \u_cpu.ALU.u_wallace._4291_ ;
 wire \u_cpu.ALU.u_wallace._4292_ ;
 wire \u_cpu.ALU.u_wallace._4293_ ;
 wire \u_cpu.ALU.u_wallace._4294_ ;
 wire \u_cpu.ALU.u_wallace._4295_ ;
 wire \u_cpu.ALU.u_wallace._4296_ ;
 wire \u_cpu.ALU.u_wallace._4297_ ;
 wire \u_cpu.ALU.u_wallace._4298_ ;
 wire \u_cpu.ALU.u_wallace._4299_ ;
 wire \u_cpu.ALU.u_wallace._4300_ ;
 wire \u_cpu.ALU.u_wallace._4301_ ;
 wire \u_cpu.ALU.u_wallace._4302_ ;
 wire \u_cpu.ALU.u_wallace._4303_ ;
 wire \u_cpu.ALU.u_wallace._4304_ ;
 wire \u_cpu.ALU.u_wallace._4305_ ;
 wire \u_cpu.ALU.u_wallace._4306_ ;
 wire \u_cpu.ALU.u_wallace._4307_ ;
 wire \u_cpu.ALU.u_wallace._4308_ ;
 wire \u_cpu.ALU.u_wallace._4309_ ;
 wire \u_cpu.ALU.u_wallace._4310_ ;
 wire \u_cpu.ALU.u_wallace._4311_ ;
 wire \u_cpu.ALU.u_wallace._4312_ ;
 wire \u_cpu.ALU.u_wallace._4313_ ;
 wire \u_cpu.ALU.u_wallace._4314_ ;
 wire \u_cpu.ALU.u_wallace._4315_ ;
 wire \u_cpu.ALU.u_wallace._4316_ ;
 wire \u_cpu.ALU.u_wallace._4317_ ;
 wire \u_cpu.ALU.u_wallace._4318_ ;
 wire \u_cpu.ALU.u_wallace._4319_ ;
 wire \u_cpu.ALU.u_wallace._4320_ ;
 wire \u_cpu.ALU.u_wallace._4321_ ;
 wire \u_cpu.ALU.u_wallace._4322_ ;
 wire \u_cpu.ALU.u_wallace._4323_ ;
 wire \u_cpu.ALU.u_wallace._4324_ ;
 wire \u_cpu.ALU.u_wallace._4325_ ;
 wire \u_cpu.ALU.u_wallace._4326_ ;
 wire \u_cpu.ALU.u_wallace._4327_ ;
 wire \u_cpu.ALU.u_wallace._4328_ ;
 wire \u_cpu.ALU.u_wallace._4329_ ;
 wire \u_cpu.ALU.u_wallace._4330_ ;
 wire \u_cpu.ALU.u_wallace._4331_ ;
 wire \u_cpu.ALU.u_wallace._4332_ ;
 wire \u_cpu.ALU.u_wallace._4333_ ;
 wire \u_cpu.ALU.u_wallace._4334_ ;
 wire \u_cpu.ALU.u_wallace._4335_ ;
 wire \u_cpu.ALU.u_wallace._4336_ ;
 wire \u_cpu.ALU.u_wallace._4337_ ;
 wire \u_cpu.ALU.u_wallace._4338_ ;
 wire \u_cpu.ALU.u_wallace._4339_ ;
 wire \u_cpu.ALU.u_wallace._4340_ ;
 wire \u_cpu.ALU.u_wallace._4341_ ;
 wire \u_cpu.ALU.u_wallace._4342_ ;
 wire \u_cpu.ALU.u_wallace._4343_ ;
 wire \u_cpu.ALU.u_wallace._4344_ ;
 wire \u_cpu.ALU.u_wallace._4345_ ;
 wire \u_cpu.ALU.u_wallace._4346_ ;
 wire \u_cpu.ALU.u_wallace._4347_ ;
 wire \u_cpu.ALU.u_wallace._4348_ ;
 wire \u_cpu.ALU.u_wallace._4349_ ;
 wire \u_cpu.ALU.u_wallace._4350_ ;
 wire \u_cpu.ALU.u_wallace._4351_ ;
 wire \u_cpu.ALU.u_wallace._4352_ ;
 wire \u_cpu.ALU.u_wallace._4353_ ;
 wire \u_cpu.ALU.u_wallace._4354_ ;
 wire \u_cpu.ALU.u_wallace._4355_ ;
 wire \u_cpu.ALU.u_wallace._4356_ ;
 wire \u_cpu.ALU.u_wallace._4357_ ;
 wire \u_cpu.ALU.u_wallace._4358_ ;
 wire \u_cpu.ALU.u_wallace._4359_ ;
 wire \u_cpu.ALU.u_wallace._4360_ ;
 wire \u_cpu.ALU.u_wallace._4361_ ;
 wire \u_cpu.ALU.u_wallace._4362_ ;
 wire \u_cpu.ALU.u_wallace._4363_ ;
 wire \u_cpu.ALU.u_wallace._4364_ ;
 wire \u_cpu.ALU.u_wallace._4365_ ;
 wire \u_cpu.ALU.u_wallace._4366_ ;
 wire \u_cpu.ALU.u_wallace._4367_ ;
 wire \u_cpu.ALU.u_wallace._4368_ ;
 wire \u_cpu.ALU.u_wallace._4369_ ;
 wire \u_cpu.ALU.u_wallace._4370_ ;
 wire \u_cpu.ALU.u_wallace._4371_ ;
 wire \u_cpu.ALU.u_wallace._4372_ ;
 wire \u_cpu.ALU.u_wallace._4373_ ;
 wire \u_cpu.ALU.u_wallace._4374_ ;
 wire \u_cpu.ALU.u_wallace._4375_ ;
 wire \u_cpu.ALU.u_wallace._4376_ ;
 wire \u_cpu.ALU.u_wallace._4377_ ;
 wire \u_cpu.ALU.u_wallace._4378_ ;
 wire \u_cpu.ALU.u_wallace._4379_ ;
 wire \u_cpu.ALU.u_wallace._4380_ ;
 wire \u_cpu.ALU.u_wallace._4381_ ;
 wire \u_cpu.ALU.u_wallace._4382_ ;
 wire \u_cpu.ALU.u_wallace._4383_ ;
 wire \u_cpu.ALU.u_wallace._4384_ ;
 wire \u_cpu.ALU.u_wallace._4385_ ;
 wire \u_cpu.ALU.u_wallace._4386_ ;
 wire \u_cpu.ALU.u_wallace._4387_ ;
 wire \u_cpu.ALU.u_wallace._4388_ ;
 wire \u_cpu.ALU.u_wallace._4389_ ;
 wire \u_cpu.ALU.u_wallace._4390_ ;
 wire \u_cpu.ALU.u_wallace._4391_ ;
 wire \u_cpu.ALU.u_wallace._4392_ ;
 wire \u_cpu.ALU.u_wallace._4393_ ;
 wire \u_cpu.ALU.u_wallace._4394_ ;
 wire \u_cpu.ALU.u_wallace._4395_ ;
 wire \u_cpu.ALU.u_wallace._4396_ ;
 wire \u_cpu.ALU.u_wallace._4397_ ;
 wire \u_cpu.ALU.u_wallace._4398_ ;
 wire \u_cpu.ALU.u_wallace._4399_ ;
 wire \u_cpu.ALU.u_wallace._4400_ ;
 wire \u_cpu.ALU.u_wallace._4401_ ;
 wire \u_cpu.ALU.u_wallace._4402_ ;
 wire \u_cpu.ALU.u_wallace._4403_ ;
 wire \u_cpu.ALU.u_wallace._4404_ ;
 wire \u_cpu.ALU.u_wallace._4405_ ;
 wire \u_cpu.ALU.u_wallace._4406_ ;
 wire \u_cpu.ALU.u_wallace._4407_ ;
 wire \u_cpu.ALU.u_wallace._4408_ ;
 wire \u_cpu.ALU.u_wallace._4409_ ;
 wire \u_cpu.ALU.u_wallace._4410_ ;
 wire \u_cpu.ALU.u_wallace._4411_ ;
 wire \u_cpu.ALU.u_wallace._4412_ ;
 wire \u_cpu.ALU.u_wallace._4413_ ;
 wire \u_cpu.ALU.u_wallace._4414_ ;
 wire \u_cpu.ALU.u_wallace._4415_ ;
 wire \u_cpu.ALU.u_wallace._4416_ ;
 wire \u_cpu.ALU.u_wallace._4417_ ;
 wire \u_cpu.ALU.u_wallace._4418_ ;
 wire \u_cpu.ALU.u_wallace._4419_ ;
 wire \u_cpu.ALU.u_wallace._4420_ ;
 wire \u_cpu.ALU.u_wallace._4421_ ;
 wire \u_cpu.ALU.u_wallace._4422_ ;
 wire \u_cpu.ALU.u_wallace._4423_ ;
 wire \u_cpu.ALU.u_wallace._4424_ ;
 wire \u_cpu.ALU.u_wallace._4425_ ;
 wire \u_cpu.ALU.u_wallace._4426_ ;
 wire \u_cpu.ALU.u_wallace._4427_ ;
 wire \u_cpu.ALU.u_wallace._4428_ ;
 wire \u_cpu.ALU.u_wallace._4429_ ;
 wire \u_cpu.ALU.u_wallace._4430_ ;
 wire \u_cpu.ALU.u_wallace._4431_ ;
 wire \u_cpu.ALU.u_wallace._4432_ ;
 wire \u_cpu.ALU.u_wallace._4433_ ;
 wire \u_cpu.ALU.u_wallace._4434_ ;
 wire \u_cpu.ALU.u_wallace._4435_ ;
 wire \u_cpu.ALU.u_wallace._4436_ ;
 wire \u_cpu.ALU.u_wallace._4437_ ;
 wire \u_cpu.ALU.u_wallace._4438_ ;
 wire \u_cpu.ALU.u_wallace._4439_ ;
 wire \u_cpu.ALU.u_wallace._4440_ ;
 wire \u_cpu.ALU.u_wallace._4441_ ;
 wire \u_cpu.ALU.u_wallace._4442_ ;
 wire \u_cpu.ALU.u_wallace._4443_ ;
 wire \u_cpu.ALU.u_wallace._4444_ ;
 wire \u_cpu.ALU.u_wallace._4445_ ;
 wire \u_cpu.ALU.u_wallace._4446_ ;
 wire \u_cpu.ALU.u_wallace._4447_ ;
 wire \u_cpu.ALU.u_wallace._4448_ ;
 wire \u_cpu.ALU.u_wallace._4449_ ;
 wire \u_cpu.ALU.u_wallace._4450_ ;
 wire \u_cpu.ALU.u_wallace._4451_ ;
 wire \u_cpu.ALU.u_wallace._4452_ ;
 wire \u_cpu.ALU.u_wallace._4453_ ;
 wire \u_cpu.ALU.u_wallace._4454_ ;
 wire \u_cpu.ALU.u_wallace._4455_ ;
 wire \u_cpu.ALU.u_wallace._4456_ ;
 wire \u_cpu.ALU.u_wallace._4457_ ;
 wire \u_cpu.ALU.u_wallace._4458_ ;
 wire \u_cpu.ALU.u_wallace._4459_ ;
 wire \u_cpu.ALU.u_wallace._4460_ ;
 wire \u_cpu.ALU.u_wallace._4461_ ;
 wire \u_cpu.ALU.u_wallace._4462_ ;
 wire \u_cpu.ALU.u_wallace._4463_ ;
 wire \u_cpu.ALU.u_wallace._4464_ ;
 wire \u_cpu.ALU.u_wallace._4465_ ;
 wire \u_cpu.ALU.u_wallace._4466_ ;
 wire \u_cpu.ALU.u_wallace._4467_ ;
 wire \u_cpu.ALU.u_wallace._4468_ ;
 wire \u_cpu.ALU.u_wallace._4469_ ;
 wire \u_cpu.ALU.u_wallace._4470_ ;
 wire \u_cpu.ALU.u_wallace._4471_ ;
 wire \u_cpu.ALU.u_wallace._4472_ ;
 wire \u_cpu.ALU.u_wallace._4473_ ;
 wire \u_cpu.ALU.u_wallace._4474_ ;
 wire \u_cpu.ALU.u_wallace._4475_ ;
 wire \u_cpu.ALU.u_wallace._4476_ ;
 wire \u_cpu.ALU.u_wallace._4477_ ;
 wire \u_cpu.ALU.u_wallace._4478_ ;
 wire \u_cpu.ALU.u_wallace._4479_ ;
 wire \u_cpu.ALU.u_wallace._4480_ ;
 wire \u_cpu.ALU.u_wallace._4481_ ;
 wire \u_cpu.ALU.u_wallace._4482_ ;
 wire \u_cpu.ALU.u_wallace._4483_ ;
 wire \u_cpu.ALU.u_wallace._4484_ ;
 wire \u_cpu.ALU.u_wallace._4485_ ;
 wire \u_cpu.ALU.u_wallace._4486_ ;
 wire \u_cpu.ALU.u_wallace._4487_ ;
 wire \u_cpu.ALU.u_wallace._4488_ ;
 wire \u_cpu.ALU.u_wallace._4489_ ;
 wire \u_cpu.ALU.u_wallace._4490_ ;
 wire \u_cpu.ALU.u_wallace._4491_ ;
 wire \u_cpu.ALU.u_wallace._4492_ ;
 wire \u_cpu.ALU.u_wallace._4493_ ;
 wire \u_cpu.ALU.u_wallace._4494_ ;
 wire \u_cpu.ALU.u_wallace._4495_ ;
 wire \u_cpu.ALU.u_wallace._4496_ ;
 wire \u_cpu.ALU.u_wallace._4497_ ;
 wire \u_cpu.ALU.u_wallace._4498_ ;
 wire \u_cpu.ALU.u_wallace._4499_ ;
 wire \u_cpu.ALU.u_wallace._4500_ ;
 wire \u_cpu.ALU.u_wallace._4501_ ;
 wire \u_cpu.ALU.u_wallace._4502_ ;
 wire \u_cpu.ALU.u_wallace._4503_ ;
 wire \u_cpu.ALU.u_wallace._4504_ ;
 wire \u_cpu.ALU.u_wallace._4505_ ;
 wire \u_cpu.ALU.u_wallace._4506_ ;
 wire \u_cpu.ALU.u_wallace._4507_ ;
 wire \u_cpu.ALU.u_wallace._4508_ ;
 wire \u_cpu.ALU.u_wallace._4509_ ;
 wire \u_cpu.ALU.u_wallace._4510_ ;
 wire \u_cpu.ALU.u_wallace._4511_ ;
 wire \u_cpu.ALU.u_wallace._4512_ ;
 wire \u_cpu.ALU.u_wallace._4513_ ;
 wire \u_cpu.ALU.u_wallace._4514_ ;
 wire \u_cpu.ALU.u_wallace._4515_ ;
 wire \u_cpu.ALU.u_wallace._4516_ ;
 wire \u_cpu.ALU.u_wallace._4517_ ;
 wire \u_cpu.ALU.u_wallace._4518_ ;
 wire \u_cpu.ALU.u_wallace._4519_ ;
 wire \u_cpu.ALU.u_wallace._4520_ ;
 wire \u_cpu.ALU.u_wallace._4521_ ;
 wire \u_cpu.ALU.u_wallace._4522_ ;
 wire \u_cpu.ALU.u_wallace._4523_ ;
 wire \u_cpu.ALU.u_wallace._4524_ ;
 wire \u_cpu.ALU.u_wallace._4525_ ;
 wire \u_cpu.ALU.u_wallace._4526_ ;
 wire \u_cpu.ALU.u_wallace._4527_ ;
 wire \u_cpu.ALU.u_wallace._4528_ ;
 wire \u_cpu.ALU.u_wallace._4529_ ;
 wire \u_cpu.ALU.u_wallace._4530_ ;
 wire \u_cpu.ALU.u_wallace._4531_ ;
 wire \u_cpu.ALU.u_wallace._4532_ ;
 wire \u_cpu.ALU.u_wallace._4533_ ;
 wire \u_cpu.ALU.u_wallace._4534_ ;
 wire \u_cpu.ALU.u_wallace._4535_ ;
 wire \u_cpu.ALU.u_wallace._4536_ ;
 wire \u_cpu.ALU.u_wallace._4537_ ;
 wire \u_cpu.ALU.u_wallace._4538_ ;
 wire \u_cpu.ALU.u_wallace._4539_ ;
 wire \u_cpu.ALU.u_wallace._4540_ ;
 wire \u_cpu.ALU.u_wallace._4541_ ;
 wire \u_cpu.ALU.u_wallace._4542_ ;
 wire \u_cpu.ALU.u_wallace._4543_ ;
 wire \u_cpu.ALU.u_wallace._4544_ ;
 wire \u_cpu.ALU.u_wallace._4545_ ;
 wire \u_cpu.ALU.u_wallace._4546_ ;
 wire \u_cpu.ALU.u_wallace._4547_ ;
 wire \u_cpu.ALU.u_wallace._4548_ ;
 wire \u_cpu.ALU.u_wallace._4549_ ;
 wire \u_cpu.ALU.u_wallace._4550_ ;
 wire \u_cpu.ALU.u_wallace._4551_ ;
 wire \u_cpu.ALU.u_wallace._4552_ ;
 wire \u_cpu.ALU.u_wallace._4553_ ;
 wire \u_cpu.ALU.u_wallace._4554_ ;
 wire \u_cpu.ALU.u_wallace._4555_ ;
 wire \u_cpu.ALU.u_wallace._4556_ ;
 wire \u_cpu.ALU.u_wallace._4557_ ;
 wire \u_cpu.ALU.u_wallace._4558_ ;
 wire \u_cpu.ALU.u_wallace._4559_ ;
 wire \u_cpu.ALU.u_wallace._4560_ ;
 wire \u_cpu.ALU.u_wallace._4561_ ;
 wire \u_cpu.ALU.u_wallace._4562_ ;
 wire \u_cpu.ALU.u_wallace._4563_ ;
 wire \u_cpu.ALU.u_wallace._4564_ ;
 wire \u_cpu.ALU.u_wallace._4565_ ;
 wire \u_cpu.ALU.u_wallace._4566_ ;
 wire \u_cpu.ALU.u_wallace._4567_ ;
 wire \u_cpu.ALU.u_wallace._4568_ ;
 wire \u_cpu.ALU.u_wallace._4569_ ;
 wire \u_cpu.ALU.u_wallace._4570_ ;
 wire \u_cpu.ALU.u_wallace._4571_ ;
 wire \u_cpu.ALU.u_wallace._4572_ ;
 wire \u_cpu.ALU.u_wallace._4573_ ;
 wire \u_cpu.ALU.u_wallace._4574_ ;
 wire \u_cpu.ALU.u_wallace._4575_ ;
 wire \u_cpu.ALU.u_wallace._4576_ ;
 wire \u_cpu.ALU.u_wallace._4577_ ;
 wire \u_cpu.ALU.u_wallace._4578_ ;
 wire \u_cpu.ALU.u_wallace._4579_ ;
 wire \u_cpu.ALU.u_wallace._4580_ ;
 wire \u_cpu.ALU.u_wallace._4581_ ;
 wire \u_cpu.ALU.u_wallace._4582_ ;
 wire \u_cpu.ALU.u_wallace._4583_ ;
 wire \u_cpu.ALU.u_wallace._4584_ ;
 wire \u_cpu.ALU.u_wallace._4585_ ;
 wire \u_cpu.ALU.u_wallace._4586_ ;
 wire \u_cpu.ALU.u_wallace._4587_ ;
 wire \u_cpu.ALU.u_wallace._4588_ ;
 wire \u_cpu.ALU.u_wallace._4589_ ;
 wire \u_cpu.ALU.u_wallace._4590_ ;
 wire \u_cpu.ALU.u_wallace._4591_ ;
 wire \u_cpu.ALU.u_wallace._4592_ ;
 wire \u_cpu.ALU.u_wallace._4593_ ;
 wire \u_cpu.ALU.u_wallace._4594_ ;
 wire \u_cpu.ALU.u_wallace._4595_ ;
 wire \u_cpu.ALU.u_wallace._4596_ ;
 wire \u_cpu.ALU.u_wallace._4597_ ;
 wire \u_cpu.ALU.u_wallace._4598_ ;
 wire \u_cpu.ALU.u_wallace._4599_ ;
 wire \u_cpu.ALU.u_wallace._4600_ ;
 wire \u_cpu.ALU.u_wallace._4601_ ;
 wire \u_cpu.ALU.u_wallace._4602_ ;
 wire \u_cpu.ALU.u_wallace._4603_ ;
 wire \u_cpu.ALU.u_wallace._4604_ ;
 wire \u_cpu.ALU.u_wallace._4605_ ;
 wire \u_cpu.ALU.u_wallace._4606_ ;
 wire \u_cpu.ALU.u_wallace._4607_ ;
 wire \u_cpu.ALU.u_wallace._4608_ ;
 wire \u_cpu.ALU.u_wallace._4609_ ;
 wire \u_cpu.ALU.u_wallace._4610_ ;
 wire \u_cpu.ALU.u_wallace._4611_ ;
 wire \u_cpu.ALU.u_wallace._4612_ ;
 wire \u_cpu.ALU.u_wallace._4613_ ;
 wire \u_cpu.ALU.u_wallace._4614_ ;
 wire \u_cpu.ALU.u_wallace._4615_ ;
 wire \u_cpu.ALU.u_wallace._4616_ ;
 wire \u_cpu.ALU.u_wallace._4617_ ;
 wire \u_cpu.ALU.u_wallace._4618_ ;
 wire \u_cpu.ALU.u_wallace._4619_ ;
 wire \u_cpu.ALU.u_wallace._4620_ ;
 wire \u_cpu.ALU.u_wallace._4621_ ;
 wire \u_cpu.ALU.u_wallace._4622_ ;
 wire \u_cpu.ALU.u_wallace._4623_ ;
 wire \u_cpu.ALU.u_wallace._4624_ ;
 wire \u_cpu.ALU.u_wallace._4625_ ;
 wire \u_cpu.ALU.u_wallace._4626_ ;
 wire \u_cpu.ALU.u_wallace._4627_ ;
 wire \u_cpu.ALU.u_wallace._4628_ ;
 wire \u_cpu.ALU.u_wallace._4629_ ;
 wire \u_cpu.ALU.u_wallace._4630_ ;
 wire \u_cpu.ALU.u_wallace._4631_ ;
 wire \u_cpu.ALU.u_wallace._4632_ ;
 wire \u_cpu.ALU.u_wallace._4633_ ;
 wire \u_cpu.ALU.u_wallace._4634_ ;
 wire \u_cpu.ALU.u_wallace._4635_ ;
 wire \u_cpu.ALU.u_wallace._4636_ ;
 wire \u_cpu.ALU.u_wallace._4637_ ;
 wire \u_cpu.ALU.u_wallace._4638_ ;
 wire \u_cpu.ALU.u_wallace._4639_ ;
 wire \u_cpu.ALU.u_wallace._4640_ ;
 wire \u_cpu.ALU.u_wallace._4641_ ;
 wire \u_cpu.ALU.u_wallace._4642_ ;
 wire \u_cpu.ALU.u_wallace._4643_ ;
 wire \u_cpu.ALU.u_wallace._4644_ ;
 wire \u_cpu.ALU.u_wallace._4645_ ;
 wire \u_cpu.ALU.u_wallace._4646_ ;
 wire \u_cpu.ALU.u_wallace._4647_ ;
 wire \u_cpu.ALU.u_wallace._4648_ ;
 wire \u_cpu.ALU.u_wallace._4649_ ;
 wire \u_cpu.ALU.u_wallace._4650_ ;
 wire \u_cpu.ALU.u_wallace._4651_ ;
 wire \u_cpu.ALU.u_wallace._4652_ ;
 wire \u_cpu.ALU.u_wallace._4653_ ;
 wire \u_cpu.ALU.u_wallace._4654_ ;
 wire \u_cpu.ALU.u_wallace._4655_ ;
 wire \u_cpu.ALU.u_wallace._4656_ ;
 wire \u_cpu.ALU.u_wallace._4657_ ;
 wire \u_cpu.ALU.u_wallace._4658_ ;
 wire \u_cpu.ALU.u_wallace._4659_ ;
 wire \u_cpu.ALU.u_wallace._4660_ ;
 wire \u_cpu.ALU.u_wallace._4661_ ;
 wire \u_cpu.ALU.u_wallace._4662_ ;
 wire \u_cpu.ALU.u_wallace._4663_ ;
 wire \u_cpu.ALU.u_wallace._4664_ ;
 wire \u_cpu.ALU.u_wallace._4665_ ;
 wire \u_cpu.ALU.u_wallace._4666_ ;
 wire \u_cpu.ALU.u_wallace._4667_ ;
 wire \u_cpu.ALU.u_wallace._4668_ ;
 wire \u_cpu.ALU.u_wallace._4669_ ;
 wire \u_cpu.ALU.u_wallace._4670_ ;
 wire \u_cpu.ALU.u_wallace._4671_ ;
 wire \u_cpu.ALU.u_wallace._4672_ ;
 wire \u_cpu.ALU.u_wallace._4673_ ;
 wire \u_cpu.ALU.u_wallace._4674_ ;
 wire \u_cpu.ALU.u_wallace._4675_ ;
 wire \u_cpu.ALU.u_wallace._4676_ ;
 wire \u_cpu.ALU.u_wallace._4677_ ;
 wire \u_cpu.ALU.u_wallace._4678_ ;
 wire \u_cpu.ALU.u_wallace._4679_ ;
 wire \u_cpu.ALU.u_wallace._4680_ ;
 wire \u_cpu.ALU.u_wallace._4681_ ;
 wire \u_cpu.ALU.u_wallace._4682_ ;
 wire \u_cpu.ALU.u_wallace._4683_ ;
 wire \u_cpu.ALU.u_wallace._4684_ ;
 wire \u_cpu.ALU.u_wallace._4685_ ;
 wire \u_cpu.ALU.u_wallace._4686_ ;
 wire \u_cpu.ALU.u_wallace._4687_ ;
 wire \u_cpu.ALU.u_wallace._4688_ ;
 wire \u_cpu.ALU.u_wallace._4689_ ;
 wire \u_cpu.ALU.u_wallace._4690_ ;
 wire \u_cpu.ALU.u_wallace._4691_ ;
 wire \u_cpu.ALU.u_wallace._4692_ ;
 wire \u_cpu.ALU.u_wallace._4693_ ;
 wire \u_cpu.ALU.u_wallace._4694_ ;
 wire \u_cpu.ALU.u_wallace._4695_ ;
 wire \u_cpu.ALU.u_wallace._4696_ ;
 wire \u_cpu.ALU.u_wallace._4697_ ;
 wire \u_cpu.ALU.u_wallace._4698_ ;
 wire \u_cpu.ALU.u_wallace._4699_ ;
 wire \u_cpu.ALU.u_wallace._4700_ ;
 wire \u_cpu.ALU.u_wallace._4701_ ;
 wire \u_cpu.ALU.u_wallace._4702_ ;
 wire \u_cpu.ALU.u_wallace._4703_ ;
 wire \u_cpu.ALU.u_wallace._4704_ ;
 wire \u_cpu.ALU.u_wallace._4705_ ;
 wire \u_cpu.ALU.u_wallace._4706_ ;
 wire \u_cpu.ALU.u_wallace._4707_ ;
 wire \u_cpu.ALU.u_wallace._4708_ ;
 wire \u_cpu.ALU.u_wallace._4709_ ;
 wire \u_cpu.ALU.u_wallace._4710_ ;
 wire \u_cpu.ALU.u_wallace._4711_ ;
 wire \u_cpu.ALU.u_wallace._4712_ ;
 wire \u_cpu.ALU.u_wallace._4713_ ;
 wire \u_cpu.ALU.u_wallace._4714_ ;
 wire \u_cpu.ALU.u_wallace._4715_ ;
 wire \u_cpu.ALU.u_wallace._4716_ ;
 wire \u_cpu.ALU.u_wallace._4717_ ;
 wire \u_cpu.ALU.u_wallace._4718_ ;
 wire \u_cpu.ALU.u_wallace._4719_ ;
 wire \u_cpu.ALU.u_wallace._4720_ ;
 wire \u_cpu.ALU.u_wallace._4721_ ;
 wire \u_cpu.ALU.u_wallace._4722_ ;
 wire \u_cpu.ALU.u_wallace._4723_ ;
 wire \u_cpu.ALU.u_wallace._4724_ ;
 wire \u_cpu.ALU.u_wallace._4725_ ;
 wire \u_cpu.ALU.u_wallace._4726_ ;
 wire \u_cpu.ALU.u_wallace._4727_ ;
 wire \u_cpu.ALU.u_wallace._4728_ ;
 wire \u_cpu.ALU.u_wallace._4729_ ;
 wire \u_cpu.ALU.u_wallace._4730_ ;
 wire \u_cpu.ALU.u_wallace._4731_ ;
 wire \u_cpu.ALU.u_wallace._4732_ ;
 wire \u_cpu.ALU.u_wallace._4733_ ;
 wire \u_cpu.ALU.u_wallace._4734_ ;
 wire \u_cpu.ALU.u_wallace._4735_ ;
 wire \u_cpu.ALU.u_wallace._4736_ ;
 wire \u_cpu.ALU.u_wallace._4737_ ;
 wire \u_cpu.ALU.u_wallace._4738_ ;
 wire \u_cpu.ALU.u_wallace._4739_ ;
 wire \u_cpu.ALU.u_wallace._4740_ ;
 wire \u_cpu.ALU.u_wallace._4741_ ;
 wire \u_cpu.ALU.u_wallace._4742_ ;
 wire \u_cpu.ALU.u_wallace._4743_ ;
 wire \u_cpu.ALU.u_wallace._4744_ ;
 wire \u_cpu.ALU.u_wallace._4745_ ;
 wire \u_cpu.ALU.u_wallace._4746_ ;
 wire \u_cpu.ALU.u_wallace._4747_ ;
 wire \u_cpu.ALU.u_wallace._4748_ ;
 wire \u_cpu.ALU.u_wallace._4749_ ;
 wire \u_cpu.ALU.u_wallace._4750_ ;
 wire \u_cpu.ALU.u_wallace._4751_ ;
 wire \u_cpu.ALU.u_wallace._4752_ ;
 wire \u_cpu.ALU.u_wallace._4753_ ;
 wire \u_cpu.ALU.u_wallace._4754_ ;
 wire \u_cpu.ALU.u_wallace._4755_ ;
 wire \u_cpu.ALU.u_wallace._4756_ ;
 wire \u_cpu.ALU.u_wallace._4757_ ;
 wire \u_cpu.ALU.u_wallace._4758_ ;
 wire \u_cpu.ALU.u_wallace._4759_ ;
 wire \u_cpu.ALU.u_wallace._4760_ ;
 wire \u_cpu.ALU.u_wallace._4761_ ;
 wire \u_cpu.ALU.u_wallace._4762_ ;
 wire \u_cpu.ALU.u_wallace._4763_ ;
 wire \u_cpu.ALU.u_wallace._4764_ ;
 wire \u_cpu.ALU.u_wallace._4765_ ;
 wire \u_cpu.ALU.u_wallace._4766_ ;
 wire \u_cpu.ALU.u_wallace._4767_ ;
 wire \u_cpu.ALU.u_wallace._4768_ ;
 wire \u_cpu.ALU.u_wallace._4769_ ;
 wire \u_cpu.ALU.u_wallace._4770_ ;
 wire \u_cpu.ALU.u_wallace._4771_ ;
 wire \u_cpu.ALU.u_wallace._4772_ ;
 wire \u_cpu.ALU.u_wallace._4773_ ;
 wire \u_cpu.ALU.u_wallace._4774_ ;
 wire \u_cpu.ALU.u_wallace._4775_ ;
 wire \u_cpu.ALU.u_wallace._4776_ ;
 wire \u_cpu.ALU.u_wallace._4777_ ;
 wire \u_cpu.ALU.u_wallace._4778_ ;
 wire \u_cpu.ALU.u_wallace._4779_ ;
 wire \u_cpu.ALU.u_wallace._4780_ ;
 wire \u_cpu.ALU.u_wallace._4781_ ;
 wire \u_cpu.ALU.u_wallace._4782_ ;
 wire \u_cpu.ALU.u_wallace._4783_ ;
 wire \u_cpu.ALU.u_wallace._4784_ ;
 wire \u_cpu.ALU.u_wallace._4785_ ;
 wire \u_cpu.ALU.u_wallace._4786_ ;
 wire \u_cpu.ALU.u_wallace._4787_ ;
 wire \u_cpu.ALU.u_wallace._4788_ ;
 wire \u_cpu.ALU.u_wallace._4789_ ;
 wire \u_cpu.ALU.u_wallace._4790_ ;
 wire \u_cpu.ALU.u_wallace._4791_ ;
 wire \u_cpu.ALU.u_wallace._4792_ ;
 wire \u_cpu.ALU.u_wallace._4793_ ;
 wire \u_cpu.ALU.u_wallace._4794_ ;
 wire \u_cpu.ALU.u_wallace._4795_ ;
 wire \u_cpu.ALU.u_wallace._4796_ ;
 wire \u_cpu.ALU.u_wallace._4797_ ;
 wire \u_cpu.ALU.u_wallace._4798_ ;
 wire \u_cpu.ALU.u_wallace._4799_ ;
 wire \u_cpu.ALU.u_wallace._4800_ ;
 wire \u_cpu.ALU.u_wallace._4801_ ;
 wire \u_cpu.ALU.u_wallace._4802_ ;
 wire \u_cpu.ALU.u_wallace._4803_ ;
 wire \u_cpu.ALU.u_wallace._4804_ ;
 wire \u_cpu.ALU.u_wallace._4805_ ;
 wire \u_cpu.ALU.u_wallace._4806_ ;
 wire \u_cpu.ALU.u_wallace._4807_ ;
 wire \u_cpu.ALU.u_wallace._4808_ ;
 wire \u_cpu.ALU.u_wallace._4809_ ;
 wire \u_cpu.ALU.u_wallace._4810_ ;
 wire \u_cpu.ALU.u_wallace._4811_ ;
 wire \u_cpu.ALU.u_wallace._4812_ ;
 wire \u_cpu.ALU.u_wallace._4813_ ;
 wire \u_cpu.ALU.u_wallace._4814_ ;
 wire \u_cpu.ALU.u_wallace._4815_ ;
 wire \u_cpu.ALU.u_wallace._4816_ ;
 wire \u_cpu.ALU.u_wallace._4817_ ;
 wire \u_cpu.ALU.u_wallace._4818_ ;
 wire \u_cpu.ALU.u_wallace._4819_ ;
 wire \u_cpu.ALU.u_wallace._4820_ ;
 wire \u_cpu.ALU.u_wallace._4821_ ;
 wire \u_cpu.ALU.u_wallace._4822_ ;
 wire \u_cpu.ALU.u_wallace._4823_ ;
 wire \u_cpu.ALU.u_wallace._4824_ ;
 wire \u_cpu.ALU.u_wallace._4825_ ;
 wire \u_cpu.ALU.u_wallace._4826_ ;
 wire \u_cpu.ALU.u_wallace._4827_ ;
 wire \u_cpu.ALU.u_wallace._4828_ ;
 wire \u_cpu.ALU.u_wallace._4829_ ;
 wire \u_cpu.ALU.u_wallace._4830_ ;
 wire \u_cpu.ALU.u_wallace._4831_ ;
 wire \u_cpu.ALU.u_wallace._4832_ ;
 wire \u_cpu.ALU.u_wallace._4833_ ;
 wire \u_cpu.ALU.u_wallace._4834_ ;
 wire \u_cpu.ALU.u_wallace._4835_ ;
 wire \u_cpu.ALU.u_wallace._4836_ ;
 wire \u_cpu.ALU.u_wallace._4837_ ;
 wire \u_cpu.ALU.u_wallace._4838_ ;
 wire \u_cpu.ALU.u_wallace._4839_ ;
 wire \u_cpu.ALU.u_wallace._4840_ ;
 wire \u_cpu.ALU.u_wallace._4841_ ;
 wire \u_cpu.ALU.u_wallace._4842_ ;
 wire \u_cpu.ALU.u_wallace._4843_ ;
 wire \u_cpu.ALU.u_wallace._4844_ ;
 wire \u_cpu.ALU.u_wallace._4845_ ;
 wire \u_cpu.ALU.u_wallace._4846_ ;
 wire \u_cpu.ALU.u_wallace._4847_ ;
 wire \u_cpu.ALU.u_wallace._4848_ ;
 wire \u_cpu.ALU.u_wallace._4849_ ;
 wire \u_cpu.ALU.u_wallace._4850_ ;
 wire \u_cpu.ALU.u_wallace._4851_ ;
 wire \u_cpu.ALU.u_wallace._4852_ ;
 wire \u_cpu.ALU.u_wallace._4853_ ;
 wire \u_cpu.ALU.u_wallace._4854_ ;
 wire \u_cpu.ALU.u_wallace._4855_ ;
 wire \u_cpu.ALU.u_wallace._4856_ ;
 wire \u_cpu.ALU.u_wallace._4857_ ;
 wire \u_cpu.ALU.u_wallace._4858_ ;
 wire \u_cpu.ALU.u_wallace._4859_ ;
 wire \u_cpu.ALU.u_wallace._4860_ ;
 wire \u_cpu.ALU.u_wallace._4861_ ;
 wire \u_cpu.ALU.u_wallace._4862_ ;
 wire \u_cpu.ALU.u_wallace._4863_ ;
 wire \u_cpu.ALU.u_wallace._4864_ ;
 wire \u_cpu.ALU.u_wallace._4865_ ;
 wire \u_cpu.ALU.u_wallace._4866_ ;
 wire \u_cpu.ALU.u_wallace._4867_ ;
 wire \u_cpu.ALU.u_wallace._4868_ ;
 wire \u_cpu.ALU.u_wallace._4869_ ;
 wire \u_cpu.ALU.u_wallace._4870_ ;
 wire \u_cpu.ALU.u_wallace._4871_ ;
 wire \u_cpu.ALU.u_wallace._4872_ ;
 wire \u_cpu.ALU.u_wallace._4873_ ;
 wire \u_cpu.ALU.u_wallace._4874_ ;
 wire \u_cpu.ALU.u_wallace._4875_ ;
 wire \u_cpu.ALU.u_wallace._4876_ ;
 wire \u_cpu.ALU.u_wallace._4877_ ;
 wire \u_cpu.ALU.u_wallace._4878_ ;
 wire \u_cpu.ALU.u_wallace._4879_ ;
 wire \u_cpu.ALU.u_wallace._4880_ ;
 wire \u_cpu.ALU.u_wallace._4881_ ;
 wire \u_cpu.ALU.u_wallace._4882_ ;
 wire \u_cpu.ALU.u_wallace._4883_ ;
 wire \u_cpu.ALU.u_wallace._4884_ ;
 wire \u_cpu.ALU.u_wallace._4885_ ;
 wire \u_cpu.ALU.u_wallace._4886_ ;
 wire \u_cpu.ALU.u_wallace._4887_ ;
 wire \u_cpu.ALU.u_wallace._4888_ ;
 wire \u_cpu.ALU.u_wallace._4889_ ;
 wire \u_cpu.ALU.u_wallace._4890_ ;
 wire \u_cpu.ALU.u_wallace._4891_ ;
 wire \u_cpu.ALU.u_wallace._4892_ ;
 wire \u_cpu.ALU.u_wallace._4893_ ;
 wire \u_cpu.ALU.u_wallace._4894_ ;
 wire \u_cpu.ALU.u_wallace._4895_ ;
 wire \u_cpu.ALU.u_wallace._4896_ ;
 wire \u_cpu.ALU.u_wallace._4897_ ;
 wire \u_cpu.ALU.u_wallace._4898_ ;
 wire \u_cpu.ALU.u_wallace._4899_ ;
 wire \u_cpu.ALU.u_wallace._4900_ ;
 wire \u_cpu.ALU.u_wallace._4901_ ;
 wire \u_cpu.ALU.u_wallace._4902_ ;
 wire \u_cpu.ALU.u_wallace._4903_ ;
 wire \u_cpu.ALU.u_wallace._4904_ ;
 wire \u_cpu.ALU.u_wallace._4905_ ;
 wire \u_cpu.ALU.u_wallace._4906_ ;
 wire \u_cpu.ALU.u_wallace._4907_ ;
 wire \u_cpu.ALU.u_wallace._4908_ ;
 wire \u_cpu.ALU.u_wallace._4909_ ;
 wire \u_cpu.ALU.u_wallace._4910_ ;
 wire \u_cpu.ALU.u_wallace._4911_ ;
 wire \u_cpu.ALU.u_wallace._4912_ ;
 wire \u_cpu.ALU.u_wallace._4913_ ;
 wire \u_cpu.ALU.u_wallace._4914_ ;
 wire \u_cpu.ALU.u_wallace._4915_ ;
 wire \u_cpu.ALU.u_wallace._4916_ ;
 wire \u_cpu.ALU.u_wallace._4917_ ;
 wire \u_cpu.ALU.u_wallace._4918_ ;
 wire \u_cpu.ALU.u_wallace._4919_ ;
 wire \u_cpu.ALU.u_wallace._4920_ ;
 wire \u_cpu.ALU.u_wallace._4921_ ;
 wire \u_cpu.ALU.u_wallace._4922_ ;
 wire \u_cpu.ALU.u_wallace._4923_ ;
 wire \u_cpu.ALU.u_wallace._4924_ ;
 wire \u_cpu.ALU.u_wallace._4925_ ;
 wire \u_cpu.ALU.u_wallace._4926_ ;
 wire \u_cpu.ALU.u_wallace._4927_ ;
 wire \u_cpu.ALU.u_wallace._4928_ ;
 wire \u_cpu.ALU.u_wallace._4929_ ;
 wire \u_cpu.ALU.u_wallace._4930_ ;
 wire \u_cpu.ALU.u_wallace._4931_ ;
 wire \u_cpu.ALU.u_wallace._4932_ ;
 wire \u_cpu.ALU.u_wallace._4933_ ;
 wire \u_cpu.ALU.u_wallace._4934_ ;
 wire \u_cpu.ALUResult_W_Reg[0] ;
 wire \u_cpu.ALUResult_W_Reg[10] ;
 wire \u_cpu.ALUResult_W_Reg[11] ;
 wire \u_cpu.ALUResult_W_Reg[12] ;
 wire \u_cpu.ALUResult_W_Reg[13] ;
 wire \u_cpu.ALUResult_W_Reg[14] ;
 wire \u_cpu.ALUResult_W_Reg[15] ;
 wire \u_cpu.ALUResult_W_Reg[16] ;
 wire \u_cpu.ALUResult_W_Reg[17] ;
 wire \u_cpu.ALUResult_W_Reg[18] ;
 wire \u_cpu.ALUResult_W_Reg[19] ;
 wire \u_cpu.ALUResult_W_Reg[20] ;
 wire \u_cpu.ALUResult_W_Reg[21] ;
 wire \u_cpu.ALUResult_W_Reg[22] ;
 wire \u_cpu.ALUResult_W_Reg[23] ;
 wire \u_cpu.ALUResult_W_Reg[24] ;
 wire \u_cpu.ALUResult_W_Reg[25] ;
 wire \u_cpu.ALUResult_W_Reg[26] ;
 wire \u_cpu.ALUResult_W_Reg[27] ;
 wire \u_cpu.ALUResult_W_Reg[28] ;
 wire \u_cpu.ALUResult_W_Reg[29] ;
 wire \u_cpu.ALUResult_W_Reg[30] ;
 wire \u_cpu.ALUResult_W_Reg[31] ;
 wire \u_cpu.IMEM._0000_ ;
 wire \u_cpu.IMEM._0001_ ;
 wire \u_cpu.IMEM._0002_ ;
 wire \u_cpu.IMEM._0003_ ;
 wire \u_cpu.IMEM._0004_ ;
 wire \u_cpu.IMEM._0005_ ;
 wire \u_cpu.IMEM._0006_ ;
 wire \u_cpu.IMEM._0007_ ;
 wire \u_cpu.IMEM._0008_ ;
 wire \u_cpu.IMEM._0009_ ;
 wire \u_cpu.IMEM._0010_ ;
 wire \u_cpu.IMEM._0011_ ;
 wire \u_cpu.IMEM._0012_ ;
 wire \u_cpu.IMEM._0013_ ;
 wire \u_cpu.IMEM._0014_ ;
 wire \u_cpu.IMEM._0015_ ;
 wire \u_cpu.IMEM._0016_ ;
 wire \u_cpu.IMEM._0017_ ;
 wire \u_cpu.IMEM._0018_ ;
 wire \u_cpu.IMEM._0019_ ;
 wire \u_cpu.IMEM._0020_ ;
 wire \u_cpu.IMEM._0021_ ;
 wire \u_cpu.IMEM._0022_ ;
 wire \u_cpu.IMEM._0023_ ;
 wire \u_cpu.IMEM._0024_ ;
 wire \u_cpu.IMEM._0025_ ;
 wire \u_cpu.IMEM._0026_ ;
 wire \u_cpu.IMEM._0027_ ;
 wire \u_cpu.IMEM._0028_ ;
 wire \u_cpu.IMEM._0029_ ;
 wire \u_cpu.IMEM._0030_ ;
 wire \u_cpu.IMEM._0031_ ;
 wire \u_cpu.IMEM._0032_ ;
 wire \u_cpu.IMEM._0033_ ;
 wire \u_cpu.IMEM._0034_ ;
 wire \u_cpu.IMEM._0035_ ;
 wire \u_cpu.IMEM._0036_ ;
 wire \u_cpu.IMEM._0037_ ;
 wire \u_cpu.IMEM._0038_ ;
 wire \u_cpu.IMEM._0039_ ;
 wire \u_cpu.IMEM._0040_ ;
 wire \u_cpu.IMEM._0041_ ;
 wire \u_cpu.IMEM._0042_ ;
 wire \u_cpu.IMEM._0043_ ;
 wire \u_cpu.IMEM._0044_ ;
 wire \u_cpu.IMEM._0045_ ;
 wire \u_cpu.IMEM._0046_ ;
 wire \u_cpu.IMEM._0047_ ;
 wire \u_cpu.IMEM._0048_ ;
 wire \u_cpu.IMEM._0049_ ;
 wire \u_cpu.IMEM._0050_ ;
 wire \u_cpu.IMEM._0051_ ;
 wire \u_cpu.IMEM._0052_ ;
 wire \u_cpu.IMEM._0053_ ;
 wire \u_cpu.IMEM._0054_ ;
 wire \u_cpu.IMEM._0055_ ;
 wire \u_cpu.IMEM._0056_ ;
 wire \u_cpu.IMEM._0057_ ;
 wire \u_cpu.IMEM._0058_ ;
 wire \u_cpu.IMEM._0059_ ;
 wire \u_cpu.IMEM._0060_ ;
 wire \u_cpu.IMEM._0061_ ;
 wire \u_cpu.IMEM._0062_ ;
 wire \u_cpu.IMEM._0063_ ;
 wire \u_cpu.IMEM._0064_ ;
 wire \u_cpu.IMEM._0065_ ;
 wire \u_cpu.IMEM._0066_ ;
 wire \u_cpu.IMEM._0067_ ;
 wire \u_cpu.IMEM._0068_ ;
 wire \u_cpu.IMEM._0069_ ;
 wire \u_cpu.IMEM._0070_ ;
 wire \u_cpu.IMEM._0071_ ;
 wire \u_cpu.IMEM._0072_ ;
 wire \u_cpu.IMEM._0073_ ;
 wire \u_cpu.IMEM._0074_ ;
 wire \u_cpu.IMEM._0075_ ;
 wire \u_cpu.IMEM._0076_ ;
 wire \u_cpu.IMEM._0077_ ;
 wire \u_cpu.IMEM._0078_ ;
 wire \u_cpu.IMEM._0079_ ;
 wire \u_cpu.IMEM._0080_ ;
 wire \u_cpu.IMEM._0081_ ;
 wire \u_cpu.IMEM._0082_ ;
 wire \u_cpu.IMEM._0083_ ;
 wire \u_cpu.IMEM._0084_ ;
 wire \u_cpu.IMEM._0085_ ;
 wire \u_cpu.IMEM._0086_ ;
 wire \u_cpu.IMEM._0087_ ;
 wire \u_cpu.IMEM._0088_ ;
 wire \u_cpu.IMEM._0089_ ;
 wire \u_cpu.IMEM._0090_ ;
 wire \u_cpu.IMEM._0091_ ;
 wire \u_cpu.IMEM._0092_ ;
 wire \u_cpu.IMEM._0093_ ;
 wire \u_cpu.IMEM._0094_ ;
 wire \u_cpu.IMEM._0095_ ;
 wire \u_cpu.IMEM._0096_ ;
 wire \u_cpu.IMEM._0097_ ;
 wire \u_cpu.IMEM._0098_ ;
 wire \u_cpu.IMEM._0099_ ;
 wire \u_cpu.IMEM._0100_ ;
 wire \u_cpu.IMEM._0101_ ;
 wire \u_cpu.IMEM._0102_ ;
 wire \u_cpu.IMEM._0103_ ;
 wire \u_cpu.IMEM._0104_ ;
 wire \u_cpu.IMEM._0105_ ;
 wire \u_cpu.IMEM._0106_ ;
 wire \u_cpu.IMEM._0107_ ;
 wire \u_cpu.IMEM._0108_ ;
 wire \u_cpu.IMEM._0109_ ;
 wire \u_cpu.IMEM._0110_ ;
 wire \u_cpu.IMEM._0111_ ;
 wire \u_cpu.IMEM._0112_ ;
 wire \u_cpu.IMEM._0113_ ;
 wire \u_cpu.IMEM._0114_ ;
 wire \u_cpu.IMEM._0115_ ;
 wire \u_cpu.IMEM._0116_ ;
 wire \u_cpu.IMEM._0117_ ;
 wire \u_cpu.IMEM._0118_ ;
 wire \u_cpu.IMEM._0119_ ;
 wire \u_cpu.IMEM._0120_ ;
 wire \u_cpu.IMEM._0121_ ;
 wire \u_cpu.IMEM._0122_ ;
 wire \u_cpu.IMEM._0123_ ;
 wire \u_cpu.IMEM._0124_ ;
 wire \u_cpu.IMEM._0125_ ;
 wire \u_cpu.IMEM._0126_ ;
 wire \u_cpu.IMEM._0127_ ;
 wire \u_cpu.IMEM._0128_ ;
 wire \u_cpu.IMEM._0129_ ;
 wire \u_cpu.IMEM._0130_ ;
 wire \u_cpu.IMEM._0131_ ;
 wire \u_cpu.IMEM._0132_ ;
 wire \u_cpu.IMEM._0133_ ;
 wire \u_cpu.IMEM._0134_ ;
 wire \u_cpu.IMEM._0135_ ;
 wire \u_cpu.IMEM._0136_ ;
 wire \u_cpu.IMEM._0137_ ;
 wire \u_cpu.IMEM._0138_ ;
 wire \u_cpu.IMEM._0139_ ;
 wire \u_cpu.IMEM._0140_ ;
 wire \u_cpu.IMEM._0141_ ;
 wire \u_cpu.IMEM._0142_ ;
 wire \u_cpu.IMEM._0143_ ;
 wire \u_cpu.IMEM._0144_ ;
 wire \u_cpu.IMEM._0145_ ;
 wire \u_cpu.IMEM._0146_ ;
 wire \u_cpu.IMEM._0147_ ;
 wire \u_cpu.IMEM._0148_ ;
 wire \u_cpu.IMEM._0149_ ;
 wire \u_cpu.IMEM._0150_ ;
 wire \u_cpu.IMEM._0151_ ;
 wire \u_cpu.IMEM._0152_ ;
 wire \u_cpu.IMEM._0153_ ;
 wire \u_cpu.IMEM._0154_ ;
 wire \u_cpu.IMEM._0155_ ;
 wire \u_cpu.IMEM._0156_ ;
 wire \u_cpu.IMEM._0157_ ;
 wire \u_cpu.IMEM._0158_ ;
 wire \u_cpu.IMEM._0159_ ;
 wire \u_cpu.IMEM._0160_ ;
 wire \u_cpu.IMEM._0161_ ;
 wire \u_cpu.IMEM._0162_ ;
 wire \u_cpu.IMEM._0163_ ;
 wire \u_cpu.IMEM._0164_ ;
 wire \u_cpu.IMEM._0165_ ;
 wire \u_cpu.IMEM._0166_ ;
 wire \u_cpu.IMEM._0167_ ;
 wire \u_cpu.IMEM._0168_ ;
 wire \u_cpu.IMEM._0169_ ;
 wire \u_cpu.IMEM._0170_ ;
 wire \u_cpu.IMEM._0171_ ;
 wire \u_cpu.IMEM._0172_ ;
 wire \u_cpu.IMEM._0173_ ;
 wire \u_cpu.IMEM._0174_ ;
 wire \u_cpu.IMEM._0175_ ;
 wire \u_cpu.IMEM._0176_ ;
 wire \u_cpu.IMEM._0177_ ;
 wire \u_cpu.IMEM._0178_ ;
 wire \u_cpu.IMEM._0179_ ;
 wire \u_cpu.IMEM._0180_ ;
 wire \u_cpu.IMEM._0181_ ;
 wire \u_cpu.IMEM._0182_ ;
 wire \u_cpu.IMEM._0183_ ;
 wire \u_cpu.IMEM._0184_ ;
 wire \u_cpu.IMEM._0185_ ;
 wire \u_cpu.IMEM._0186_ ;
 wire \u_cpu.IMEM._0187_ ;
 wire \u_cpu.IMEM._0188_ ;
 wire \u_cpu.IMEM._0189_ ;
 wire \u_cpu.IMEM._0190_ ;
 wire \u_cpu.IMEM._0191_ ;
 wire \u_cpu.IMEM._0192_ ;
 wire \u_cpu.IMEM._0193_ ;
 wire \u_cpu.IMEM._0194_ ;
 wire \u_cpu.IMEM._0195_ ;
 wire \u_cpu.IMEM._0196_ ;
 wire \u_cpu.IMEM._0197_ ;
 wire \u_cpu.IMEM._0198_ ;
 wire \u_cpu.IMEM._0199_ ;
 wire \u_cpu.IMEM._0200_ ;
 wire \u_cpu.IMEM._0201_ ;
 wire \u_cpu.IMEM._0202_ ;
 wire \u_cpu.IMEM._0203_ ;
 wire \u_cpu.IMEM._0204_ ;
 wire \u_cpu.IMEM._0205_ ;
 wire \u_cpu.IMEM._0206_ ;
 wire \u_cpu.IMEM._0207_ ;
 wire \u_cpu.IMEM._0208_ ;
 wire \u_cpu.IMEM._0209_ ;
 wire \u_cpu.IMEM._0210_ ;
 wire \u_cpu.IMEM._0211_ ;
 wire \u_cpu.IMEM._0212_ ;
 wire \u_cpu.IMEM._0213_ ;
 wire \u_cpu.IMEM._0214_ ;
 wire \u_cpu.IMEM._0215_ ;
 wire \u_cpu.IMEM._0216_ ;
 wire \u_cpu.IMEM._0217_ ;
 wire \u_cpu.IMEM._0218_ ;
 wire \u_cpu.IMEM._0219_ ;
 wire \u_cpu.IMEM._0220_ ;
 wire \u_cpu.IMEM._0221_ ;
 wire \u_cpu.IMEM._0222_ ;
 wire \u_cpu.IMEM._0223_ ;
 wire \u_cpu.IMEM._0224_ ;
 wire \u_cpu.IMEM._0225_ ;
 wire \u_cpu.IMEM._0226_ ;
 wire \u_cpu.IMEM._0227_ ;
 wire \u_cpu.IMEM._0228_ ;
 wire \u_cpu.IMEM._0229_ ;
 wire \u_cpu.IMEM._0230_ ;
 wire \u_cpu.IMEM._0231_ ;
 wire \u_cpu.IMEM._0232_ ;
 wire \u_cpu.IMEM._0233_ ;
 wire \u_cpu.IMEM._0234_ ;
 wire \u_cpu.IMEM._0235_ ;
 wire \u_cpu.IMEM._0236_ ;
 wire \u_cpu.IMEM._0237_ ;
 wire \u_cpu.IMEM._0238_ ;
 wire \u_cpu.IMEM._0239_ ;
 wire \u_cpu.IMEM._0240_ ;
 wire \u_cpu.IMEM._0241_ ;
 wire \u_cpu.IMEM._0242_ ;
 wire \u_cpu.IMEM._0243_ ;
 wire \u_cpu.IMEM._0244_ ;
 wire \u_cpu.IMEM._0245_ ;
 wire \u_cpu.IMEM._0246_ ;
 wire \u_cpu.IMEM._0247_ ;
 wire \u_cpu.IMEM._0248_ ;
 wire \u_cpu.IMEM._0249_ ;
 wire \u_cpu.IMEM._0250_ ;
 wire \u_cpu.IMEM._0251_ ;
 wire \u_cpu.IMEM._0252_ ;
 wire \u_cpu.IMEM._0253_ ;
 wire \u_cpu.IMEM._0254_ ;
 wire \u_cpu.IMEM._0255_ ;
 wire \u_cpu.IMEM._0256_ ;
 wire \u_cpu.IMEM._0257_ ;
 wire \u_cpu.IMEM._0258_ ;
 wire \u_cpu.IMEM._0259_ ;
 wire \u_cpu.IMEM._0260_ ;
 wire \u_cpu.IMEM._0261_ ;
 wire \u_cpu.IMEM._0262_ ;
 wire \u_cpu.IMEM._0263_ ;
 wire \u_cpu.IMEM._0264_ ;
 wire \u_cpu.IMEM._0265_ ;
 wire \u_cpu.IMEM._0266_ ;
 wire \u_cpu.IMEM._0267_ ;
 wire \u_cpu.IMEM._0268_ ;
 wire \u_cpu.IMEM._0269_ ;
 wire \u_cpu.IMEM._0270_ ;
 wire \u_cpu.IMEM._0271_ ;
 wire \u_cpu.IMEM._0272_ ;
 wire \u_cpu.IMEM._0273_ ;
 wire \u_cpu.IMEM._0274_ ;
 wire \u_cpu.IMEM._0275_ ;
 wire \u_cpu.IMEM._0276_ ;
 wire \u_cpu.IMEM._0277_ ;
 wire \u_cpu.IMEM._0278_ ;
 wire \u_cpu.IMEM._0279_ ;
 wire \u_cpu.IMEM._0280_ ;
 wire \u_cpu.IMEM._0281_ ;
 wire \u_cpu.IMEM._0282_ ;
 wire \u_cpu.IMEM._0283_ ;
 wire \u_cpu.IMEM._0284_ ;
 wire \u_cpu.IMEM._0285_ ;
 wire \u_cpu.IMEM._0286_ ;
 wire \u_cpu.IMEM._0287_ ;
 wire \u_cpu.IMEM._0288_ ;
 wire \u_cpu.IMEM._0289_ ;
 wire \u_cpu.IMEM._0290_ ;
 wire \u_cpu.IMEM._0291_ ;
 wire \u_cpu.IMEM._0292_ ;
 wire \u_cpu.IMEM._0293_ ;
 wire \u_cpu.IMEM._0294_ ;
 wire \u_cpu.IMEM._0295_ ;
 wire \u_cpu.IMEM._0296_ ;
 wire \u_cpu.IMEM._0297_ ;
 wire \u_cpu.IMEM._0298_ ;
 wire \u_cpu.IMEM._0299_ ;
 wire \u_cpu.IMEM._0300_ ;
 wire \u_cpu.IMEM._0301_ ;
 wire \u_cpu.IMEM._0302_ ;
 wire \u_cpu.IMEM._0303_ ;
 wire \u_cpu.IMEM._0304_ ;
 wire \u_cpu.IMEM._0305_ ;
 wire \u_cpu.IMEM._0306_ ;
 wire \u_cpu.IMEM._0307_ ;
 wire \u_cpu.IMEM._0308_ ;
 wire \u_cpu.IMEM._0309_ ;
 wire \u_cpu.IMEM._0310_ ;
 wire \u_cpu.IMEM._0311_ ;
 wire \u_cpu.IMEM._0312_ ;
 wire \u_cpu.IMEM._0313_ ;
 wire \u_cpu.IMEM._0314_ ;
 wire \u_cpu.IMEM._0315_ ;
 wire \u_cpu.IMEM._0316_ ;
 wire \u_cpu.IMEM._0317_ ;
 wire \u_cpu.IMEM._0318_ ;
 wire \u_cpu.IMEM._0319_ ;
 wire \u_cpu.IMEM._0320_ ;
 wire \u_cpu.IMEM._0321_ ;
 wire \u_cpu.IMEM._0322_ ;
 wire \u_cpu.IMEM._0323_ ;
 wire \u_cpu.IMEM._0324_ ;
 wire \u_cpu.IMEM._0325_ ;
 wire \u_cpu.IMEM._0326_ ;
 wire \u_cpu.IMEM._0327_ ;
 wire \u_cpu.IMEM._0328_ ;
 wire \u_cpu.IMEM._0329_ ;
 wire \u_cpu.IMEM._0330_ ;
 wire \u_cpu.IMEM._0331_ ;
 wire \u_cpu.IMEM._0332_ ;
 wire \u_cpu.IMEM._0333_ ;
 wire \u_cpu.IMEM._0334_ ;
 wire \u_cpu.IMEM._0335_ ;
 wire \u_cpu.IMEM._0336_ ;
 wire \u_cpu.IMEM._0337_ ;
 wire \u_cpu.IMEM._0338_ ;
 wire \u_cpu.IMEM._0339_ ;
 wire \u_cpu.IMEM._0340_ ;
 wire \u_cpu.IMEM._0341_ ;
 wire \u_cpu.IMEM._0342_ ;
 wire \u_cpu.IMEM._0343_ ;
 wire \u_cpu.IMEM._0344_ ;
 wire \u_cpu.IMEM._0345_ ;
 wire \u_cpu.IMEM._0346_ ;
 wire \u_cpu.IMEM._0347_ ;
 wire \u_cpu.IMEM._0348_ ;
 wire \u_cpu.IMEM._0349_ ;
 wire \u_cpu.IMEM._0350_ ;
 wire \u_cpu.IMEM._0351_ ;
 wire \u_cpu.IMEM._0352_ ;
 wire \u_cpu.IMEM._0353_ ;
 wire \u_cpu.IMEM._0354_ ;
 wire \u_cpu.IMEM._0355_ ;
 wire \u_cpu.IMEM._0356_ ;
 wire \u_cpu.IMEM._0357_ ;
 wire \u_cpu.IMEM._0358_ ;
 wire \u_cpu.IMEM._0359_ ;
 wire \u_cpu.IMEM._0360_ ;
 wire \u_cpu.IMEM._0361_ ;
 wire \u_cpu.IMEM._0362_ ;
 wire \u_cpu.IMEM._0363_ ;
 wire \u_cpu.IMEM._0364_ ;
 wire \u_cpu.IMEM._0365_ ;
 wire \u_cpu.IMEM._0366_ ;
 wire \u_cpu.IMEM._0367_ ;
 wire \u_cpu.IMEM._0368_ ;
 wire \u_cpu.IMEM._0369_ ;
 wire \u_cpu.IMEM._0370_ ;
 wire \u_cpu.IMEM._0371_ ;
 wire \u_cpu.IMEM._0372_ ;
 wire \u_cpu.IMEM._0373_ ;
 wire \u_cpu.IMEM._0374_ ;
 wire \u_cpu.IMEM._0375_ ;
 wire \u_cpu.IMEM._0376_ ;
 wire \u_cpu.IMEM._0377_ ;
 wire \u_cpu.IMEM._0378_ ;
 wire \u_cpu.IMEM._0379_ ;
 wire \u_cpu.IMEM._0380_ ;
 wire \u_cpu.IMEM._0381_ ;
 wire \u_cpu.IMEM._0382_ ;
 wire \u_cpu.IMEM._0383_ ;
 wire \u_cpu.IMEM._0384_ ;
 wire \u_cpu.IMEM._0385_ ;
 wire \u_cpu.IMEM._0386_ ;
 wire \u_cpu.IMEM._0387_ ;
 wire \u_cpu.IMEM._0388_ ;
 wire \u_cpu.IMEM._0389_ ;
 wire \u_cpu.IMEM._0390_ ;
 wire \u_cpu.IMEM._0391_ ;
 wire \u_cpu.IMEM._0392_ ;
 wire \u_cpu.IMEM._0393_ ;
 wire \u_cpu.IMEM._0394_ ;
 wire \u_cpu.IMEM._0395_ ;
 wire \u_cpu.IMEM._0396_ ;
 wire \u_cpu.IMEM._0397_ ;
 wire \u_cpu.IMEM._0398_ ;
 wire \u_cpu.IMEM._0399_ ;
 wire \u_cpu.IMEM._0400_ ;
 wire \u_cpu.IMEM._0401_ ;
 wire \u_cpu.IMEM._0402_ ;
 wire \u_cpu.IMEM._0403_ ;
 wire \u_cpu.IMEM._0404_ ;
 wire \u_cpu.IMEM._0405_ ;
 wire \u_cpu.IMEM._0406_ ;
 wire \u_cpu.IMEM._0407_ ;
 wire \u_cpu.IMEM._0408_ ;
 wire \u_cpu.IMEM._0409_ ;
 wire \u_cpu.IMEM._0410_ ;
 wire \u_cpu.IMEM._0411_ ;
 wire \u_cpu.IMEM._0412_ ;
 wire \u_cpu.IMEM._0413_ ;
 wire \u_cpu.IMEM._0414_ ;
 wire \u_cpu.IMEM._0415_ ;
 wire \u_cpu.IMEM._0416_ ;
 wire \u_cpu.IMEM._0417_ ;
 wire \u_cpu.IMEM._0418_ ;
 wire \u_cpu.IMEM._0419_ ;
 wire \u_cpu.IMEM._0420_ ;
 wire \u_cpu.IMEM._0421_ ;
 wire \u_cpu.IMEM._0422_ ;
 wire \u_cpu.IMEM._0423_ ;
 wire \u_cpu.IMEM._0424_ ;
 wire \u_cpu.IMEM._0425_ ;
 wire \u_cpu.IMEM._0426_ ;
 wire \u_cpu.IMEM._0427_ ;
 wire \u_cpu.IMEM._0428_ ;
 wire \u_cpu.IMEM._0429_ ;
 wire \u_cpu.IMEM._0430_ ;
 wire \u_cpu.IMEM._0431_ ;
 wire \u_cpu.IMEM._0432_ ;
 wire \u_cpu.IMEM._0433_ ;
 wire \u_cpu.IMEM._0434_ ;
 wire \u_cpu.IMEM._0435_ ;
 wire \u_cpu.IMEM._0436_ ;
 wire \u_cpu.IMEM._0437_ ;
 wire \u_cpu.IMEM._0438_ ;
 wire \u_cpu.IMEM._0439_ ;
 wire \u_cpu.IMEM._0440_ ;
 wire \u_cpu.IMEM._0441_ ;
 wire \u_cpu.IMEM._0442_ ;
 wire \u_cpu.IMEM._0443_ ;
 wire \u_cpu.IMEM._0444_ ;
 wire \u_cpu.IMEM._0445_ ;
 wire \u_cpu.IMEM._0446_ ;
 wire \u_cpu.IMEM._0447_ ;
 wire \u_cpu.IMEM._0448_ ;
 wire \u_cpu.IMEM._0449_ ;
 wire \u_cpu.IMEM._0450_ ;
 wire \u_cpu.IMEM._0451_ ;
 wire \u_cpu.IMEM._0452_ ;
 wire \u_cpu.IMEM._0453_ ;
 wire \u_cpu.IMEM._0454_ ;
 wire \u_cpu.IMEM._0455_ ;
 wire \u_cpu.IMEM._0456_ ;
 wire \u_cpu.IMEM._0457_ ;
 wire \u_cpu.IMEM._0458_ ;
 wire \u_cpu.IMEM._0459_ ;
 wire \u_cpu.IMEM._0460_ ;
 wire \u_cpu.IMEM._0461_ ;
 wire \u_cpu.IMEM._0462_ ;
 wire \u_cpu.IMEM._0463_ ;
 wire \u_cpu.IMEM._0464_ ;
 wire \u_cpu.IMEM._0465_ ;
 wire \u_cpu.IMEM._0466_ ;
 wire \u_cpu.IMEM._0467_ ;
 wire \u_cpu.IMEM._0468_ ;
 wire \u_cpu.IMEM._0469_ ;
 wire \u_cpu.IMEM._0470_ ;
 wire \u_cpu.IMEM._0471_ ;
 wire \u_cpu.IMEM._0472_ ;
 wire \u_cpu.IMEM._0473_ ;
 wire \u_cpu.IMEM._0474_ ;
 wire \u_cpu.IMEM._0475_ ;
 wire \u_cpu.IMEM._0476_ ;
 wire \u_cpu.IMEM._0477_ ;
 wire \u_cpu.IMEM._0478_ ;
 wire \u_cpu.IMEM._0479_ ;
 wire \u_cpu.IMEM._0480_ ;
 wire \u_cpu.IMEM._0481_ ;
 wire \u_cpu.IMEM._0482_ ;
 wire \u_cpu.IMEM._0483_ ;
 wire \u_cpu.IMEM._0484_ ;
 wire \u_cpu.IMEM._0485_ ;
 wire \u_cpu.IMEM._0486_ ;
 wire \u_cpu.IMEM._0487_ ;
 wire \u_cpu.IMEM._0488_ ;
 wire \u_cpu.IMEM._0489_ ;
 wire \u_cpu.IMEM._0490_ ;
 wire \u_cpu.IMEM._0491_ ;
 wire \u_cpu.IMEM._0492_ ;
 wire \u_cpu.IMEM._0493_ ;
 wire \u_cpu.IMEM._0494_ ;
 wire \u_cpu.IMEM._0495_ ;
 wire \u_cpu.IMEM._0496_ ;
 wire \u_cpu.IMEM._0497_ ;
 wire \u_cpu.IMEM._0498_ ;
 wire \u_cpu.IMEM._0499_ ;
 wire \u_cpu.IMEM._0500_ ;
 wire \u_cpu.IMEM._0501_ ;
 wire \u_cpu.IMEM._0502_ ;
 wire \u_cpu.IMEM._0503_ ;
 wire \u_cpu.IMEM._0504_ ;
 wire \u_cpu.IMEM._0505_ ;
 wire \u_cpu.IMEM._0506_ ;
 wire \u_cpu.IMEM._0507_ ;
 wire \u_cpu.IMEM._0508_ ;
 wire \u_cpu.IMEM._0509_ ;
 wire \u_cpu.IMEM._0510_ ;
 wire \u_cpu.IMEM._0511_ ;
 wire \u_cpu.IMEM._0512_ ;
 wire \u_cpu.IMEM._0513_ ;
 wire \u_cpu.IMEM._0514_ ;
 wire \u_cpu.IMEM._0515_ ;
 wire \u_cpu.IMEM._0516_ ;
 wire \u_cpu.IMEM._0517_ ;
 wire \u_cpu.IMEM._0518_ ;
 wire \u_cpu.IMEM._0519_ ;
 wire \u_cpu.IMEM._0520_ ;
 wire \u_cpu.IMEM._0521_ ;
 wire \u_cpu.IMEM._0522_ ;
 wire \u_cpu.IMEM._0523_ ;
 wire \u_cpu.IMEM._0524_ ;
 wire \u_cpu.IMEM._0525_ ;
 wire \u_cpu.IMEM._0526_ ;
 wire \u_cpu.IMEM._0527_ ;
 wire \u_cpu.IMEM._0528_ ;
 wire \u_cpu.IMEM._0529_ ;
 wire \u_cpu.IMEM._0530_ ;
 wire \u_cpu.IMEM._0531_ ;
 wire \u_cpu.IMEM._0532_ ;
 wire \u_cpu.IMEM._0533_ ;
 wire \u_cpu.IMEM._0534_ ;
 wire \u_cpu.IMEM._0535_ ;
 wire \u_cpu.IMEM._0536_ ;
 wire \u_cpu.IMEM._0537_ ;
 wire \u_cpu.IMEM._0538_ ;
 wire \u_cpu.IMEM._0539_ ;
 wire \u_cpu.IMEM._0540_ ;
 wire \u_cpu.IMEM._0541_ ;
 wire \u_cpu.IMEM._0542_ ;
 wire \u_cpu.IMEM._0543_ ;
 wire \u_cpu.IMEM._0544_ ;
 wire \u_cpu.IMEM._0545_ ;
 wire \u_cpu.IMEM._0546_ ;
 wire \u_cpu.IMEM._0547_ ;
 wire \u_cpu.IMEM._0548_ ;
 wire \u_cpu.IMEM._0549_ ;
 wire \u_cpu.IMEM._0550_ ;
 wire \u_cpu.IMEM._0551_ ;
 wire \u_cpu.IMEM._0552_ ;
 wire \u_cpu.IMEM._0553_ ;
 wire \u_cpu.IMEM._0554_ ;
 wire \u_cpu.IMEM._0555_ ;
 wire \u_cpu.IMEM._0556_ ;
 wire \u_cpu.IMEM._0557_ ;
 wire \u_cpu.IMEM._0558_ ;
 wire \u_cpu.IMEM._0559_ ;
 wire \u_cpu.IMEM._0560_ ;
 wire \u_cpu.IMEM._0561_ ;
 wire \u_cpu.IMEM._0562_ ;
 wire \u_cpu.IMEM._0563_ ;
 wire \u_cpu.IMEM._0564_ ;
 wire \u_cpu.IMEM._0565_ ;
 wire \u_cpu.IMEM._0566_ ;
 wire \u_cpu.IMEM._0567_ ;
 wire \u_cpu.IMEM._0568_ ;
 wire \u_cpu.IMEM._0569_ ;
 wire \u_cpu.IMEM._0570_ ;
 wire \u_cpu.IMEM._0571_ ;
 wire \u_cpu.IMEM._0572_ ;
 wire \u_cpu.IMEM._0573_ ;
 wire \u_cpu.IMEM._0574_ ;
 wire \u_cpu.IMEM._0575_ ;
 wire \u_cpu.IMEM._0576_ ;
 wire \u_cpu.IMEM._0577_ ;
 wire \u_cpu.IMEM._0578_ ;
 wire \u_cpu.IMEM._0579_ ;
 wire \u_cpu.IMEM._0580_ ;
 wire \u_cpu.IMEM._0581_ ;
 wire \u_cpu.IMEM._0582_ ;
 wire \u_cpu.IMEM._0583_ ;
 wire \u_cpu.IMEM._0584_ ;
 wire \u_cpu.IMEM._0585_ ;
 wire \u_cpu.IMEM._0586_ ;
 wire \u_cpu.IMEM._0587_ ;
 wire \u_cpu.IMEM._0588_ ;
 wire \u_cpu.IMEM._0589_ ;
 wire \u_cpu.IMEM._0590_ ;
 wire \u_cpu.IMEM._0591_ ;
 wire \u_cpu.IMEM._0592_ ;
 wire \u_cpu.IMEM._0593_ ;
 wire \u_cpu.IMEM._0594_ ;
 wire \u_cpu.IMEM._0595_ ;
 wire \u_cpu.IMEM._0596_ ;
 wire \u_cpu.IMEM._0597_ ;
 wire \u_cpu.IMEM._0598_ ;
 wire \u_cpu.IMEM._0599_ ;
 wire \u_cpu.IMEM._0600_ ;
 wire \u_cpu.IMEM._0601_ ;
 wire \u_cpu.IMEM._0602_ ;
 wire \u_cpu.IMEM._0603_ ;
 wire \u_cpu.IMEM._0604_ ;
 wire \u_cpu.IMEM._0605_ ;
 wire \u_cpu.IMEM._0606_ ;
 wire \u_cpu.IMEM._0607_ ;
 wire \u_cpu.IMEM._0608_ ;
 wire \u_cpu.IMEM._0609_ ;
 wire \u_cpu.IMEM._0610_ ;
 wire \u_cpu.IMEM._0611_ ;
 wire \u_cpu.IMEM._0612_ ;
 wire \u_cpu.IMEM._0613_ ;
 wire \u_cpu.IMEM._0614_ ;
 wire \u_cpu.IMEM._0615_ ;
 wire \u_cpu.IMEM._0616_ ;
 wire \u_cpu.IMEM._0617_ ;
 wire \u_cpu.IMEM._0618_ ;
 wire \u_cpu.IMEM._0619_ ;
 wire \u_cpu.IMEM._0620_ ;
 wire \u_cpu.IMEM._0621_ ;
 wire \u_cpu.IMEM._0622_ ;
 wire \u_cpu.IMEM._0623_ ;
 wire \u_cpu.IMEM._0624_ ;
 wire \u_cpu.IMEM._0625_ ;
 wire \u_cpu.IMEM._0626_ ;
 wire \u_cpu.IMEM._0627_ ;
 wire \u_cpu.IMEM._0628_ ;
 wire \u_cpu.IMEM._0629_ ;
 wire \u_cpu.IMEM._0630_ ;
 wire \u_cpu.IMEM._0631_ ;
 wire \u_cpu.IMEM._0632_ ;
 wire \u_cpu.IMEM._0633_ ;
 wire \u_cpu.IMEM._0634_ ;
 wire \u_cpu.IMEM._0635_ ;
 wire \u_cpu.IMEM._0636_ ;
 wire \u_cpu.IMEM._0637_ ;
 wire \u_cpu.IMEM._0638_ ;
 wire \u_cpu.IMEM._0639_ ;
 wire \u_cpu.IMEM._0640_ ;
 wire \u_cpu.IMEM._0641_ ;
 wire \u_cpu.IMEM._0642_ ;
 wire \u_cpu.IMEM._0643_ ;
 wire \u_cpu.IMEM._0644_ ;
 wire \u_cpu.IMEM._0645_ ;
 wire \u_cpu.IMEM._0646_ ;
 wire \u_cpu.IMEM._0647_ ;
 wire \u_cpu.IMEM._0648_ ;
 wire \u_cpu.IMEM._0649_ ;
 wire \u_cpu.IMEM._0650_ ;
 wire \u_cpu.IMEM._0651_ ;
 wire \u_cpu.IMEM._0652_ ;
 wire \u_cpu.IMEM._0653_ ;
 wire \u_cpu.IMEM._0654_ ;
 wire \u_cpu.IMEM._0655_ ;
 wire \u_cpu.IMEM._0656_ ;
 wire \u_cpu.IMEM._0657_ ;
 wire \u_cpu.IMEM._0658_ ;
 wire \u_cpu.IMEM._0659_ ;
 wire \u_cpu.IMEM._0660_ ;
 wire \u_cpu.IMEM._0661_ ;
 wire \u_cpu.IMEM._0662_ ;
 wire \u_cpu.IMEM._0663_ ;
 wire \u_cpu.IMEM._0664_ ;
 wire \u_cpu.IMEM._0665_ ;
 wire \u_cpu.IMEM._0666_ ;
 wire \u_cpu.IMEM._0667_ ;
 wire \u_cpu.IMEM._0668_ ;
 wire \u_cpu.IMEM._0669_ ;
 wire \u_cpu.IMEM._0670_ ;
 wire \u_cpu.IMEM._0671_ ;
 wire \u_cpu.IMEM._0672_ ;
 wire \u_cpu.IMEM._0673_ ;
 wire \u_cpu.IMEM._0674_ ;
 wire \u_cpu.IMEM._0675_ ;
 wire \u_cpu.IMEM._0676_ ;
 wire \u_cpu.IMEM._0677_ ;
 wire \u_cpu.IMEM._0678_ ;
 wire \u_cpu.IMEM._0679_ ;
 wire \u_cpu.IMEM._0680_ ;
 wire \u_cpu.IMEM._0681_ ;
 wire \u_cpu.IMEM._0682_ ;
 wire \u_cpu.IMEM._0683_ ;
 wire \u_cpu.IMEM._0684_ ;
 wire \u_cpu.IMEM._0685_ ;
 wire \u_cpu.IMEM._0686_ ;
 wire \u_cpu.IMEM._0687_ ;
 wire \u_cpu.IMEM._0688_ ;
 wire \u_cpu.IMEM._0689_ ;
 wire \u_cpu.IMEM._0690_ ;
 wire \u_cpu.IMEM._0691_ ;
 wire \u_cpu.IMEM._0692_ ;
 wire \u_cpu.IMEM._0693_ ;
 wire \u_cpu.IMEM._0694_ ;
 wire \u_cpu.IMEM._0695_ ;
 wire \u_cpu.IMEM._0696_ ;
 wire \u_cpu.IMEM._0697_ ;
 wire \u_cpu.IMEM._0698_ ;
 wire \u_cpu.IMEM._0699_ ;
 wire \u_cpu.IMEM._0700_ ;
 wire \u_cpu.IMEM._0701_ ;
 wire \u_cpu.IMEM._0702_ ;
 wire \u_cpu.IMEM._0703_ ;
 wire \u_cpu.IMEM._0704_ ;
 wire \u_cpu.IMEM._0705_ ;
 wire \u_cpu.IMEM._0706_ ;
 wire \u_cpu.IMEM._0707_ ;
 wire \u_cpu.IMEM._0708_ ;
 wire \u_cpu.IMEM._0709_ ;
 wire \u_cpu.IMEM._0710_ ;
 wire \u_cpu.IMEM._0711_ ;
 wire \u_cpu.IMEM._0712_ ;
 wire \u_cpu.IMEM._0713_ ;
 wire \u_cpu.IMEM._0714_ ;
 wire \u_cpu.IMEM._0715_ ;
 wire \u_cpu.IMEM._0716_ ;
 wire \u_cpu.IMEM._0717_ ;
 wire \u_cpu.IMEM._0718_ ;
 wire \u_cpu.IMEM._0719_ ;
 wire \u_cpu.IMEM._0720_ ;
 wire \u_cpu.IMEM._0721_ ;
 wire \u_cpu.IMEM._0722_ ;
 wire \u_cpu.IMEM._0723_ ;
 wire \u_cpu.IMEM._0724_ ;
 wire \u_cpu.IMEM._0725_ ;
 wire \u_cpu.IMEM._0726_ ;
 wire \u_cpu.IMEM._0727_ ;
 wire \u_cpu.IMEM._0728_ ;
 wire \u_cpu.IMEM._0729_ ;
 wire \u_cpu.IMEM._0730_ ;
 wire \u_cpu.IMEM._0731_ ;
 wire \u_cpu.IMEM._0732_ ;
 wire \u_cpu.IMEM._0733_ ;
 wire \u_cpu.IMEM._0734_ ;
 wire \u_cpu.IMEM._0735_ ;
 wire \u_cpu.IMEM._0736_ ;
 wire \u_cpu.IMEM._0737_ ;
 wire \u_cpu.IMEM._0738_ ;
 wire \u_cpu.IMEM._0739_ ;
 wire \u_cpu.IMEM._0740_ ;
 wire \u_cpu.IMEM._0741_ ;
 wire \u_cpu.IMEM._0742_ ;
 wire \u_cpu.IMEM._0743_ ;
 wire \u_cpu.IMEM._0744_ ;
 wire \u_cpu.IMEM._0745_ ;
 wire \u_cpu.IMEM._0746_ ;
 wire \u_cpu.IMEM._0747_ ;
 wire \u_cpu.IMEM._0748_ ;
 wire \u_cpu.IMEM._0749_ ;
 wire \u_cpu.IMEM._0750_ ;
 wire \u_cpu.IMEM._0751_ ;
 wire \u_cpu.IMEM._0752_ ;
 wire \u_cpu.IMEM._0753_ ;
 wire \u_cpu.IMEM._0754_ ;
 wire \u_cpu.IMEM._0755_ ;
 wire \u_cpu.IMEM._0756_ ;
 wire \u_cpu.IMEM._0757_ ;
 wire \u_cpu.IMEM._0758_ ;
 wire \u_cpu.IMEM._0759_ ;
 wire \u_cpu.IMEM._0760_ ;
 wire \u_cpu.IMEM._0761_ ;
 wire \u_cpu.IMEM._0762_ ;
 wire \u_cpu.IMEM._0763_ ;
 wire \u_cpu.IMEM._0764_ ;
 wire \u_cpu.IMEM._0765_ ;
 wire \u_cpu.IMEM._0766_ ;
 wire \u_cpu.IMEM._0767_ ;
 wire \u_cpu.IMEM._0768_ ;
 wire \u_cpu.IMEM._0769_ ;
 wire \u_cpu.IMEM._0770_ ;
 wire \u_cpu.IMEM._0771_ ;
 wire \u_cpu.IMEM._0772_ ;
 wire \u_cpu.IMEM._0773_ ;
 wire \u_cpu.IMEM._0774_ ;
 wire \u_cpu.IMEM._0775_ ;
 wire \u_cpu.IMEM._0776_ ;
 wire \u_cpu.IMEM._0777_ ;
 wire \u_cpu.IMEM._0778_ ;
 wire \u_cpu.IMEM._0779_ ;
 wire \u_cpu.IMEM._0780_ ;
 wire \u_cpu.IMEM._0781_ ;
 wire \u_cpu.IMEM._0782_ ;
 wire \u_cpu.IMEM._0783_ ;
 wire \u_cpu.IMEM._0784_ ;
 wire \u_cpu.IMEM._0785_ ;
 wire \u_cpu.IMEM._0786_ ;
 wire \u_cpu.IMEM._0787_ ;
 wire \u_cpu.IMEM._0788_ ;
 wire \u_cpu.IMEM._0789_ ;
 wire \u_cpu.IMEM._0790_ ;
 wire \u_cpu.IMEM._0791_ ;
 wire \u_cpu.IMEM._0792_ ;
 wire \u_cpu.IMEM._0793_ ;
 wire \u_cpu.IMEM._0794_ ;
 wire \u_cpu.IMEM._0795_ ;
 wire \u_cpu.IMEM._0796_ ;
 wire \u_cpu.IMEM._0797_ ;
 wire \u_cpu.IMEM._0798_ ;
 wire \u_cpu.IMEM._0799_ ;
 wire \u_cpu.IMEM._0800_ ;
 wire \u_cpu.IMEM._0801_ ;
 wire \u_cpu.IMEM._0802_ ;
 wire \u_cpu.IMEM._0803_ ;
 wire \u_cpu.IMEM._0804_ ;
 wire \u_cpu.IMEM._0805_ ;
 wire \u_cpu.IMEM._0806_ ;
 wire \u_cpu.IMEM._0807_ ;
 wire \u_cpu.IMEM._0808_ ;
 wire \u_cpu.IMEM._0809_ ;
 wire \u_cpu.IMEM._0810_ ;
 wire \u_cpu.IMEM._0811_ ;
 wire \u_cpu.IMEM._0812_ ;
 wire \u_cpu.IMEM._0813_ ;
 wire \u_cpu.IMEM._0814_ ;
 wire \u_cpu.IMEM._0815_ ;
 wire \u_cpu.IMEM._0816_ ;
 wire \u_cpu.IMEM._0817_ ;
 wire \u_cpu.IMEM._0818_ ;
 wire \u_cpu.IMEM._0819_ ;
 wire \u_cpu.IMEM._0820_ ;
 wire \u_cpu.IMEM._0821_ ;
 wire \u_cpu.IMEM._0822_ ;
 wire \u_cpu.IMEM._0823_ ;
 wire \u_cpu.IMEM._0824_ ;
 wire \u_cpu.IMEM._0825_ ;
 wire \u_cpu.IMEM._0826_ ;
 wire \u_cpu.IMEM._0827_ ;
 wire \u_cpu.IMEM._0828_ ;
 wire \u_cpu.IMEM._0829_ ;
 wire \u_cpu.IMEM._0830_ ;
 wire \u_cpu.IMEM._0831_ ;
 wire \u_cpu.IMEM._0832_ ;
 wire \u_cpu.IMEM._0833_ ;
 wire \u_cpu.IMEM._0834_ ;
 wire \u_cpu.IMEM._0835_ ;
 wire \u_cpu.IMEM._0836_ ;
 wire \u_cpu.IMEM._0837_ ;
 wire \u_cpu.IMEM._0838_ ;
 wire \u_cpu.IMEM._0839_ ;
 wire \u_cpu.IMEM._0840_ ;
 wire \u_cpu.IMEM._0841_ ;
 wire \u_cpu.IMEM._0842_ ;
 wire \u_cpu.IMEM._0843_ ;
 wire \u_cpu.IMEM._0844_ ;
 wire \u_cpu.IMEM._0845_ ;
 wire \u_cpu.IMEM._0846_ ;
 wire \u_cpu.IMEM._0847_ ;
 wire \u_cpu.IMEM._0848_ ;
 wire \u_cpu.IMEM._0849_ ;
 wire \u_cpu.IMEM._0850_ ;
 wire \u_cpu.IMEM._0851_ ;
 wire \u_cpu.IMEM._0852_ ;
 wire \u_cpu.IMEM._0853_ ;
 wire \u_cpu.IMEM._0854_ ;
 wire \u_cpu.IMEM._0855_ ;
 wire \u_cpu.IMEM._0856_ ;
 wire \u_cpu.IMEM._0857_ ;
 wire \u_cpu.IMEM._0858_ ;
 wire \u_cpu.IMEM._0859_ ;
 wire \u_cpu.IMEM._0860_ ;
 wire \u_cpu.IMEM._0861_ ;
 wire \u_cpu.IMEM._0862_ ;
 wire \u_cpu.IMEM._0863_ ;
 wire \u_cpu.IMEM._0864_ ;
 wire \u_cpu.IMEM._0865_ ;
 wire \u_cpu.IMEM._0866_ ;
 wire \u_cpu.IMEM._0867_ ;
 wire \u_cpu.IMEM._0868_ ;
 wire \u_cpu.IMEM._0869_ ;
 wire \u_cpu.IMEM._0870_ ;
 wire \u_cpu.IMEM._0871_ ;
 wire \u_cpu.IMEM._0872_ ;
 wire \u_cpu.IMEM._0873_ ;
 wire \u_cpu.IMEM._0874_ ;
 wire \u_cpu.IMEM._0875_ ;
 wire \u_cpu.IMEM._0876_ ;
 wire \u_cpu.IMEM._0877_ ;
 wire \u_cpu.IMEM._0878_ ;
 wire \u_cpu.IMEM._0879_ ;
 wire \u_cpu.IMEM._0880_ ;
 wire \u_cpu.IMEM._0881_ ;
 wire \u_cpu.IMEM._0882_ ;
 wire \u_cpu.IMEM._0883_ ;
 wire \u_cpu.IMEM._0884_ ;
 wire \u_cpu.IMEM._0885_ ;
 wire \u_cpu.IMEM._0886_ ;
 wire \u_cpu.IMEM._0887_ ;
 wire \u_cpu.IMEM._0888_ ;
 wire \u_cpu.IMEM._0889_ ;
 wire \u_cpu.IMEM._0890_ ;
 wire \u_cpu.IMEM._0891_ ;
 wire \u_cpu.IMEM._0892_ ;
 wire \u_cpu.IMEM._0893_ ;
 wire \u_cpu.IMEM._0894_ ;
 wire \u_cpu.IMEM._0895_ ;
 wire \u_cpu.IMEM._0896_ ;
 wire \u_cpu.IMEM._0897_ ;
 wire \u_cpu.IMEM._0898_ ;
 wire \u_cpu.IMEM._0899_ ;
 wire \u_cpu.IMEM._0900_ ;
 wire \u_cpu.IMEM._0901_ ;
 wire \u_cpu.IMEM._0902_ ;
 wire \u_cpu.IMEM._0903_ ;
 wire \u_cpu.IMEM._0904_ ;
 wire \u_cpu.IMEM._0905_ ;
 wire \u_cpu.IMEM._0906_ ;
 wire \u_cpu.IMEM._0907_ ;
 wire \u_cpu.IMEM._0908_ ;
 wire \u_cpu.IMEM._0909_ ;
 wire \u_cpu.IMEM._0910_ ;
 wire \u_cpu.IMEM._0911_ ;
 wire \u_cpu.IMEM._0912_ ;
 wire \u_cpu.IMEM._0913_ ;
 wire \u_cpu.IMEM._0914_ ;
 wire \u_cpu.IMEM._0915_ ;
 wire \u_cpu.IMEM._0916_ ;
 wire \u_cpu.IMEM._0917_ ;
 wire \u_cpu.IMEM._0918_ ;
 wire \u_cpu.IMEM._0919_ ;
 wire \u_cpu.IMEM._0920_ ;
 wire \u_cpu.IMEM._0921_ ;
 wire \u_cpu.IMEM._0922_ ;
 wire \u_cpu.IMEM._0923_ ;
 wire \u_cpu.IMEM._0924_ ;
 wire \u_cpu.IMEM._0925_ ;
 wire \u_cpu.IMEM._0926_ ;
 wire \u_cpu.IMEM._0927_ ;
 wire \u_cpu.IMEM.a[10] ;
 wire \u_cpu.IMEM.a[11] ;
 wire \u_cpu.IMEM.a[12] ;
 wire \u_cpu.IMEM.a[13] ;
 wire \u_cpu.IMEM.a[14] ;
 wire \u_cpu.IMEM.a[15] ;
 wire \u_cpu.IMEM.a[16] ;
 wire \u_cpu.IMEM.a[17] ;
 wire \u_cpu.IMEM.a[18] ;
 wire \u_cpu.IMEM.a[19] ;
 wire \u_cpu.IMEM.a[20] ;
 wire \u_cpu.IMEM.a[21] ;
 wire \u_cpu.IMEM.a[22] ;
 wire \u_cpu.IMEM.a[23] ;
 wire \u_cpu.IMEM.a[24] ;
 wire \u_cpu.IMEM.a[25] ;
 wire \u_cpu.IMEM.a[26] ;
 wire \u_cpu.IMEM.a[27] ;
 wire \u_cpu.IMEM.a[28] ;
 wire \u_cpu.IMEM.a[29] ;
 wire \u_cpu.IMEM.a[2] ;
 wire \u_cpu.IMEM.a[30] ;
 wire \u_cpu.IMEM.a[31] ;
 wire \u_cpu.IMEM.a[3] ;
 wire \u_cpu.IMEM.a[4] ;
 wire \u_cpu.IMEM.a[5] ;
 wire \u_cpu.IMEM.a[6] ;
 wire \u_cpu.IMEM.a[7] ;
 wire \u_cpu.IMEM.a[8] ;
 wire \u_cpu.IMEM.a[9] ;
 wire \u_cpu.IMEM.rd[0] ;
 wire \u_cpu.IMEM.rd[10] ;
 wire \u_cpu.IMEM.rd[11] ;
 wire \u_cpu.IMEM.rd[12] ;
 wire \u_cpu.IMEM.rd[13] ;
 wire \u_cpu.IMEM.rd[14] ;
 wire \u_cpu.IMEM.rd[15] ;
 wire \u_cpu.IMEM.rd[16] ;
 wire \u_cpu.IMEM.rd[17] ;
 wire \u_cpu.IMEM.rd[18] ;
 wire \u_cpu.IMEM.rd[19] ;
 wire \u_cpu.IMEM.rd[1] ;
 wire \u_cpu.IMEM.rd[20] ;
 wire \u_cpu.IMEM.rd[21] ;
 wire \u_cpu.IMEM.rd[22] ;
 wire \u_cpu.IMEM.rd[23] ;
 wire \u_cpu.IMEM.rd[24] ;
 wire \u_cpu.IMEM.rd[25] ;
 wire \u_cpu.IMEM.rd[26] ;
 wire \u_cpu.IMEM.rd[27] ;
 wire \u_cpu.IMEM.rd[28] ;
 wire \u_cpu.IMEM.rd[29] ;
 wire \u_cpu.IMEM.rd[2] ;
 wire \u_cpu.IMEM.rd[30] ;
 wire \u_cpu.IMEM.rd[31] ;
 wire \u_cpu.IMEM.rd[3] ;
 wire \u_cpu.IMEM.rd[4] ;
 wire \u_cpu.IMEM.rd[5] ;
 wire \u_cpu.IMEM.rd[6] ;
 wire \u_cpu.IMEM.rd[7] ;
 wire \u_cpu.IMEM.rd[8] ;
 wire \u_cpu.IMEM.rd[9] ;
 wire \u_cpu.M_AXI_AWADDR[0] ;
 wire \u_cpu.M_AXI_AWADDR[10] ;
 wire \u_cpu.M_AXI_AWADDR[11] ;
 wire \u_cpu.M_AXI_AWADDR[12] ;
 wire \u_cpu.M_AXI_AWADDR[13] ;
 wire \u_cpu.M_AXI_AWADDR[14] ;
 wire \u_cpu.M_AXI_AWADDR[15] ;
 wire \u_cpu.M_AXI_AWADDR[16] ;
 wire \u_cpu.M_AXI_AWADDR[17] ;
 wire \u_cpu.M_AXI_AWADDR[18] ;
 wire \u_cpu.M_AXI_AWADDR[19] ;
 wire \u_cpu.M_AXI_AWADDR[1] ;
 wire \u_cpu.M_AXI_AWADDR[20] ;
 wire \u_cpu.M_AXI_AWADDR[21] ;
 wire \u_cpu.M_AXI_AWADDR[22] ;
 wire \u_cpu.M_AXI_AWADDR[23] ;
 wire \u_cpu.M_AXI_AWADDR[24] ;
 wire \u_cpu.M_AXI_AWADDR[25] ;
 wire \u_cpu.M_AXI_AWADDR[26] ;
 wire \u_cpu.M_AXI_AWADDR[27] ;
 wire \u_cpu.M_AXI_AWADDR[28] ;
 wire \u_cpu.M_AXI_AWADDR[29] ;
 wire \u_cpu.M_AXI_AWADDR[2] ;
 wire \u_cpu.M_AXI_AWADDR[30] ;
 wire \u_cpu.M_AXI_AWADDR[31] ;
 wire \u_cpu.M_AXI_AWADDR[3] ;
 wire \u_cpu.M_AXI_AWADDR[4] ;
 wire \u_cpu.M_AXI_AWADDR[5] ;
 wire \u_cpu.M_AXI_AWADDR[6] ;
 wire \u_cpu.M_AXI_AWADDR[7] ;
 wire \u_cpu.M_AXI_AWADDR[8] ;
 wire \u_cpu.M_AXI_AWADDR[9] ;
 wire \u_cpu.M_AXI_WDATA[0] ;
 wire \u_cpu.M_AXI_WDATA[10] ;
 wire \u_cpu.M_AXI_WDATA[11] ;
 wire \u_cpu.M_AXI_WDATA[12] ;
 wire \u_cpu.M_AXI_WDATA[13] ;
 wire \u_cpu.M_AXI_WDATA[14] ;
 wire \u_cpu.M_AXI_WDATA[15] ;
 wire \u_cpu.M_AXI_WDATA[16] ;
 wire \u_cpu.M_AXI_WDATA[17] ;
 wire \u_cpu.M_AXI_WDATA[18] ;
 wire \u_cpu.M_AXI_WDATA[19] ;
 wire \u_cpu.M_AXI_WDATA[1] ;
 wire \u_cpu.M_AXI_WDATA[20] ;
 wire \u_cpu.M_AXI_WDATA[21] ;
 wire \u_cpu.M_AXI_WDATA[22] ;
 wire \u_cpu.M_AXI_WDATA[23] ;
 wire \u_cpu.M_AXI_WDATA[24] ;
 wire \u_cpu.M_AXI_WDATA[25] ;
 wire \u_cpu.M_AXI_WDATA[26] ;
 wire \u_cpu.M_AXI_WDATA[27] ;
 wire \u_cpu.M_AXI_WDATA[28] ;
 wire \u_cpu.M_AXI_WDATA[29] ;
 wire \u_cpu.M_AXI_WDATA[2] ;
 wire \u_cpu.M_AXI_WDATA[30] ;
 wire \u_cpu.M_AXI_WDATA[31] ;
 wire \u_cpu.M_AXI_WDATA[3] ;
 wire \u_cpu.M_AXI_WDATA[4] ;
 wire \u_cpu.M_AXI_WDATA[5] ;
 wire \u_cpu.M_AXI_WDATA[6] ;
 wire \u_cpu.M_AXI_WDATA[7] ;
 wire \u_cpu.M_AXI_WDATA[8] ;
 wire \u_cpu.M_AXI_WDATA[9] ;
 wire \u_cpu.REG_FILE._00000_ ;
 wire \u_cpu.REG_FILE._00001_ ;
 wire \u_cpu.REG_FILE._00002_ ;
 wire \u_cpu.REG_FILE._00003_ ;
 wire \u_cpu.REG_FILE._00004_ ;
 wire \u_cpu.REG_FILE._00005_ ;
 wire \u_cpu.REG_FILE._00006_ ;
 wire \u_cpu.REG_FILE._00007_ ;
 wire \u_cpu.REG_FILE._00008_ ;
 wire \u_cpu.REG_FILE._00009_ ;
 wire \u_cpu.REG_FILE._00010_ ;
 wire \u_cpu.REG_FILE._00011_ ;
 wire \u_cpu.REG_FILE._00012_ ;
 wire \u_cpu.REG_FILE._00013_ ;
 wire \u_cpu.REG_FILE._00014_ ;
 wire \u_cpu.REG_FILE._00015_ ;
 wire \u_cpu.REG_FILE._00016_ ;
 wire \u_cpu.REG_FILE._00017_ ;
 wire \u_cpu.REG_FILE._00018_ ;
 wire \u_cpu.REG_FILE._00019_ ;
 wire \u_cpu.REG_FILE._00020_ ;
 wire \u_cpu.REG_FILE._00021_ ;
 wire \u_cpu.REG_FILE._00022_ ;
 wire \u_cpu.REG_FILE._00023_ ;
 wire \u_cpu.REG_FILE._00024_ ;
 wire \u_cpu.REG_FILE._00025_ ;
 wire \u_cpu.REG_FILE._00026_ ;
 wire \u_cpu.REG_FILE._00027_ ;
 wire \u_cpu.REG_FILE._00028_ ;
 wire \u_cpu.REG_FILE._00029_ ;
 wire \u_cpu.REG_FILE._00030_ ;
 wire \u_cpu.REG_FILE._00031_ ;
 wire \u_cpu.REG_FILE._00032_ ;
 wire \u_cpu.REG_FILE._00033_ ;
 wire \u_cpu.REG_FILE._00034_ ;
 wire \u_cpu.REG_FILE._00035_ ;
 wire \u_cpu.REG_FILE._00036_ ;
 wire \u_cpu.REG_FILE._00037_ ;
 wire \u_cpu.REG_FILE._00038_ ;
 wire \u_cpu.REG_FILE._00039_ ;
 wire \u_cpu.REG_FILE._00040_ ;
 wire \u_cpu.REG_FILE._00041_ ;
 wire \u_cpu.REG_FILE._00042_ ;
 wire \u_cpu.REG_FILE._00043_ ;
 wire \u_cpu.REG_FILE._00044_ ;
 wire \u_cpu.REG_FILE._00045_ ;
 wire \u_cpu.REG_FILE._00046_ ;
 wire \u_cpu.REG_FILE._00047_ ;
 wire \u_cpu.REG_FILE._00048_ ;
 wire \u_cpu.REG_FILE._00049_ ;
 wire \u_cpu.REG_FILE._00050_ ;
 wire \u_cpu.REG_FILE._00051_ ;
 wire \u_cpu.REG_FILE._00052_ ;
 wire \u_cpu.REG_FILE._00053_ ;
 wire \u_cpu.REG_FILE._00054_ ;
 wire \u_cpu.REG_FILE._00055_ ;
 wire \u_cpu.REG_FILE._00056_ ;
 wire \u_cpu.REG_FILE._00057_ ;
 wire \u_cpu.REG_FILE._00058_ ;
 wire \u_cpu.REG_FILE._00059_ ;
 wire \u_cpu.REG_FILE._00060_ ;
 wire \u_cpu.REG_FILE._00061_ ;
 wire \u_cpu.REG_FILE._00062_ ;
 wire \u_cpu.REG_FILE._00063_ ;
 wire \u_cpu.REG_FILE._00064_ ;
 wire \u_cpu.REG_FILE._00065_ ;
 wire \u_cpu.REG_FILE._00066_ ;
 wire \u_cpu.REG_FILE._00067_ ;
 wire \u_cpu.REG_FILE._00068_ ;
 wire \u_cpu.REG_FILE._00069_ ;
 wire \u_cpu.REG_FILE._00070_ ;
 wire \u_cpu.REG_FILE._00071_ ;
 wire \u_cpu.REG_FILE._00072_ ;
 wire \u_cpu.REG_FILE._00073_ ;
 wire \u_cpu.REG_FILE._00074_ ;
 wire \u_cpu.REG_FILE._00075_ ;
 wire \u_cpu.REG_FILE._00076_ ;
 wire \u_cpu.REG_FILE._00077_ ;
 wire \u_cpu.REG_FILE._00078_ ;
 wire \u_cpu.REG_FILE._00079_ ;
 wire \u_cpu.REG_FILE._00080_ ;
 wire \u_cpu.REG_FILE._00081_ ;
 wire \u_cpu.REG_FILE._00082_ ;
 wire \u_cpu.REG_FILE._00083_ ;
 wire \u_cpu.REG_FILE._00084_ ;
 wire \u_cpu.REG_FILE._00085_ ;
 wire \u_cpu.REG_FILE._00086_ ;
 wire \u_cpu.REG_FILE._00087_ ;
 wire \u_cpu.REG_FILE._00088_ ;
 wire \u_cpu.REG_FILE._00089_ ;
 wire \u_cpu.REG_FILE._00090_ ;
 wire \u_cpu.REG_FILE._00091_ ;
 wire \u_cpu.REG_FILE._00092_ ;
 wire \u_cpu.REG_FILE._00093_ ;
 wire \u_cpu.REG_FILE._00094_ ;
 wire \u_cpu.REG_FILE._00095_ ;
 wire \u_cpu.REG_FILE._00096_ ;
 wire \u_cpu.REG_FILE._00097_ ;
 wire \u_cpu.REG_FILE._00098_ ;
 wire \u_cpu.REG_FILE._00099_ ;
 wire \u_cpu.REG_FILE._00100_ ;
 wire \u_cpu.REG_FILE._00101_ ;
 wire \u_cpu.REG_FILE._00102_ ;
 wire \u_cpu.REG_FILE._00103_ ;
 wire \u_cpu.REG_FILE._00104_ ;
 wire \u_cpu.REG_FILE._00105_ ;
 wire \u_cpu.REG_FILE._00106_ ;
 wire \u_cpu.REG_FILE._00107_ ;
 wire \u_cpu.REG_FILE._00108_ ;
 wire \u_cpu.REG_FILE._00109_ ;
 wire \u_cpu.REG_FILE._00110_ ;
 wire \u_cpu.REG_FILE._00111_ ;
 wire \u_cpu.REG_FILE._00112_ ;
 wire \u_cpu.REG_FILE._00113_ ;
 wire \u_cpu.REG_FILE._00114_ ;
 wire \u_cpu.REG_FILE._00115_ ;
 wire \u_cpu.REG_FILE._00116_ ;
 wire \u_cpu.REG_FILE._00117_ ;
 wire \u_cpu.REG_FILE._00118_ ;
 wire \u_cpu.REG_FILE._00119_ ;
 wire \u_cpu.REG_FILE._00120_ ;
 wire \u_cpu.REG_FILE._00121_ ;
 wire \u_cpu.REG_FILE._00122_ ;
 wire \u_cpu.REG_FILE._00123_ ;
 wire \u_cpu.REG_FILE._00124_ ;
 wire \u_cpu.REG_FILE._00125_ ;
 wire \u_cpu.REG_FILE._00126_ ;
 wire \u_cpu.REG_FILE._00127_ ;
 wire \u_cpu.REG_FILE._00128_ ;
 wire \u_cpu.REG_FILE._00129_ ;
 wire \u_cpu.REG_FILE._00130_ ;
 wire \u_cpu.REG_FILE._00131_ ;
 wire \u_cpu.REG_FILE._00132_ ;
 wire \u_cpu.REG_FILE._00133_ ;
 wire \u_cpu.REG_FILE._00134_ ;
 wire \u_cpu.REG_FILE._00135_ ;
 wire \u_cpu.REG_FILE._00136_ ;
 wire \u_cpu.REG_FILE._00137_ ;
 wire \u_cpu.REG_FILE._00138_ ;
 wire \u_cpu.REG_FILE._00139_ ;
 wire \u_cpu.REG_FILE._00140_ ;
 wire \u_cpu.REG_FILE._00141_ ;
 wire \u_cpu.REG_FILE._00142_ ;
 wire \u_cpu.REG_FILE._00143_ ;
 wire \u_cpu.REG_FILE._00144_ ;
 wire \u_cpu.REG_FILE._00145_ ;
 wire \u_cpu.REG_FILE._00146_ ;
 wire \u_cpu.REG_FILE._00147_ ;
 wire \u_cpu.REG_FILE._00148_ ;
 wire \u_cpu.REG_FILE._00149_ ;
 wire \u_cpu.REG_FILE._00150_ ;
 wire \u_cpu.REG_FILE._00151_ ;
 wire \u_cpu.REG_FILE._00152_ ;
 wire \u_cpu.REG_FILE._00153_ ;
 wire \u_cpu.REG_FILE._00154_ ;
 wire \u_cpu.REG_FILE._00155_ ;
 wire \u_cpu.REG_FILE._00156_ ;
 wire \u_cpu.REG_FILE._00157_ ;
 wire \u_cpu.REG_FILE._00158_ ;
 wire \u_cpu.REG_FILE._00159_ ;
 wire \u_cpu.REG_FILE._00160_ ;
 wire \u_cpu.REG_FILE._00161_ ;
 wire \u_cpu.REG_FILE._00162_ ;
 wire \u_cpu.REG_FILE._00163_ ;
 wire \u_cpu.REG_FILE._00164_ ;
 wire \u_cpu.REG_FILE._00165_ ;
 wire \u_cpu.REG_FILE._00166_ ;
 wire \u_cpu.REG_FILE._00167_ ;
 wire \u_cpu.REG_FILE._00168_ ;
 wire \u_cpu.REG_FILE._00169_ ;
 wire \u_cpu.REG_FILE._00170_ ;
 wire \u_cpu.REG_FILE._00171_ ;
 wire \u_cpu.REG_FILE._00172_ ;
 wire \u_cpu.REG_FILE._00173_ ;
 wire \u_cpu.REG_FILE._00174_ ;
 wire \u_cpu.REG_FILE._00175_ ;
 wire \u_cpu.REG_FILE._00176_ ;
 wire \u_cpu.REG_FILE._00177_ ;
 wire \u_cpu.REG_FILE._00178_ ;
 wire \u_cpu.REG_FILE._00179_ ;
 wire \u_cpu.REG_FILE._00180_ ;
 wire \u_cpu.REG_FILE._00181_ ;
 wire \u_cpu.REG_FILE._00182_ ;
 wire \u_cpu.REG_FILE._00183_ ;
 wire \u_cpu.REG_FILE._00184_ ;
 wire \u_cpu.REG_FILE._00185_ ;
 wire \u_cpu.REG_FILE._00186_ ;
 wire \u_cpu.REG_FILE._00187_ ;
 wire \u_cpu.REG_FILE._00188_ ;
 wire \u_cpu.REG_FILE._00189_ ;
 wire \u_cpu.REG_FILE._00190_ ;
 wire \u_cpu.REG_FILE._00191_ ;
 wire \u_cpu.REG_FILE._00192_ ;
 wire \u_cpu.REG_FILE._00193_ ;
 wire \u_cpu.REG_FILE._00194_ ;
 wire \u_cpu.REG_FILE._00195_ ;
 wire \u_cpu.REG_FILE._00196_ ;
 wire \u_cpu.REG_FILE._00197_ ;
 wire \u_cpu.REG_FILE._00198_ ;
 wire \u_cpu.REG_FILE._00199_ ;
 wire \u_cpu.REG_FILE._00200_ ;
 wire \u_cpu.REG_FILE._00201_ ;
 wire \u_cpu.REG_FILE._00202_ ;
 wire \u_cpu.REG_FILE._00203_ ;
 wire \u_cpu.REG_FILE._00204_ ;
 wire \u_cpu.REG_FILE._00205_ ;
 wire \u_cpu.REG_FILE._00206_ ;
 wire \u_cpu.REG_FILE._00207_ ;
 wire \u_cpu.REG_FILE._00208_ ;
 wire \u_cpu.REG_FILE._00209_ ;
 wire \u_cpu.REG_FILE._00210_ ;
 wire \u_cpu.REG_FILE._00211_ ;
 wire \u_cpu.REG_FILE._00212_ ;
 wire \u_cpu.REG_FILE._00213_ ;
 wire \u_cpu.REG_FILE._00214_ ;
 wire \u_cpu.REG_FILE._00215_ ;
 wire \u_cpu.REG_FILE._00216_ ;
 wire \u_cpu.REG_FILE._00217_ ;
 wire \u_cpu.REG_FILE._00218_ ;
 wire \u_cpu.REG_FILE._00219_ ;
 wire \u_cpu.REG_FILE._00220_ ;
 wire \u_cpu.REG_FILE._00221_ ;
 wire \u_cpu.REG_FILE._00222_ ;
 wire \u_cpu.REG_FILE._00223_ ;
 wire \u_cpu.REG_FILE._00224_ ;
 wire \u_cpu.REG_FILE._00225_ ;
 wire \u_cpu.REG_FILE._00226_ ;
 wire \u_cpu.REG_FILE._00227_ ;
 wire \u_cpu.REG_FILE._00228_ ;
 wire \u_cpu.REG_FILE._00229_ ;
 wire \u_cpu.REG_FILE._00230_ ;
 wire \u_cpu.REG_FILE._00231_ ;
 wire \u_cpu.REG_FILE._00232_ ;
 wire \u_cpu.REG_FILE._00233_ ;
 wire \u_cpu.REG_FILE._00234_ ;
 wire \u_cpu.REG_FILE._00235_ ;
 wire \u_cpu.REG_FILE._00236_ ;
 wire \u_cpu.REG_FILE._00237_ ;
 wire \u_cpu.REG_FILE._00238_ ;
 wire \u_cpu.REG_FILE._00239_ ;
 wire \u_cpu.REG_FILE._00240_ ;
 wire \u_cpu.REG_FILE._00241_ ;
 wire \u_cpu.REG_FILE._00242_ ;
 wire \u_cpu.REG_FILE._00243_ ;
 wire \u_cpu.REG_FILE._00244_ ;
 wire \u_cpu.REG_FILE._00245_ ;
 wire \u_cpu.REG_FILE._00246_ ;
 wire \u_cpu.REG_FILE._00247_ ;
 wire \u_cpu.REG_FILE._00248_ ;
 wire \u_cpu.REG_FILE._00249_ ;
 wire \u_cpu.REG_FILE._00250_ ;
 wire \u_cpu.REG_FILE._00251_ ;
 wire \u_cpu.REG_FILE._00252_ ;
 wire \u_cpu.REG_FILE._00253_ ;
 wire \u_cpu.REG_FILE._00254_ ;
 wire \u_cpu.REG_FILE._00255_ ;
 wire \u_cpu.REG_FILE._00256_ ;
 wire \u_cpu.REG_FILE._00257_ ;
 wire \u_cpu.REG_FILE._00258_ ;
 wire \u_cpu.REG_FILE._00259_ ;
 wire \u_cpu.REG_FILE._00260_ ;
 wire \u_cpu.REG_FILE._00261_ ;
 wire \u_cpu.REG_FILE._00262_ ;
 wire \u_cpu.REG_FILE._00263_ ;
 wire \u_cpu.REG_FILE._00264_ ;
 wire \u_cpu.REG_FILE._00265_ ;
 wire \u_cpu.REG_FILE._00266_ ;
 wire \u_cpu.REG_FILE._00267_ ;
 wire \u_cpu.REG_FILE._00268_ ;
 wire \u_cpu.REG_FILE._00269_ ;
 wire \u_cpu.REG_FILE._00270_ ;
 wire \u_cpu.REG_FILE._00271_ ;
 wire \u_cpu.REG_FILE._00272_ ;
 wire \u_cpu.REG_FILE._00273_ ;
 wire \u_cpu.REG_FILE._00274_ ;
 wire \u_cpu.REG_FILE._00275_ ;
 wire \u_cpu.REG_FILE._00276_ ;
 wire \u_cpu.REG_FILE._00277_ ;
 wire \u_cpu.REG_FILE._00278_ ;
 wire \u_cpu.REG_FILE._00279_ ;
 wire \u_cpu.REG_FILE._00280_ ;
 wire \u_cpu.REG_FILE._00281_ ;
 wire \u_cpu.REG_FILE._00282_ ;
 wire \u_cpu.REG_FILE._00283_ ;
 wire \u_cpu.REG_FILE._00284_ ;
 wire \u_cpu.REG_FILE._00285_ ;
 wire \u_cpu.REG_FILE._00286_ ;
 wire \u_cpu.REG_FILE._00287_ ;
 wire \u_cpu.REG_FILE._00288_ ;
 wire \u_cpu.REG_FILE._00289_ ;
 wire \u_cpu.REG_FILE._00290_ ;
 wire \u_cpu.REG_FILE._00291_ ;
 wire \u_cpu.REG_FILE._00292_ ;
 wire \u_cpu.REG_FILE._00293_ ;
 wire \u_cpu.REG_FILE._00294_ ;
 wire \u_cpu.REG_FILE._00295_ ;
 wire \u_cpu.REG_FILE._00296_ ;
 wire \u_cpu.REG_FILE._00297_ ;
 wire \u_cpu.REG_FILE._00298_ ;
 wire \u_cpu.REG_FILE._00299_ ;
 wire \u_cpu.REG_FILE._00300_ ;
 wire \u_cpu.REG_FILE._00301_ ;
 wire \u_cpu.REG_FILE._00302_ ;
 wire \u_cpu.REG_FILE._00303_ ;
 wire \u_cpu.REG_FILE._00304_ ;
 wire \u_cpu.REG_FILE._00305_ ;
 wire \u_cpu.REG_FILE._00306_ ;
 wire \u_cpu.REG_FILE._00307_ ;
 wire \u_cpu.REG_FILE._00308_ ;
 wire \u_cpu.REG_FILE._00309_ ;
 wire \u_cpu.REG_FILE._00310_ ;
 wire \u_cpu.REG_FILE._00311_ ;
 wire \u_cpu.REG_FILE._00312_ ;
 wire \u_cpu.REG_FILE._00313_ ;
 wire \u_cpu.REG_FILE._00314_ ;
 wire \u_cpu.REG_FILE._00315_ ;
 wire \u_cpu.REG_FILE._00316_ ;
 wire \u_cpu.REG_FILE._00317_ ;
 wire \u_cpu.REG_FILE._00318_ ;
 wire \u_cpu.REG_FILE._00319_ ;
 wire \u_cpu.REG_FILE._00320_ ;
 wire \u_cpu.REG_FILE._00321_ ;
 wire \u_cpu.REG_FILE._00322_ ;
 wire \u_cpu.REG_FILE._00323_ ;
 wire \u_cpu.REG_FILE._00324_ ;
 wire \u_cpu.REG_FILE._00325_ ;
 wire \u_cpu.REG_FILE._00326_ ;
 wire \u_cpu.REG_FILE._00327_ ;
 wire \u_cpu.REG_FILE._00328_ ;
 wire \u_cpu.REG_FILE._00329_ ;
 wire \u_cpu.REG_FILE._00330_ ;
 wire \u_cpu.REG_FILE._00331_ ;
 wire \u_cpu.REG_FILE._00332_ ;
 wire \u_cpu.REG_FILE._00333_ ;
 wire \u_cpu.REG_FILE._00334_ ;
 wire \u_cpu.REG_FILE._00335_ ;
 wire \u_cpu.REG_FILE._00336_ ;
 wire \u_cpu.REG_FILE._00337_ ;
 wire \u_cpu.REG_FILE._00338_ ;
 wire \u_cpu.REG_FILE._00339_ ;
 wire \u_cpu.REG_FILE._00340_ ;
 wire \u_cpu.REG_FILE._00341_ ;
 wire \u_cpu.REG_FILE._00342_ ;
 wire \u_cpu.REG_FILE._00343_ ;
 wire \u_cpu.REG_FILE._00344_ ;
 wire \u_cpu.REG_FILE._00345_ ;
 wire \u_cpu.REG_FILE._00346_ ;
 wire \u_cpu.REG_FILE._00347_ ;
 wire \u_cpu.REG_FILE._00348_ ;
 wire \u_cpu.REG_FILE._00349_ ;
 wire \u_cpu.REG_FILE._00350_ ;
 wire \u_cpu.REG_FILE._00351_ ;
 wire \u_cpu.REG_FILE._00352_ ;
 wire \u_cpu.REG_FILE._00353_ ;
 wire \u_cpu.REG_FILE._00354_ ;
 wire \u_cpu.REG_FILE._00355_ ;
 wire \u_cpu.REG_FILE._00356_ ;
 wire \u_cpu.REG_FILE._00357_ ;
 wire \u_cpu.REG_FILE._00358_ ;
 wire \u_cpu.REG_FILE._00359_ ;
 wire \u_cpu.REG_FILE._00360_ ;
 wire \u_cpu.REG_FILE._00361_ ;
 wire \u_cpu.REG_FILE._00362_ ;
 wire \u_cpu.REG_FILE._00363_ ;
 wire \u_cpu.REG_FILE._00364_ ;
 wire \u_cpu.REG_FILE._00365_ ;
 wire \u_cpu.REG_FILE._00366_ ;
 wire \u_cpu.REG_FILE._00367_ ;
 wire \u_cpu.REG_FILE._00368_ ;
 wire \u_cpu.REG_FILE._00369_ ;
 wire \u_cpu.REG_FILE._00370_ ;
 wire \u_cpu.REG_FILE._00371_ ;
 wire \u_cpu.REG_FILE._00372_ ;
 wire \u_cpu.REG_FILE._00373_ ;
 wire \u_cpu.REG_FILE._00374_ ;
 wire \u_cpu.REG_FILE._00375_ ;
 wire \u_cpu.REG_FILE._00376_ ;
 wire \u_cpu.REG_FILE._00377_ ;
 wire \u_cpu.REG_FILE._00378_ ;
 wire \u_cpu.REG_FILE._00379_ ;
 wire \u_cpu.REG_FILE._00380_ ;
 wire \u_cpu.REG_FILE._00381_ ;
 wire \u_cpu.REG_FILE._00382_ ;
 wire \u_cpu.REG_FILE._00383_ ;
 wire \u_cpu.REG_FILE._00384_ ;
 wire \u_cpu.REG_FILE._00385_ ;
 wire \u_cpu.REG_FILE._00386_ ;
 wire \u_cpu.REG_FILE._00387_ ;
 wire \u_cpu.REG_FILE._00388_ ;
 wire \u_cpu.REG_FILE._00389_ ;
 wire \u_cpu.REG_FILE._00390_ ;
 wire \u_cpu.REG_FILE._00391_ ;
 wire \u_cpu.REG_FILE._00392_ ;
 wire \u_cpu.REG_FILE._00393_ ;
 wire \u_cpu.REG_FILE._00394_ ;
 wire \u_cpu.REG_FILE._00395_ ;
 wire \u_cpu.REG_FILE._00396_ ;
 wire \u_cpu.REG_FILE._00397_ ;
 wire \u_cpu.REG_FILE._00398_ ;
 wire \u_cpu.REG_FILE._00399_ ;
 wire \u_cpu.REG_FILE._00400_ ;
 wire \u_cpu.REG_FILE._00401_ ;
 wire \u_cpu.REG_FILE._00402_ ;
 wire \u_cpu.REG_FILE._00403_ ;
 wire \u_cpu.REG_FILE._00404_ ;
 wire \u_cpu.REG_FILE._00405_ ;
 wire \u_cpu.REG_FILE._00406_ ;
 wire \u_cpu.REG_FILE._00407_ ;
 wire \u_cpu.REG_FILE._00408_ ;
 wire \u_cpu.REG_FILE._00409_ ;
 wire \u_cpu.REG_FILE._00410_ ;
 wire \u_cpu.REG_FILE._00411_ ;
 wire \u_cpu.REG_FILE._00412_ ;
 wire \u_cpu.REG_FILE._00413_ ;
 wire \u_cpu.REG_FILE._00414_ ;
 wire \u_cpu.REG_FILE._00415_ ;
 wire \u_cpu.REG_FILE._00416_ ;
 wire \u_cpu.REG_FILE._00417_ ;
 wire \u_cpu.REG_FILE._00418_ ;
 wire \u_cpu.REG_FILE._00419_ ;
 wire \u_cpu.REG_FILE._00420_ ;
 wire \u_cpu.REG_FILE._00421_ ;
 wire \u_cpu.REG_FILE._00422_ ;
 wire \u_cpu.REG_FILE._00423_ ;
 wire \u_cpu.REG_FILE._00424_ ;
 wire \u_cpu.REG_FILE._00425_ ;
 wire \u_cpu.REG_FILE._00426_ ;
 wire \u_cpu.REG_FILE._00427_ ;
 wire \u_cpu.REG_FILE._00428_ ;
 wire \u_cpu.REG_FILE._00429_ ;
 wire \u_cpu.REG_FILE._00430_ ;
 wire \u_cpu.REG_FILE._00431_ ;
 wire \u_cpu.REG_FILE._00432_ ;
 wire \u_cpu.REG_FILE._00433_ ;
 wire \u_cpu.REG_FILE._00434_ ;
 wire \u_cpu.REG_FILE._00435_ ;
 wire \u_cpu.REG_FILE._00436_ ;
 wire \u_cpu.REG_FILE._00437_ ;
 wire \u_cpu.REG_FILE._00438_ ;
 wire \u_cpu.REG_FILE._00439_ ;
 wire \u_cpu.REG_FILE._00440_ ;
 wire \u_cpu.REG_FILE._00441_ ;
 wire \u_cpu.REG_FILE._00442_ ;
 wire \u_cpu.REG_FILE._00443_ ;
 wire \u_cpu.REG_FILE._00444_ ;
 wire \u_cpu.REG_FILE._00445_ ;
 wire \u_cpu.REG_FILE._00446_ ;
 wire \u_cpu.REG_FILE._00447_ ;
 wire \u_cpu.REG_FILE._00448_ ;
 wire \u_cpu.REG_FILE._00449_ ;
 wire \u_cpu.REG_FILE._00450_ ;
 wire \u_cpu.REG_FILE._00451_ ;
 wire \u_cpu.REG_FILE._00452_ ;
 wire \u_cpu.REG_FILE._00453_ ;
 wire \u_cpu.REG_FILE._00454_ ;
 wire \u_cpu.REG_FILE._00455_ ;
 wire \u_cpu.REG_FILE._00456_ ;
 wire \u_cpu.REG_FILE._00457_ ;
 wire \u_cpu.REG_FILE._00458_ ;
 wire \u_cpu.REG_FILE._00459_ ;
 wire \u_cpu.REG_FILE._00460_ ;
 wire \u_cpu.REG_FILE._00461_ ;
 wire \u_cpu.REG_FILE._00462_ ;
 wire \u_cpu.REG_FILE._00463_ ;
 wire \u_cpu.REG_FILE._00464_ ;
 wire \u_cpu.REG_FILE._00465_ ;
 wire \u_cpu.REG_FILE._00466_ ;
 wire \u_cpu.REG_FILE._00467_ ;
 wire \u_cpu.REG_FILE._00468_ ;
 wire \u_cpu.REG_FILE._00469_ ;
 wire \u_cpu.REG_FILE._00470_ ;
 wire \u_cpu.REG_FILE._00471_ ;
 wire \u_cpu.REG_FILE._00472_ ;
 wire \u_cpu.REG_FILE._00473_ ;
 wire \u_cpu.REG_FILE._00474_ ;
 wire \u_cpu.REG_FILE._00475_ ;
 wire \u_cpu.REG_FILE._00476_ ;
 wire \u_cpu.REG_FILE._00477_ ;
 wire \u_cpu.REG_FILE._00478_ ;
 wire \u_cpu.REG_FILE._00479_ ;
 wire \u_cpu.REG_FILE._00480_ ;
 wire \u_cpu.REG_FILE._00481_ ;
 wire \u_cpu.REG_FILE._00482_ ;
 wire \u_cpu.REG_FILE._00483_ ;
 wire \u_cpu.REG_FILE._00484_ ;
 wire \u_cpu.REG_FILE._00485_ ;
 wire \u_cpu.REG_FILE._00486_ ;
 wire \u_cpu.REG_FILE._00487_ ;
 wire \u_cpu.REG_FILE._00488_ ;
 wire \u_cpu.REG_FILE._00489_ ;
 wire \u_cpu.REG_FILE._00490_ ;
 wire \u_cpu.REG_FILE._00491_ ;
 wire \u_cpu.REG_FILE._00492_ ;
 wire \u_cpu.REG_FILE._00493_ ;
 wire \u_cpu.REG_FILE._00494_ ;
 wire \u_cpu.REG_FILE._00495_ ;
 wire \u_cpu.REG_FILE._00496_ ;
 wire \u_cpu.REG_FILE._00497_ ;
 wire \u_cpu.REG_FILE._00498_ ;
 wire \u_cpu.REG_FILE._00499_ ;
 wire \u_cpu.REG_FILE._00500_ ;
 wire \u_cpu.REG_FILE._00501_ ;
 wire \u_cpu.REG_FILE._00502_ ;
 wire \u_cpu.REG_FILE._00503_ ;
 wire \u_cpu.REG_FILE._00504_ ;
 wire \u_cpu.REG_FILE._00505_ ;
 wire \u_cpu.REG_FILE._00506_ ;
 wire \u_cpu.REG_FILE._00507_ ;
 wire \u_cpu.REG_FILE._00508_ ;
 wire \u_cpu.REG_FILE._00509_ ;
 wire \u_cpu.REG_FILE._00510_ ;
 wire \u_cpu.REG_FILE._00511_ ;
 wire \u_cpu.REG_FILE._00512_ ;
 wire \u_cpu.REG_FILE._00513_ ;
 wire \u_cpu.REG_FILE._00514_ ;
 wire \u_cpu.REG_FILE._00515_ ;
 wire \u_cpu.REG_FILE._00516_ ;
 wire \u_cpu.REG_FILE._00517_ ;
 wire \u_cpu.REG_FILE._00518_ ;
 wire \u_cpu.REG_FILE._00519_ ;
 wire \u_cpu.REG_FILE._00520_ ;
 wire \u_cpu.REG_FILE._00521_ ;
 wire \u_cpu.REG_FILE._00522_ ;
 wire \u_cpu.REG_FILE._00523_ ;
 wire \u_cpu.REG_FILE._00524_ ;
 wire \u_cpu.REG_FILE._00525_ ;
 wire \u_cpu.REG_FILE._00526_ ;
 wire \u_cpu.REG_FILE._00527_ ;
 wire \u_cpu.REG_FILE._00528_ ;
 wire \u_cpu.REG_FILE._00529_ ;
 wire \u_cpu.REG_FILE._00530_ ;
 wire \u_cpu.REG_FILE._00531_ ;
 wire \u_cpu.REG_FILE._00532_ ;
 wire \u_cpu.REG_FILE._00533_ ;
 wire \u_cpu.REG_FILE._00534_ ;
 wire \u_cpu.REG_FILE._00535_ ;
 wire \u_cpu.REG_FILE._00536_ ;
 wire \u_cpu.REG_FILE._00537_ ;
 wire \u_cpu.REG_FILE._00538_ ;
 wire \u_cpu.REG_FILE._00539_ ;
 wire \u_cpu.REG_FILE._00540_ ;
 wire \u_cpu.REG_FILE._00541_ ;
 wire \u_cpu.REG_FILE._00542_ ;
 wire \u_cpu.REG_FILE._00543_ ;
 wire \u_cpu.REG_FILE._00544_ ;
 wire \u_cpu.REG_FILE._00545_ ;
 wire \u_cpu.REG_FILE._00546_ ;
 wire \u_cpu.REG_FILE._00547_ ;
 wire \u_cpu.REG_FILE._00548_ ;
 wire \u_cpu.REG_FILE._00549_ ;
 wire \u_cpu.REG_FILE._00550_ ;
 wire \u_cpu.REG_FILE._00551_ ;
 wire \u_cpu.REG_FILE._00552_ ;
 wire \u_cpu.REG_FILE._00553_ ;
 wire \u_cpu.REG_FILE._00554_ ;
 wire \u_cpu.REG_FILE._00555_ ;
 wire \u_cpu.REG_FILE._00556_ ;
 wire \u_cpu.REG_FILE._00557_ ;
 wire \u_cpu.REG_FILE._00558_ ;
 wire \u_cpu.REG_FILE._00559_ ;
 wire \u_cpu.REG_FILE._00560_ ;
 wire \u_cpu.REG_FILE._00561_ ;
 wire \u_cpu.REG_FILE._00562_ ;
 wire \u_cpu.REG_FILE._00563_ ;
 wire \u_cpu.REG_FILE._00564_ ;
 wire \u_cpu.REG_FILE._00565_ ;
 wire \u_cpu.REG_FILE._00566_ ;
 wire \u_cpu.REG_FILE._00567_ ;
 wire \u_cpu.REG_FILE._00568_ ;
 wire \u_cpu.REG_FILE._00569_ ;
 wire \u_cpu.REG_FILE._00570_ ;
 wire \u_cpu.REG_FILE._00571_ ;
 wire \u_cpu.REG_FILE._00572_ ;
 wire \u_cpu.REG_FILE._00573_ ;
 wire \u_cpu.REG_FILE._00574_ ;
 wire \u_cpu.REG_FILE._00575_ ;
 wire \u_cpu.REG_FILE._00576_ ;
 wire \u_cpu.REG_FILE._00577_ ;
 wire \u_cpu.REG_FILE._00578_ ;
 wire \u_cpu.REG_FILE._00579_ ;
 wire \u_cpu.REG_FILE._00580_ ;
 wire \u_cpu.REG_FILE._00581_ ;
 wire \u_cpu.REG_FILE._00582_ ;
 wire \u_cpu.REG_FILE._00583_ ;
 wire \u_cpu.REG_FILE._00584_ ;
 wire \u_cpu.REG_FILE._00585_ ;
 wire \u_cpu.REG_FILE._00586_ ;
 wire \u_cpu.REG_FILE._00587_ ;
 wire \u_cpu.REG_FILE._00588_ ;
 wire \u_cpu.REG_FILE._00589_ ;
 wire \u_cpu.REG_FILE._00590_ ;
 wire \u_cpu.REG_FILE._00591_ ;
 wire \u_cpu.REG_FILE._00592_ ;
 wire \u_cpu.REG_FILE._00593_ ;
 wire \u_cpu.REG_FILE._00594_ ;
 wire \u_cpu.REG_FILE._00595_ ;
 wire \u_cpu.REG_FILE._00596_ ;
 wire \u_cpu.REG_FILE._00597_ ;
 wire \u_cpu.REG_FILE._00598_ ;
 wire \u_cpu.REG_FILE._00599_ ;
 wire \u_cpu.REG_FILE._00600_ ;
 wire \u_cpu.REG_FILE._00601_ ;
 wire \u_cpu.REG_FILE._00602_ ;
 wire \u_cpu.REG_FILE._00603_ ;
 wire \u_cpu.REG_FILE._00604_ ;
 wire \u_cpu.REG_FILE._00605_ ;
 wire \u_cpu.REG_FILE._00606_ ;
 wire \u_cpu.REG_FILE._00607_ ;
 wire \u_cpu.REG_FILE._00608_ ;
 wire \u_cpu.REG_FILE._00609_ ;
 wire \u_cpu.REG_FILE._00610_ ;
 wire \u_cpu.REG_FILE._00611_ ;
 wire \u_cpu.REG_FILE._00612_ ;
 wire \u_cpu.REG_FILE._00613_ ;
 wire \u_cpu.REG_FILE._00614_ ;
 wire \u_cpu.REG_FILE._00615_ ;
 wire \u_cpu.REG_FILE._00616_ ;
 wire \u_cpu.REG_FILE._00617_ ;
 wire \u_cpu.REG_FILE._00618_ ;
 wire \u_cpu.REG_FILE._00619_ ;
 wire \u_cpu.REG_FILE._00620_ ;
 wire \u_cpu.REG_FILE._00621_ ;
 wire \u_cpu.REG_FILE._00622_ ;
 wire \u_cpu.REG_FILE._00623_ ;
 wire \u_cpu.REG_FILE._00624_ ;
 wire \u_cpu.REG_FILE._00625_ ;
 wire \u_cpu.REG_FILE._00626_ ;
 wire \u_cpu.REG_FILE._00627_ ;
 wire \u_cpu.REG_FILE._00628_ ;
 wire \u_cpu.REG_FILE._00629_ ;
 wire \u_cpu.REG_FILE._00630_ ;
 wire \u_cpu.REG_FILE._00631_ ;
 wire \u_cpu.REG_FILE._00632_ ;
 wire \u_cpu.REG_FILE._00633_ ;
 wire \u_cpu.REG_FILE._00634_ ;
 wire \u_cpu.REG_FILE._00635_ ;
 wire \u_cpu.REG_FILE._00636_ ;
 wire \u_cpu.REG_FILE._00637_ ;
 wire \u_cpu.REG_FILE._00638_ ;
 wire \u_cpu.REG_FILE._00639_ ;
 wire \u_cpu.REG_FILE._00640_ ;
 wire \u_cpu.REG_FILE._00641_ ;
 wire \u_cpu.REG_FILE._00642_ ;
 wire \u_cpu.REG_FILE._00643_ ;
 wire \u_cpu.REG_FILE._00644_ ;
 wire \u_cpu.REG_FILE._00645_ ;
 wire \u_cpu.REG_FILE._00646_ ;
 wire \u_cpu.REG_FILE._00647_ ;
 wire \u_cpu.REG_FILE._00648_ ;
 wire \u_cpu.REG_FILE._00649_ ;
 wire \u_cpu.REG_FILE._00650_ ;
 wire \u_cpu.REG_FILE._00651_ ;
 wire \u_cpu.REG_FILE._00652_ ;
 wire \u_cpu.REG_FILE._00653_ ;
 wire \u_cpu.REG_FILE._00654_ ;
 wire \u_cpu.REG_FILE._00655_ ;
 wire \u_cpu.REG_FILE._00656_ ;
 wire \u_cpu.REG_FILE._00657_ ;
 wire \u_cpu.REG_FILE._00658_ ;
 wire \u_cpu.REG_FILE._00659_ ;
 wire \u_cpu.REG_FILE._00660_ ;
 wire \u_cpu.REG_FILE._00661_ ;
 wire \u_cpu.REG_FILE._00662_ ;
 wire \u_cpu.REG_FILE._00663_ ;
 wire \u_cpu.REG_FILE._00664_ ;
 wire \u_cpu.REG_FILE._00665_ ;
 wire \u_cpu.REG_FILE._00666_ ;
 wire \u_cpu.REG_FILE._00667_ ;
 wire \u_cpu.REG_FILE._00668_ ;
 wire \u_cpu.REG_FILE._00669_ ;
 wire \u_cpu.REG_FILE._00670_ ;
 wire \u_cpu.REG_FILE._00671_ ;
 wire \u_cpu.REG_FILE._00672_ ;
 wire \u_cpu.REG_FILE._00673_ ;
 wire \u_cpu.REG_FILE._00674_ ;
 wire \u_cpu.REG_FILE._00675_ ;
 wire \u_cpu.REG_FILE._00676_ ;
 wire \u_cpu.REG_FILE._00677_ ;
 wire \u_cpu.REG_FILE._00678_ ;
 wire \u_cpu.REG_FILE._00679_ ;
 wire \u_cpu.REG_FILE._00680_ ;
 wire \u_cpu.REG_FILE._00681_ ;
 wire \u_cpu.REG_FILE._00682_ ;
 wire \u_cpu.REG_FILE._00683_ ;
 wire \u_cpu.REG_FILE._00684_ ;
 wire \u_cpu.REG_FILE._00685_ ;
 wire \u_cpu.REG_FILE._00686_ ;
 wire \u_cpu.REG_FILE._00687_ ;
 wire \u_cpu.REG_FILE._00688_ ;
 wire \u_cpu.REG_FILE._00689_ ;
 wire \u_cpu.REG_FILE._00690_ ;
 wire \u_cpu.REG_FILE._00691_ ;
 wire \u_cpu.REG_FILE._00692_ ;
 wire \u_cpu.REG_FILE._00693_ ;
 wire \u_cpu.REG_FILE._00694_ ;
 wire \u_cpu.REG_FILE._00695_ ;
 wire \u_cpu.REG_FILE._00696_ ;
 wire \u_cpu.REG_FILE._00697_ ;
 wire \u_cpu.REG_FILE._00698_ ;
 wire \u_cpu.REG_FILE._00699_ ;
 wire \u_cpu.REG_FILE._00700_ ;
 wire \u_cpu.REG_FILE._00701_ ;
 wire \u_cpu.REG_FILE._00702_ ;
 wire \u_cpu.REG_FILE._00703_ ;
 wire \u_cpu.REG_FILE._00704_ ;
 wire \u_cpu.REG_FILE._00705_ ;
 wire \u_cpu.REG_FILE._00706_ ;
 wire \u_cpu.REG_FILE._00707_ ;
 wire \u_cpu.REG_FILE._00708_ ;
 wire \u_cpu.REG_FILE._00709_ ;
 wire \u_cpu.REG_FILE._00710_ ;
 wire \u_cpu.REG_FILE._00711_ ;
 wire \u_cpu.REG_FILE._00712_ ;
 wire \u_cpu.REG_FILE._00713_ ;
 wire \u_cpu.REG_FILE._00714_ ;
 wire \u_cpu.REG_FILE._00715_ ;
 wire \u_cpu.REG_FILE._00716_ ;
 wire \u_cpu.REG_FILE._00717_ ;
 wire \u_cpu.REG_FILE._00718_ ;
 wire \u_cpu.REG_FILE._00719_ ;
 wire \u_cpu.REG_FILE._00720_ ;
 wire \u_cpu.REG_FILE._00721_ ;
 wire \u_cpu.REG_FILE._00722_ ;
 wire \u_cpu.REG_FILE._00723_ ;
 wire \u_cpu.REG_FILE._00724_ ;
 wire \u_cpu.REG_FILE._00725_ ;
 wire \u_cpu.REG_FILE._00726_ ;
 wire \u_cpu.REG_FILE._00727_ ;
 wire \u_cpu.REG_FILE._00728_ ;
 wire \u_cpu.REG_FILE._00729_ ;
 wire \u_cpu.REG_FILE._00730_ ;
 wire \u_cpu.REG_FILE._00731_ ;
 wire \u_cpu.REG_FILE._00732_ ;
 wire \u_cpu.REG_FILE._00733_ ;
 wire \u_cpu.REG_FILE._00734_ ;
 wire \u_cpu.REG_FILE._00735_ ;
 wire \u_cpu.REG_FILE._00736_ ;
 wire \u_cpu.REG_FILE._00737_ ;
 wire \u_cpu.REG_FILE._00738_ ;
 wire \u_cpu.REG_FILE._00739_ ;
 wire \u_cpu.REG_FILE._00740_ ;
 wire \u_cpu.REG_FILE._00741_ ;
 wire \u_cpu.REG_FILE._00742_ ;
 wire \u_cpu.REG_FILE._00743_ ;
 wire \u_cpu.REG_FILE._00744_ ;
 wire \u_cpu.REG_FILE._00745_ ;
 wire \u_cpu.REG_FILE._00746_ ;
 wire \u_cpu.REG_FILE._00747_ ;
 wire \u_cpu.REG_FILE._00748_ ;
 wire \u_cpu.REG_FILE._00749_ ;
 wire \u_cpu.REG_FILE._00750_ ;
 wire \u_cpu.REG_FILE._00751_ ;
 wire \u_cpu.REG_FILE._00752_ ;
 wire \u_cpu.REG_FILE._00753_ ;
 wire \u_cpu.REG_FILE._00754_ ;
 wire \u_cpu.REG_FILE._00755_ ;
 wire \u_cpu.REG_FILE._00756_ ;
 wire \u_cpu.REG_FILE._00757_ ;
 wire \u_cpu.REG_FILE._00758_ ;
 wire \u_cpu.REG_FILE._00759_ ;
 wire \u_cpu.REG_FILE._00760_ ;
 wire \u_cpu.REG_FILE._00761_ ;
 wire \u_cpu.REG_FILE._00762_ ;
 wire \u_cpu.REG_FILE._00763_ ;
 wire \u_cpu.REG_FILE._00764_ ;
 wire \u_cpu.REG_FILE._00765_ ;
 wire \u_cpu.REG_FILE._00766_ ;
 wire \u_cpu.REG_FILE._00767_ ;
 wire \u_cpu.REG_FILE._00768_ ;
 wire \u_cpu.REG_FILE._00769_ ;
 wire \u_cpu.REG_FILE._00770_ ;
 wire \u_cpu.REG_FILE._00771_ ;
 wire \u_cpu.REG_FILE._00772_ ;
 wire \u_cpu.REG_FILE._00773_ ;
 wire \u_cpu.REG_FILE._00774_ ;
 wire \u_cpu.REG_FILE._00775_ ;
 wire \u_cpu.REG_FILE._00776_ ;
 wire \u_cpu.REG_FILE._00777_ ;
 wire \u_cpu.REG_FILE._00778_ ;
 wire \u_cpu.REG_FILE._00779_ ;
 wire \u_cpu.REG_FILE._00780_ ;
 wire \u_cpu.REG_FILE._00781_ ;
 wire \u_cpu.REG_FILE._00782_ ;
 wire \u_cpu.REG_FILE._00783_ ;
 wire \u_cpu.REG_FILE._00784_ ;
 wire \u_cpu.REG_FILE._00785_ ;
 wire \u_cpu.REG_FILE._00786_ ;
 wire \u_cpu.REG_FILE._00787_ ;
 wire \u_cpu.REG_FILE._00788_ ;
 wire \u_cpu.REG_FILE._00789_ ;
 wire \u_cpu.REG_FILE._00790_ ;
 wire \u_cpu.REG_FILE._00791_ ;
 wire \u_cpu.REG_FILE._00792_ ;
 wire \u_cpu.REG_FILE._00793_ ;
 wire \u_cpu.REG_FILE._00794_ ;
 wire \u_cpu.REG_FILE._00795_ ;
 wire \u_cpu.REG_FILE._00796_ ;
 wire \u_cpu.REG_FILE._00797_ ;
 wire \u_cpu.REG_FILE._00798_ ;
 wire \u_cpu.REG_FILE._00799_ ;
 wire \u_cpu.REG_FILE._00800_ ;
 wire \u_cpu.REG_FILE._00801_ ;
 wire \u_cpu.REG_FILE._00802_ ;
 wire \u_cpu.REG_FILE._00803_ ;
 wire \u_cpu.REG_FILE._00804_ ;
 wire \u_cpu.REG_FILE._00805_ ;
 wire \u_cpu.REG_FILE._00806_ ;
 wire \u_cpu.REG_FILE._00807_ ;
 wire \u_cpu.REG_FILE._00808_ ;
 wire \u_cpu.REG_FILE._00809_ ;
 wire \u_cpu.REG_FILE._00810_ ;
 wire \u_cpu.REG_FILE._00811_ ;
 wire \u_cpu.REG_FILE._00812_ ;
 wire \u_cpu.REG_FILE._00813_ ;
 wire \u_cpu.REG_FILE._00814_ ;
 wire \u_cpu.REG_FILE._00815_ ;
 wire \u_cpu.REG_FILE._00816_ ;
 wire \u_cpu.REG_FILE._00817_ ;
 wire \u_cpu.REG_FILE._00818_ ;
 wire \u_cpu.REG_FILE._00819_ ;
 wire \u_cpu.REG_FILE._00820_ ;
 wire \u_cpu.REG_FILE._00821_ ;
 wire \u_cpu.REG_FILE._00822_ ;
 wire \u_cpu.REG_FILE._00823_ ;
 wire \u_cpu.REG_FILE._00824_ ;
 wire \u_cpu.REG_FILE._00825_ ;
 wire \u_cpu.REG_FILE._00826_ ;
 wire \u_cpu.REG_FILE._00827_ ;
 wire \u_cpu.REG_FILE._00828_ ;
 wire \u_cpu.REG_FILE._00829_ ;
 wire \u_cpu.REG_FILE._00830_ ;
 wire \u_cpu.REG_FILE._00831_ ;
 wire \u_cpu.REG_FILE._00832_ ;
 wire \u_cpu.REG_FILE._00833_ ;
 wire \u_cpu.REG_FILE._00834_ ;
 wire \u_cpu.REG_FILE._00835_ ;
 wire \u_cpu.REG_FILE._00836_ ;
 wire \u_cpu.REG_FILE._00837_ ;
 wire \u_cpu.REG_FILE._00838_ ;
 wire \u_cpu.REG_FILE._00839_ ;
 wire \u_cpu.REG_FILE._00840_ ;
 wire \u_cpu.REG_FILE._00841_ ;
 wire \u_cpu.REG_FILE._00842_ ;
 wire \u_cpu.REG_FILE._00843_ ;
 wire \u_cpu.REG_FILE._00844_ ;
 wire \u_cpu.REG_FILE._00845_ ;
 wire \u_cpu.REG_FILE._00846_ ;
 wire \u_cpu.REG_FILE._00847_ ;
 wire \u_cpu.REG_FILE._00848_ ;
 wire \u_cpu.REG_FILE._00849_ ;
 wire \u_cpu.REG_FILE._00850_ ;
 wire \u_cpu.REG_FILE._00851_ ;
 wire \u_cpu.REG_FILE._00852_ ;
 wire \u_cpu.REG_FILE._00853_ ;
 wire \u_cpu.REG_FILE._00854_ ;
 wire \u_cpu.REG_FILE._00855_ ;
 wire \u_cpu.REG_FILE._00856_ ;
 wire \u_cpu.REG_FILE._00857_ ;
 wire \u_cpu.REG_FILE._00858_ ;
 wire \u_cpu.REG_FILE._00859_ ;
 wire \u_cpu.REG_FILE._00860_ ;
 wire \u_cpu.REG_FILE._00861_ ;
 wire \u_cpu.REG_FILE._00862_ ;
 wire \u_cpu.REG_FILE._00863_ ;
 wire \u_cpu.REG_FILE._00864_ ;
 wire \u_cpu.REG_FILE._00865_ ;
 wire \u_cpu.REG_FILE._00866_ ;
 wire \u_cpu.REG_FILE._00867_ ;
 wire \u_cpu.REG_FILE._00868_ ;
 wire \u_cpu.REG_FILE._00869_ ;
 wire \u_cpu.REG_FILE._00870_ ;
 wire \u_cpu.REG_FILE._00871_ ;
 wire \u_cpu.REG_FILE._00872_ ;
 wire \u_cpu.REG_FILE._00873_ ;
 wire \u_cpu.REG_FILE._00874_ ;
 wire \u_cpu.REG_FILE._00875_ ;
 wire \u_cpu.REG_FILE._00876_ ;
 wire \u_cpu.REG_FILE._00877_ ;
 wire \u_cpu.REG_FILE._00878_ ;
 wire \u_cpu.REG_FILE._00879_ ;
 wire \u_cpu.REG_FILE._00880_ ;
 wire \u_cpu.REG_FILE._00881_ ;
 wire \u_cpu.REG_FILE._00882_ ;
 wire \u_cpu.REG_FILE._00883_ ;
 wire \u_cpu.REG_FILE._00884_ ;
 wire \u_cpu.REG_FILE._00885_ ;
 wire \u_cpu.REG_FILE._00886_ ;
 wire \u_cpu.REG_FILE._00887_ ;
 wire \u_cpu.REG_FILE._00888_ ;
 wire \u_cpu.REG_FILE._00889_ ;
 wire \u_cpu.REG_FILE._00890_ ;
 wire \u_cpu.REG_FILE._00891_ ;
 wire \u_cpu.REG_FILE._00892_ ;
 wire \u_cpu.REG_FILE._00893_ ;
 wire \u_cpu.REG_FILE._00894_ ;
 wire \u_cpu.REG_FILE._00895_ ;
 wire \u_cpu.REG_FILE._00896_ ;
 wire \u_cpu.REG_FILE._00897_ ;
 wire \u_cpu.REG_FILE._00898_ ;
 wire \u_cpu.REG_FILE._00899_ ;
 wire \u_cpu.REG_FILE._00900_ ;
 wire \u_cpu.REG_FILE._00901_ ;
 wire \u_cpu.REG_FILE._00902_ ;
 wire \u_cpu.REG_FILE._00903_ ;
 wire \u_cpu.REG_FILE._00904_ ;
 wire \u_cpu.REG_FILE._00905_ ;
 wire \u_cpu.REG_FILE._00906_ ;
 wire \u_cpu.REG_FILE._00907_ ;
 wire \u_cpu.REG_FILE._00908_ ;
 wire \u_cpu.REG_FILE._00909_ ;
 wire \u_cpu.REG_FILE._00910_ ;
 wire \u_cpu.REG_FILE._00911_ ;
 wire \u_cpu.REG_FILE._00912_ ;
 wire \u_cpu.REG_FILE._00913_ ;
 wire \u_cpu.REG_FILE._00914_ ;
 wire \u_cpu.REG_FILE._00915_ ;
 wire \u_cpu.REG_FILE._00916_ ;
 wire \u_cpu.REG_FILE._00917_ ;
 wire \u_cpu.REG_FILE._00918_ ;
 wire \u_cpu.REG_FILE._00919_ ;
 wire \u_cpu.REG_FILE._00920_ ;
 wire \u_cpu.REG_FILE._00921_ ;
 wire \u_cpu.REG_FILE._00922_ ;
 wire \u_cpu.REG_FILE._00923_ ;
 wire \u_cpu.REG_FILE._00924_ ;
 wire \u_cpu.REG_FILE._00925_ ;
 wire \u_cpu.REG_FILE._00926_ ;
 wire \u_cpu.REG_FILE._00927_ ;
 wire \u_cpu.REG_FILE._00928_ ;
 wire \u_cpu.REG_FILE._00929_ ;
 wire \u_cpu.REG_FILE._00930_ ;
 wire \u_cpu.REG_FILE._00931_ ;
 wire \u_cpu.REG_FILE._00932_ ;
 wire \u_cpu.REG_FILE._00933_ ;
 wire \u_cpu.REG_FILE._00934_ ;
 wire \u_cpu.REG_FILE._00935_ ;
 wire \u_cpu.REG_FILE._00936_ ;
 wire \u_cpu.REG_FILE._00937_ ;
 wire \u_cpu.REG_FILE._00938_ ;
 wire \u_cpu.REG_FILE._00939_ ;
 wire \u_cpu.REG_FILE._00940_ ;
 wire \u_cpu.REG_FILE._00941_ ;
 wire \u_cpu.REG_FILE._00942_ ;
 wire \u_cpu.REG_FILE._00943_ ;
 wire \u_cpu.REG_FILE._00944_ ;
 wire \u_cpu.REG_FILE._00945_ ;
 wire \u_cpu.REG_FILE._00946_ ;
 wire \u_cpu.REG_FILE._00947_ ;
 wire \u_cpu.REG_FILE._00948_ ;
 wire \u_cpu.REG_FILE._00949_ ;
 wire \u_cpu.REG_FILE._00950_ ;
 wire \u_cpu.REG_FILE._00951_ ;
 wire \u_cpu.REG_FILE._00952_ ;
 wire \u_cpu.REG_FILE._00953_ ;
 wire \u_cpu.REG_FILE._00954_ ;
 wire \u_cpu.REG_FILE._00955_ ;
 wire \u_cpu.REG_FILE._00956_ ;
 wire \u_cpu.REG_FILE._00957_ ;
 wire \u_cpu.REG_FILE._00958_ ;
 wire \u_cpu.REG_FILE._00959_ ;
 wire \u_cpu.REG_FILE._00960_ ;
 wire \u_cpu.REG_FILE._00961_ ;
 wire \u_cpu.REG_FILE._00962_ ;
 wire \u_cpu.REG_FILE._00963_ ;
 wire \u_cpu.REG_FILE._00964_ ;
 wire \u_cpu.REG_FILE._00965_ ;
 wire \u_cpu.REG_FILE._00966_ ;
 wire \u_cpu.REG_FILE._00967_ ;
 wire \u_cpu.REG_FILE._00968_ ;
 wire \u_cpu.REG_FILE._00969_ ;
 wire \u_cpu.REG_FILE._00970_ ;
 wire \u_cpu.REG_FILE._00971_ ;
 wire \u_cpu.REG_FILE._00972_ ;
 wire \u_cpu.REG_FILE._00973_ ;
 wire \u_cpu.REG_FILE._00974_ ;
 wire \u_cpu.REG_FILE._00975_ ;
 wire \u_cpu.REG_FILE._00976_ ;
 wire \u_cpu.REG_FILE._00977_ ;
 wire \u_cpu.REG_FILE._00978_ ;
 wire \u_cpu.REG_FILE._00979_ ;
 wire \u_cpu.REG_FILE._00980_ ;
 wire \u_cpu.REG_FILE._00981_ ;
 wire \u_cpu.REG_FILE._00982_ ;
 wire \u_cpu.REG_FILE._00983_ ;
 wire \u_cpu.REG_FILE._00984_ ;
 wire \u_cpu.REG_FILE._00985_ ;
 wire \u_cpu.REG_FILE._00986_ ;
 wire \u_cpu.REG_FILE._00987_ ;
 wire \u_cpu.REG_FILE._00988_ ;
 wire \u_cpu.REG_FILE._00989_ ;
 wire \u_cpu.REG_FILE._00990_ ;
 wire \u_cpu.REG_FILE._00991_ ;
 wire \u_cpu.REG_FILE._00992_ ;
 wire \u_cpu.REG_FILE._00993_ ;
 wire \u_cpu.REG_FILE._00994_ ;
 wire \u_cpu.REG_FILE._00995_ ;
 wire \u_cpu.REG_FILE._00996_ ;
 wire \u_cpu.REG_FILE._00997_ ;
 wire \u_cpu.REG_FILE._00998_ ;
 wire \u_cpu.REG_FILE._00999_ ;
 wire \u_cpu.REG_FILE._01000_ ;
 wire \u_cpu.REG_FILE._01001_ ;
 wire \u_cpu.REG_FILE._01002_ ;
 wire \u_cpu.REG_FILE._01003_ ;
 wire \u_cpu.REG_FILE._01004_ ;
 wire \u_cpu.REG_FILE._01005_ ;
 wire \u_cpu.REG_FILE._01006_ ;
 wire \u_cpu.REG_FILE._01007_ ;
 wire \u_cpu.REG_FILE._01008_ ;
 wire \u_cpu.REG_FILE._01009_ ;
 wire \u_cpu.REG_FILE._01010_ ;
 wire \u_cpu.REG_FILE._01011_ ;
 wire \u_cpu.REG_FILE._01012_ ;
 wire \u_cpu.REG_FILE._01013_ ;
 wire \u_cpu.REG_FILE._01014_ ;
 wire \u_cpu.REG_FILE._01015_ ;
 wire \u_cpu.REG_FILE._01016_ ;
 wire \u_cpu.REG_FILE._01017_ ;
 wire \u_cpu.REG_FILE._01018_ ;
 wire \u_cpu.REG_FILE._01019_ ;
 wire \u_cpu.REG_FILE._01020_ ;
 wire \u_cpu.REG_FILE._01021_ ;
 wire \u_cpu.REG_FILE._01022_ ;
 wire \u_cpu.REG_FILE._01023_ ;
 wire \u_cpu.REG_FILE._01024_ ;
 wire \u_cpu.REG_FILE._01025_ ;
 wire \u_cpu.REG_FILE._01026_ ;
 wire \u_cpu.REG_FILE._01027_ ;
 wire \u_cpu.REG_FILE._01028_ ;
 wire \u_cpu.REG_FILE._01029_ ;
 wire \u_cpu.REG_FILE._01030_ ;
 wire \u_cpu.REG_FILE._01031_ ;
 wire \u_cpu.REG_FILE._01032_ ;
 wire \u_cpu.REG_FILE._01033_ ;
 wire \u_cpu.REG_FILE._01034_ ;
 wire \u_cpu.REG_FILE._01035_ ;
 wire \u_cpu.REG_FILE._01036_ ;
 wire \u_cpu.REG_FILE._01037_ ;
 wire \u_cpu.REG_FILE._01038_ ;
 wire \u_cpu.REG_FILE._01039_ ;
 wire \u_cpu.REG_FILE._01040_ ;
 wire \u_cpu.REG_FILE._01041_ ;
 wire \u_cpu.REG_FILE._01042_ ;
 wire \u_cpu.REG_FILE._01043_ ;
 wire \u_cpu.REG_FILE._01044_ ;
 wire \u_cpu.REG_FILE._01045_ ;
 wire \u_cpu.REG_FILE._01046_ ;
 wire \u_cpu.REG_FILE._01047_ ;
 wire \u_cpu.REG_FILE._01048_ ;
 wire \u_cpu.REG_FILE._01049_ ;
 wire \u_cpu.REG_FILE._01050_ ;
 wire \u_cpu.REG_FILE._01051_ ;
 wire \u_cpu.REG_FILE._01052_ ;
 wire \u_cpu.REG_FILE._01053_ ;
 wire \u_cpu.REG_FILE._01054_ ;
 wire \u_cpu.REG_FILE._01055_ ;
 wire \u_cpu.REG_FILE._01056_ ;
 wire \u_cpu.REG_FILE._01057_ ;
 wire \u_cpu.REG_FILE._01058_ ;
 wire \u_cpu.REG_FILE._01059_ ;
 wire \u_cpu.REG_FILE._01060_ ;
 wire \u_cpu.REG_FILE._01061_ ;
 wire \u_cpu.REG_FILE._01062_ ;
 wire \u_cpu.REG_FILE._01063_ ;
 wire \u_cpu.REG_FILE._01064_ ;
 wire \u_cpu.REG_FILE._01065_ ;
 wire \u_cpu.REG_FILE._01066_ ;
 wire \u_cpu.REG_FILE._01067_ ;
 wire \u_cpu.REG_FILE._01068_ ;
 wire \u_cpu.REG_FILE._01069_ ;
 wire \u_cpu.REG_FILE._01070_ ;
 wire \u_cpu.REG_FILE._01071_ ;
 wire \u_cpu.REG_FILE._01072_ ;
 wire \u_cpu.REG_FILE._01073_ ;
 wire \u_cpu.REG_FILE._01074_ ;
 wire \u_cpu.REG_FILE._01075_ ;
 wire \u_cpu.REG_FILE._01076_ ;
 wire \u_cpu.REG_FILE._01077_ ;
 wire \u_cpu.REG_FILE._01078_ ;
 wire \u_cpu.REG_FILE._01079_ ;
 wire \u_cpu.REG_FILE._01080_ ;
 wire \u_cpu.REG_FILE._01081_ ;
 wire \u_cpu.REG_FILE._01082_ ;
 wire \u_cpu.REG_FILE._01083_ ;
 wire \u_cpu.REG_FILE._01084_ ;
 wire \u_cpu.REG_FILE._01085_ ;
 wire \u_cpu.REG_FILE._01086_ ;
 wire \u_cpu.REG_FILE._01087_ ;
 wire \u_cpu.REG_FILE._01088_ ;
 wire \u_cpu.REG_FILE._01089_ ;
 wire \u_cpu.REG_FILE._01090_ ;
 wire \u_cpu.REG_FILE._01091_ ;
 wire \u_cpu.REG_FILE._01092_ ;
 wire \u_cpu.REG_FILE._01093_ ;
 wire \u_cpu.REG_FILE._01094_ ;
 wire \u_cpu.REG_FILE._01095_ ;
 wire \u_cpu.REG_FILE._01096_ ;
 wire \u_cpu.REG_FILE._01097_ ;
 wire \u_cpu.REG_FILE._01098_ ;
 wire \u_cpu.REG_FILE._01099_ ;
 wire \u_cpu.REG_FILE._01100_ ;
 wire \u_cpu.REG_FILE._01101_ ;
 wire \u_cpu.REG_FILE._01102_ ;
 wire \u_cpu.REG_FILE._01103_ ;
 wire \u_cpu.REG_FILE._01104_ ;
 wire \u_cpu.REG_FILE._01105_ ;
 wire \u_cpu.REG_FILE._01106_ ;
 wire \u_cpu.REG_FILE._01107_ ;
 wire \u_cpu.REG_FILE._01108_ ;
 wire \u_cpu.REG_FILE._01109_ ;
 wire \u_cpu.REG_FILE._01110_ ;
 wire \u_cpu.REG_FILE._01111_ ;
 wire \u_cpu.REG_FILE._01112_ ;
 wire \u_cpu.REG_FILE._01113_ ;
 wire \u_cpu.REG_FILE._01114_ ;
 wire \u_cpu.REG_FILE._01115_ ;
 wire \u_cpu.REG_FILE._01116_ ;
 wire \u_cpu.REG_FILE._01117_ ;
 wire \u_cpu.REG_FILE._01118_ ;
 wire \u_cpu.REG_FILE._01119_ ;
 wire \u_cpu.REG_FILE._01120_ ;
 wire \u_cpu.REG_FILE._01121_ ;
 wire \u_cpu.REG_FILE._01122_ ;
 wire \u_cpu.REG_FILE._01123_ ;
 wire \u_cpu.REG_FILE._01124_ ;
 wire \u_cpu.REG_FILE._01125_ ;
 wire \u_cpu.REG_FILE._01126_ ;
 wire \u_cpu.REG_FILE._01127_ ;
 wire \u_cpu.REG_FILE._01128_ ;
 wire \u_cpu.REG_FILE._01129_ ;
 wire \u_cpu.REG_FILE._01130_ ;
 wire \u_cpu.REG_FILE._01131_ ;
 wire \u_cpu.REG_FILE._01132_ ;
 wire \u_cpu.REG_FILE._01133_ ;
 wire \u_cpu.REG_FILE._01134_ ;
 wire \u_cpu.REG_FILE._01135_ ;
 wire \u_cpu.REG_FILE._01136_ ;
 wire \u_cpu.REG_FILE._01137_ ;
 wire \u_cpu.REG_FILE._01138_ ;
 wire \u_cpu.REG_FILE._01139_ ;
 wire \u_cpu.REG_FILE._01140_ ;
 wire \u_cpu.REG_FILE._01141_ ;
 wire \u_cpu.REG_FILE._01142_ ;
 wire \u_cpu.REG_FILE._01143_ ;
 wire \u_cpu.REG_FILE._01144_ ;
 wire \u_cpu.REG_FILE._01145_ ;
 wire \u_cpu.REG_FILE._01146_ ;
 wire \u_cpu.REG_FILE._01147_ ;
 wire \u_cpu.REG_FILE._01148_ ;
 wire \u_cpu.REG_FILE._01149_ ;
 wire \u_cpu.REG_FILE._01150_ ;
 wire \u_cpu.REG_FILE._01151_ ;
 wire \u_cpu.REG_FILE._01152_ ;
 wire \u_cpu.REG_FILE._01153_ ;
 wire \u_cpu.REG_FILE._01154_ ;
 wire \u_cpu.REG_FILE._01155_ ;
 wire \u_cpu.REG_FILE._01156_ ;
 wire \u_cpu.REG_FILE._01157_ ;
 wire \u_cpu.REG_FILE._01158_ ;
 wire \u_cpu.REG_FILE._01159_ ;
 wire \u_cpu.REG_FILE._01160_ ;
 wire \u_cpu.REG_FILE._01161_ ;
 wire \u_cpu.REG_FILE._01162_ ;
 wire \u_cpu.REG_FILE._01163_ ;
 wire \u_cpu.REG_FILE._01164_ ;
 wire \u_cpu.REG_FILE._01165_ ;
 wire \u_cpu.REG_FILE._01166_ ;
 wire \u_cpu.REG_FILE._01167_ ;
 wire \u_cpu.REG_FILE._01168_ ;
 wire \u_cpu.REG_FILE._01169_ ;
 wire \u_cpu.REG_FILE._01170_ ;
 wire \u_cpu.REG_FILE._01171_ ;
 wire \u_cpu.REG_FILE._01172_ ;
 wire \u_cpu.REG_FILE._01173_ ;
 wire \u_cpu.REG_FILE._01174_ ;
 wire \u_cpu.REG_FILE._01175_ ;
 wire \u_cpu.REG_FILE._01176_ ;
 wire \u_cpu.REG_FILE._01177_ ;
 wire \u_cpu.REG_FILE._01178_ ;
 wire \u_cpu.REG_FILE._01179_ ;
 wire \u_cpu.REG_FILE._01180_ ;
 wire \u_cpu.REG_FILE._01181_ ;
 wire \u_cpu.REG_FILE._01182_ ;
 wire \u_cpu.REG_FILE._01183_ ;
 wire \u_cpu.REG_FILE._01184_ ;
 wire \u_cpu.REG_FILE._01185_ ;
 wire \u_cpu.REG_FILE._01186_ ;
 wire \u_cpu.REG_FILE._01187_ ;
 wire \u_cpu.REG_FILE._01188_ ;
 wire \u_cpu.REG_FILE._01189_ ;
 wire \u_cpu.REG_FILE._01190_ ;
 wire \u_cpu.REG_FILE._01191_ ;
 wire \u_cpu.REG_FILE._01192_ ;
 wire \u_cpu.REG_FILE._01193_ ;
 wire \u_cpu.REG_FILE._01194_ ;
 wire \u_cpu.REG_FILE._01195_ ;
 wire \u_cpu.REG_FILE._01196_ ;
 wire \u_cpu.REG_FILE._01197_ ;
 wire \u_cpu.REG_FILE._01198_ ;
 wire \u_cpu.REG_FILE._01199_ ;
 wire \u_cpu.REG_FILE._01200_ ;
 wire \u_cpu.REG_FILE._01201_ ;
 wire \u_cpu.REG_FILE._01202_ ;
 wire \u_cpu.REG_FILE._01203_ ;
 wire \u_cpu.REG_FILE._01204_ ;
 wire \u_cpu.REG_FILE._01205_ ;
 wire \u_cpu.REG_FILE._01206_ ;
 wire \u_cpu.REG_FILE._01207_ ;
 wire \u_cpu.REG_FILE._01208_ ;
 wire \u_cpu.REG_FILE._01209_ ;
 wire \u_cpu.REG_FILE._01210_ ;
 wire \u_cpu.REG_FILE._01211_ ;
 wire \u_cpu.REG_FILE._01212_ ;
 wire \u_cpu.REG_FILE._01213_ ;
 wire \u_cpu.REG_FILE._01214_ ;
 wire \u_cpu.REG_FILE._01215_ ;
 wire \u_cpu.REG_FILE._01216_ ;
 wire \u_cpu.REG_FILE._01217_ ;
 wire \u_cpu.REG_FILE._01218_ ;
 wire \u_cpu.REG_FILE._01219_ ;
 wire \u_cpu.REG_FILE._01220_ ;
 wire \u_cpu.REG_FILE._01221_ ;
 wire \u_cpu.REG_FILE._01222_ ;
 wire \u_cpu.REG_FILE._01223_ ;
 wire \u_cpu.REG_FILE._01224_ ;
 wire \u_cpu.REG_FILE._01225_ ;
 wire \u_cpu.REG_FILE._01226_ ;
 wire \u_cpu.REG_FILE._01227_ ;
 wire \u_cpu.REG_FILE._01228_ ;
 wire \u_cpu.REG_FILE._01229_ ;
 wire \u_cpu.REG_FILE._01230_ ;
 wire \u_cpu.REG_FILE._01231_ ;
 wire \u_cpu.REG_FILE._01232_ ;
 wire \u_cpu.REG_FILE._01233_ ;
 wire \u_cpu.REG_FILE._01234_ ;
 wire \u_cpu.REG_FILE._01235_ ;
 wire \u_cpu.REG_FILE._01236_ ;
 wire \u_cpu.REG_FILE._01237_ ;
 wire \u_cpu.REG_FILE._01238_ ;
 wire \u_cpu.REG_FILE._01239_ ;
 wire \u_cpu.REG_FILE._01240_ ;
 wire \u_cpu.REG_FILE._01241_ ;
 wire \u_cpu.REG_FILE._01242_ ;
 wire \u_cpu.REG_FILE._01243_ ;
 wire \u_cpu.REG_FILE._01244_ ;
 wire \u_cpu.REG_FILE._01245_ ;
 wire \u_cpu.REG_FILE._01246_ ;
 wire \u_cpu.REG_FILE._01247_ ;
 wire \u_cpu.REG_FILE._01248_ ;
 wire \u_cpu.REG_FILE._01249_ ;
 wire \u_cpu.REG_FILE._01250_ ;
 wire \u_cpu.REG_FILE._01251_ ;
 wire \u_cpu.REG_FILE._01252_ ;
 wire \u_cpu.REG_FILE._01253_ ;
 wire \u_cpu.REG_FILE._01254_ ;
 wire \u_cpu.REG_FILE._01255_ ;
 wire \u_cpu.REG_FILE._01256_ ;
 wire \u_cpu.REG_FILE._01257_ ;
 wire \u_cpu.REG_FILE._01258_ ;
 wire \u_cpu.REG_FILE._01259_ ;
 wire \u_cpu.REG_FILE._01260_ ;
 wire \u_cpu.REG_FILE._01261_ ;
 wire \u_cpu.REG_FILE._01262_ ;
 wire \u_cpu.REG_FILE._01263_ ;
 wire \u_cpu.REG_FILE._01264_ ;
 wire \u_cpu.REG_FILE._01265_ ;
 wire \u_cpu.REG_FILE._01266_ ;
 wire \u_cpu.REG_FILE._01267_ ;
 wire \u_cpu.REG_FILE._01268_ ;
 wire \u_cpu.REG_FILE._01269_ ;
 wire \u_cpu.REG_FILE._01270_ ;
 wire \u_cpu.REG_FILE._01271_ ;
 wire \u_cpu.REG_FILE._01272_ ;
 wire \u_cpu.REG_FILE._01273_ ;
 wire \u_cpu.REG_FILE._01274_ ;
 wire \u_cpu.REG_FILE._01275_ ;
 wire \u_cpu.REG_FILE._01276_ ;
 wire \u_cpu.REG_FILE._01277_ ;
 wire \u_cpu.REG_FILE._01278_ ;
 wire \u_cpu.REG_FILE._01279_ ;
 wire \u_cpu.REG_FILE._01280_ ;
 wire \u_cpu.REG_FILE._01281_ ;
 wire \u_cpu.REG_FILE._01282_ ;
 wire \u_cpu.REG_FILE._01283_ ;
 wire \u_cpu.REG_FILE._01284_ ;
 wire \u_cpu.REG_FILE._01285_ ;
 wire \u_cpu.REG_FILE._01286_ ;
 wire \u_cpu.REG_FILE._01287_ ;
 wire \u_cpu.REG_FILE._01288_ ;
 wire \u_cpu.REG_FILE._01289_ ;
 wire \u_cpu.REG_FILE._01290_ ;
 wire \u_cpu.REG_FILE._01291_ ;
 wire \u_cpu.REG_FILE._01292_ ;
 wire \u_cpu.REG_FILE._01293_ ;
 wire \u_cpu.REG_FILE._01294_ ;
 wire \u_cpu.REG_FILE._01295_ ;
 wire \u_cpu.REG_FILE._01296_ ;
 wire \u_cpu.REG_FILE._01297_ ;
 wire \u_cpu.REG_FILE._01298_ ;
 wire \u_cpu.REG_FILE._01299_ ;
 wire \u_cpu.REG_FILE._01300_ ;
 wire \u_cpu.REG_FILE._01301_ ;
 wire \u_cpu.REG_FILE._01302_ ;
 wire \u_cpu.REG_FILE._01303_ ;
 wire \u_cpu.REG_FILE._01304_ ;
 wire \u_cpu.REG_FILE._01305_ ;
 wire \u_cpu.REG_FILE._01306_ ;
 wire \u_cpu.REG_FILE._01307_ ;
 wire \u_cpu.REG_FILE._01308_ ;
 wire \u_cpu.REG_FILE._01309_ ;
 wire \u_cpu.REG_FILE._01310_ ;
 wire \u_cpu.REG_FILE._01311_ ;
 wire \u_cpu.REG_FILE._01312_ ;
 wire \u_cpu.REG_FILE._01313_ ;
 wire \u_cpu.REG_FILE._01314_ ;
 wire \u_cpu.REG_FILE._01315_ ;
 wire \u_cpu.REG_FILE._01316_ ;
 wire \u_cpu.REG_FILE._01317_ ;
 wire \u_cpu.REG_FILE._01318_ ;
 wire \u_cpu.REG_FILE._01319_ ;
 wire \u_cpu.REG_FILE._01320_ ;
 wire \u_cpu.REG_FILE._01321_ ;
 wire \u_cpu.REG_FILE._01322_ ;
 wire \u_cpu.REG_FILE._01323_ ;
 wire \u_cpu.REG_FILE._01324_ ;
 wire \u_cpu.REG_FILE._01325_ ;
 wire \u_cpu.REG_FILE._01326_ ;
 wire \u_cpu.REG_FILE._01327_ ;
 wire \u_cpu.REG_FILE._01328_ ;
 wire \u_cpu.REG_FILE._01329_ ;
 wire \u_cpu.REG_FILE._01330_ ;
 wire \u_cpu.REG_FILE._01331_ ;
 wire \u_cpu.REG_FILE._01332_ ;
 wire \u_cpu.REG_FILE._01333_ ;
 wire \u_cpu.REG_FILE._01334_ ;
 wire \u_cpu.REG_FILE._01335_ ;
 wire \u_cpu.REG_FILE._01336_ ;
 wire \u_cpu.REG_FILE._01337_ ;
 wire \u_cpu.REG_FILE._01338_ ;
 wire \u_cpu.REG_FILE._01339_ ;
 wire \u_cpu.REG_FILE._01340_ ;
 wire \u_cpu.REG_FILE._01341_ ;
 wire \u_cpu.REG_FILE._01342_ ;
 wire \u_cpu.REG_FILE._01343_ ;
 wire \u_cpu.REG_FILE._01344_ ;
 wire \u_cpu.REG_FILE._01345_ ;
 wire \u_cpu.REG_FILE._01346_ ;
 wire \u_cpu.REG_FILE._01347_ ;
 wire \u_cpu.REG_FILE._01348_ ;
 wire \u_cpu.REG_FILE._01349_ ;
 wire \u_cpu.REG_FILE._01350_ ;
 wire \u_cpu.REG_FILE._01351_ ;
 wire \u_cpu.REG_FILE._01352_ ;
 wire \u_cpu.REG_FILE._01353_ ;
 wire \u_cpu.REG_FILE._01354_ ;
 wire \u_cpu.REG_FILE._01355_ ;
 wire \u_cpu.REG_FILE._01356_ ;
 wire \u_cpu.REG_FILE._01357_ ;
 wire \u_cpu.REG_FILE._01358_ ;
 wire \u_cpu.REG_FILE._01359_ ;
 wire \u_cpu.REG_FILE._01360_ ;
 wire \u_cpu.REG_FILE._01361_ ;
 wire \u_cpu.REG_FILE._01362_ ;
 wire \u_cpu.REG_FILE._01363_ ;
 wire \u_cpu.REG_FILE._01364_ ;
 wire \u_cpu.REG_FILE._01365_ ;
 wire \u_cpu.REG_FILE._01366_ ;
 wire \u_cpu.REG_FILE._01367_ ;
 wire \u_cpu.REG_FILE._01368_ ;
 wire \u_cpu.REG_FILE._01369_ ;
 wire \u_cpu.REG_FILE._01370_ ;
 wire \u_cpu.REG_FILE._01371_ ;
 wire \u_cpu.REG_FILE._01372_ ;
 wire \u_cpu.REG_FILE._01373_ ;
 wire \u_cpu.REG_FILE._01374_ ;
 wire \u_cpu.REG_FILE._01375_ ;
 wire \u_cpu.REG_FILE._01376_ ;
 wire \u_cpu.REG_FILE._01377_ ;
 wire \u_cpu.REG_FILE._01378_ ;
 wire \u_cpu.REG_FILE._01379_ ;
 wire \u_cpu.REG_FILE._01380_ ;
 wire \u_cpu.REG_FILE._01381_ ;
 wire \u_cpu.REG_FILE._01382_ ;
 wire \u_cpu.REG_FILE._01383_ ;
 wire \u_cpu.REG_FILE._01384_ ;
 wire \u_cpu.REG_FILE._01385_ ;
 wire \u_cpu.REG_FILE._01386_ ;
 wire \u_cpu.REG_FILE._01387_ ;
 wire \u_cpu.REG_FILE._01388_ ;
 wire \u_cpu.REG_FILE._01389_ ;
 wire \u_cpu.REG_FILE._01390_ ;
 wire \u_cpu.REG_FILE._01391_ ;
 wire \u_cpu.REG_FILE._01392_ ;
 wire \u_cpu.REG_FILE._01393_ ;
 wire \u_cpu.REG_FILE._01394_ ;
 wire \u_cpu.REG_FILE._01395_ ;
 wire \u_cpu.REG_FILE._01396_ ;
 wire \u_cpu.REG_FILE._01397_ ;
 wire \u_cpu.REG_FILE._01398_ ;
 wire \u_cpu.REG_FILE._01399_ ;
 wire \u_cpu.REG_FILE._01400_ ;
 wire \u_cpu.REG_FILE._01401_ ;
 wire \u_cpu.REG_FILE._01402_ ;
 wire \u_cpu.REG_FILE._01403_ ;
 wire \u_cpu.REG_FILE._01404_ ;
 wire \u_cpu.REG_FILE._01405_ ;
 wire \u_cpu.REG_FILE._01406_ ;
 wire \u_cpu.REG_FILE._01407_ ;
 wire \u_cpu.REG_FILE._01408_ ;
 wire \u_cpu.REG_FILE._01409_ ;
 wire \u_cpu.REG_FILE._01410_ ;
 wire \u_cpu.REG_FILE._01411_ ;
 wire \u_cpu.REG_FILE._01412_ ;
 wire \u_cpu.REG_FILE._01413_ ;
 wire \u_cpu.REG_FILE._01414_ ;
 wire \u_cpu.REG_FILE._01415_ ;
 wire \u_cpu.REG_FILE._01416_ ;
 wire \u_cpu.REG_FILE._01417_ ;
 wire \u_cpu.REG_FILE._01418_ ;
 wire \u_cpu.REG_FILE._01419_ ;
 wire \u_cpu.REG_FILE._01420_ ;
 wire \u_cpu.REG_FILE._01421_ ;
 wire \u_cpu.REG_FILE._01422_ ;
 wire \u_cpu.REG_FILE._01423_ ;
 wire \u_cpu.REG_FILE._01424_ ;
 wire \u_cpu.REG_FILE._01425_ ;
 wire \u_cpu.REG_FILE._01426_ ;
 wire \u_cpu.REG_FILE._01427_ ;
 wire \u_cpu.REG_FILE._01428_ ;
 wire \u_cpu.REG_FILE._01429_ ;
 wire \u_cpu.REG_FILE._01430_ ;
 wire \u_cpu.REG_FILE._01431_ ;
 wire \u_cpu.REG_FILE._01432_ ;
 wire \u_cpu.REG_FILE._01433_ ;
 wire \u_cpu.REG_FILE._01434_ ;
 wire \u_cpu.REG_FILE._01435_ ;
 wire \u_cpu.REG_FILE._01436_ ;
 wire \u_cpu.REG_FILE._01437_ ;
 wire \u_cpu.REG_FILE._01438_ ;
 wire \u_cpu.REG_FILE._01439_ ;
 wire \u_cpu.REG_FILE._01440_ ;
 wire \u_cpu.REG_FILE._01441_ ;
 wire \u_cpu.REG_FILE._01442_ ;
 wire \u_cpu.REG_FILE._01443_ ;
 wire \u_cpu.REG_FILE._01444_ ;
 wire \u_cpu.REG_FILE._01445_ ;
 wire \u_cpu.REG_FILE._01446_ ;
 wire \u_cpu.REG_FILE._01447_ ;
 wire \u_cpu.REG_FILE._01448_ ;
 wire \u_cpu.REG_FILE._01449_ ;
 wire \u_cpu.REG_FILE._01450_ ;
 wire \u_cpu.REG_FILE._01451_ ;
 wire \u_cpu.REG_FILE._01452_ ;
 wire \u_cpu.REG_FILE._01453_ ;
 wire \u_cpu.REG_FILE._01454_ ;
 wire \u_cpu.REG_FILE._01455_ ;
 wire \u_cpu.REG_FILE._01456_ ;
 wire \u_cpu.REG_FILE._01457_ ;
 wire \u_cpu.REG_FILE._01458_ ;
 wire \u_cpu.REG_FILE._01459_ ;
 wire \u_cpu.REG_FILE._01460_ ;
 wire \u_cpu.REG_FILE._01461_ ;
 wire \u_cpu.REG_FILE._01462_ ;
 wire \u_cpu.REG_FILE._01463_ ;
 wire \u_cpu.REG_FILE._01464_ ;
 wire \u_cpu.REG_FILE._01465_ ;
 wire \u_cpu.REG_FILE._01466_ ;
 wire \u_cpu.REG_FILE._01467_ ;
 wire \u_cpu.REG_FILE._01468_ ;
 wire \u_cpu.REG_FILE._01469_ ;
 wire \u_cpu.REG_FILE._01470_ ;
 wire \u_cpu.REG_FILE._01471_ ;
 wire \u_cpu.REG_FILE._01472_ ;
 wire \u_cpu.REG_FILE._01473_ ;
 wire \u_cpu.REG_FILE._01474_ ;
 wire \u_cpu.REG_FILE._01475_ ;
 wire \u_cpu.REG_FILE._01476_ ;
 wire \u_cpu.REG_FILE._01477_ ;
 wire \u_cpu.REG_FILE._01478_ ;
 wire \u_cpu.REG_FILE._01479_ ;
 wire \u_cpu.REG_FILE._01480_ ;
 wire \u_cpu.REG_FILE._01481_ ;
 wire \u_cpu.REG_FILE._01482_ ;
 wire \u_cpu.REG_FILE._01483_ ;
 wire \u_cpu.REG_FILE._01484_ ;
 wire \u_cpu.REG_FILE._01485_ ;
 wire \u_cpu.REG_FILE._01486_ ;
 wire \u_cpu.REG_FILE._01487_ ;
 wire \u_cpu.REG_FILE._01488_ ;
 wire \u_cpu.REG_FILE._01489_ ;
 wire \u_cpu.REG_FILE._01490_ ;
 wire \u_cpu.REG_FILE._01491_ ;
 wire \u_cpu.REG_FILE._01492_ ;
 wire \u_cpu.REG_FILE._01493_ ;
 wire \u_cpu.REG_FILE._01494_ ;
 wire \u_cpu.REG_FILE._01495_ ;
 wire \u_cpu.REG_FILE._01496_ ;
 wire \u_cpu.REG_FILE._01497_ ;
 wire \u_cpu.REG_FILE._01498_ ;
 wire \u_cpu.REG_FILE._01499_ ;
 wire \u_cpu.REG_FILE._01500_ ;
 wire \u_cpu.REG_FILE._01501_ ;
 wire \u_cpu.REG_FILE._01502_ ;
 wire \u_cpu.REG_FILE._01503_ ;
 wire \u_cpu.REG_FILE._01504_ ;
 wire \u_cpu.REG_FILE._01505_ ;
 wire \u_cpu.REG_FILE._01506_ ;
 wire \u_cpu.REG_FILE._01507_ ;
 wire \u_cpu.REG_FILE._01508_ ;
 wire \u_cpu.REG_FILE._01509_ ;
 wire \u_cpu.REG_FILE._01510_ ;
 wire \u_cpu.REG_FILE._01511_ ;
 wire \u_cpu.REG_FILE._01512_ ;
 wire \u_cpu.REG_FILE._01513_ ;
 wire \u_cpu.REG_FILE._01514_ ;
 wire \u_cpu.REG_FILE._01515_ ;
 wire \u_cpu.REG_FILE._01516_ ;
 wire \u_cpu.REG_FILE._01517_ ;
 wire \u_cpu.REG_FILE._01518_ ;
 wire \u_cpu.REG_FILE._01519_ ;
 wire \u_cpu.REG_FILE._01520_ ;
 wire \u_cpu.REG_FILE._01521_ ;
 wire \u_cpu.REG_FILE._01522_ ;
 wire \u_cpu.REG_FILE._01523_ ;
 wire \u_cpu.REG_FILE._01524_ ;
 wire \u_cpu.REG_FILE._01525_ ;
 wire \u_cpu.REG_FILE._01526_ ;
 wire \u_cpu.REG_FILE._01527_ ;
 wire \u_cpu.REG_FILE._01528_ ;
 wire \u_cpu.REG_FILE._01529_ ;
 wire \u_cpu.REG_FILE._01530_ ;
 wire \u_cpu.REG_FILE._01531_ ;
 wire \u_cpu.REG_FILE._01532_ ;
 wire \u_cpu.REG_FILE._01533_ ;
 wire \u_cpu.REG_FILE._01534_ ;
 wire \u_cpu.REG_FILE._01535_ ;
 wire \u_cpu.REG_FILE._01536_ ;
 wire \u_cpu.REG_FILE._01537_ ;
 wire \u_cpu.REG_FILE._01538_ ;
 wire \u_cpu.REG_FILE._01539_ ;
 wire \u_cpu.REG_FILE._01540_ ;
 wire \u_cpu.REG_FILE._01541_ ;
 wire \u_cpu.REG_FILE._01542_ ;
 wire \u_cpu.REG_FILE._01543_ ;
 wire \u_cpu.REG_FILE._01544_ ;
 wire \u_cpu.REG_FILE._01545_ ;
 wire \u_cpu.REG_FILE._01546_ ;
 wire \u_cpu.REG_FILE._01547_ ;
 wire \u_cpu.REG_FILE._01548_ ;
 wire \u_cpu.REG_FILE._01549_ ;
 wire \u_cpu.REG_FILE._01550_ ;
 wire \u_cpu.REG_FILE._01551_ ;
 wire \u_cpu.REG_FILE._01552_ ;
 wire \u_cpu.REG_FILE._01553_ ;
 wire \u_cpu.REG_FILE._01554_ ;
 wire \u_cpu.REG_FILE._01555_ ;
 wire \u_cpu.REG_FILE._01556_ ;
 wire \u_cpu.REG_FILE._01557_ ;
 wire \u_cpu.REG_FILE._01558_ ;
 wire \u_cpu.REG_FILE._01559_ ;
 wire \u_cpu.REG_FILE._01560_ ;
 wire \u_cpu.REG_FILE._01561_ ;
 wire \u_cpu.REG_FILE._01562_ ;
 wire \u_cpu.REG_FILE._01563_ ;
 wire \u_cpu.REG_FILE._01564_ ;
 wire \u_cpu.REG_FILE._01565_ ;
 wire \u_cpu.REG_FILE._01566_ ;
 wire \u_cpu.REG_FILE._01567_ ;
 wire \u_cpu.REG_FILE._01568_ ;
 wire \u_cpu.REG_FILE._01569_ ;
 wire \u_cpu.REG_FILE._01570_ ;
 wire \u_cpu.REG_FILE._01571_ ;
 wire \u_cpu.REG_FILE._01572_ ;
 wire \u_cpu.REG_FILE._01573_ ;
 wire \u_cpu.REG_FILE._01574_ ;
 wire \u_cpu.REG_FILE._01575_ ;
 wire \u_cpu.REG_FILE._01576_ ;
 wire \u_cpu.REG_FILE._01577_ ;
 wire \u_cpu.REG_FILE._01578_ ;
 wire \u_cpu.REG_FILE._01579_ ;
 wire \u_cpu.REG_FILE._01580_ ;
 wire \u_cpu.REG_FILE._01581_ ;
 wire \u_cpu.REG_FILE._01582_ ;
 wire \u_cpu.REG_FILE._01583_ ;
 wire \u_cpu.REG_FILE._01584_ ;
 wire \u_cpu.REG_FILE._01585_ ;
 wire \u_cpu.REG_FILE._01586_ ;
 wire \u_cpu.REG_FILE._01587_ ;
 wire \u_cpu.REG_FILE._01588_ ;
 wire \u_cpu.REG_FILE._01589_ ;
 wire \u_cpu.REG_FILE._01590_ ;
 wire \u_cpu.REG_FILE._01591_ ;
 wire \u_cpu.REG_FILE._01592_ ;
 wire \u_cpu.REG_FILE._01593_ ;
 wire \u_cpu.REG_FILE._01594_ ;
 wire \u_cpu.REG_FILE._01595_ ;
 wire \u_cpu.REG_FILE._01596_ ;
 wire \u_cpu.REG_FILE._01597_ ;
 wire \u_cpu.REG_FILE._01598_ ;
 wire \u_cpu.REG_FILE._01599_ ;
 wire \u_cpu.REG_FILE._01600_ ;
 wire \u_cpu.REG_FILE._01601_ ;
 wire \u_cpu.REG_FILE._01602_ ;
 wire \u_cpu.REG_FILE._01603_ ;
 wire \u_cpu.REG_FILE._01604_ ;
 wire \u_cpu.REG_FILE._01605_ ;
 wire \u_cpu.REG_FILE._01606_ ;
 wire \u_cpu.REG_FILE._01607_ ;
 wire \u_cpu.REG_FILE._01608_ ;
 wire \u_cpu.REG_FILE._01609_ ;
 wire \u_cpu.REG_FILE._01610_ ;
 wire \u_cpu.REG_FILE._01611_ ;
 wire \u_cpu.REG_FILE._01612_ ;
 wire \u_cpu.REG_FILE._01613_ ;
 wire \u_cpu.REG_FILE._01614_ ;
 wire \u_cpu.REG_FILE._01615_ ;
 wire \u_cpu.REG_FILE._01616_ ;
 wire \u_cpu.REG_FILE._01617_ ;
 wire \u_cpu.REG_FILE._01618_ ;
 wire \u_cpu.REG_FILE._01619_ ;
 wire \u_cpu.REG_FILE._01620_ ;
 wire \u_cpu.REG_FILE._01621_ ;
 wire \u_cpu.REG_FILE._01622_ ;
 wire \u_cpu.REG_FILE._01623_ ;
 wire \u_cpu.REG_FILE._01624_ ;
 wire \u_cpu.REG_FILE._01625_ ;
 wire \u_cpu.REG_FILE._01626_ ;
 wire \u_cpu.REG_FILE._01627_ ;
 wire \u_cpu.REG_FILE._01628_ ;
 wire \u_cpu.REG_FILE._01629_ ;
 wire \u_cpu.REG_FILE._01630_ ;
 wire \u_cpu.REG_FILE._01631_ ;
 wire \u_cpu.REG_FILE._01632_ ;
 wire \u_cpu.REG_FILE._01633_ ;
 wire \u_cpu.REG_FILE._01634_ ;
 wire \u_cpu.REG_FILE._01635_ ;
 wire \u_cpu.REG_FILE._01636_ ;
 wire \u_cpu.REG_FILE._01637_ ;
 wire \u_cpu.REG_FILE._01638_ ;
 wire \u_cpu.REG_FILE._01639_ ;
 wire \u_cpu.REG_FILE._01640_ ;
 wire \u_cpu.REG_FILE._01641_ ;
 wire \u_cpu.REG_FILE._01642_ ;
 wire \u_cpu.REG_FILE._01643_ ;
 wire \u_cpu.REG_FILE._01644_ ;
 wire \u_cpu.REG_FILE._01645_ ;
 wire \u_cpu.REG_FILE._01646_ ;
 wire \u_cpu.REG_FILE._01647_ ;
 wire \u_cpu.REG_FILE._01648_ ;
 wire \u_cpu.REG_FILE._01649_ ;
 wire \u_cpu.REG_FILE._01650_ ;
 wire \u_cpu.REG_FILE._01651_ ;
 wire \u_cpu.REG_FILE._01652_ ;
 wire \u_cpu.REG_FILE._01653_ ;
 wire \u_cpu.REG_FILE._01654_ ;
 wire \u_cpu.REG_FILE._01655_ ;
 wire \u_cpu.REG_FILE._01656_ ;
 wire \u_cpu.REG_FILE._01657_ ;
 wire \u_cpu.REG_FILE._01658_ ;
 wire \u_cpu.REG_FILE._01659_ ;
 wire \u_cpu.REG_FILE._01660_ ;
 wire \u_cpu.REG_FILE._01661_ ;
 wire \u_cpu.REG_FILE._01662_ ;
 wire \u_cpu.REG_FILE._01663_ ;
 wire \u_cpu.REG_FILE._01664_ ;
 wire \u_cpu.REG_FILE._01665_ ;
 wire \u_cpu.REG_FILE._01666_ ;
 wire \u_cpu.REG_FILE._01667_ ;
 wire \u_cpu.REG_FILE._01668_ ;
 wire \u_cpu.REG_FILE._01669_ ;
 wire \u_cpu.REG_FILE._01670_ ;
 wire \u_cpu.REG_FILE._01671_ ;
 wire \u_cpu.REG_FILE._01672_ ;
 wire \u_cpu.REG_FILE._01673_ ;
 wire \u_cpu.REG_FILE._01674_ ;
 wire \u_cpu.REG_FILE._01675_ ;
 wire \u_cpu.REG_FILE._01676_ ;
 wire \u_cpu.REG_FILE._01677_ ;
 wire \u_cpu.REG_FILE._01678_ ;
 wire \u_cpu.REG_FILE._01679_ ;
 wire \u_cpu.REG_FILE._01680_ ;
 wire \u_cpu.REG_FILE._01681_ ;
 wire \u_cpu.REG_FILE._01682_ ;
 wire \u_cpu.REG_FILE._01683_ ;
 wire \u_cpu.REG_FILE._01684_ ;
 wire \u_cpu.REG_FILE._01685_ ;
 wire \u_cpu.REG_FILE._01686_ ;
 wire \u_cpu.REG_FILE._01687_ ;
 wire \u_cpu.REG_FILE._01688_ ;
 wire \u_cpu.REG_FILE._01689_ ;
 wire \u_cpu.REG_FILE._01690_ ;
 wire \u_cpu.REG_FILE._01691_ ;
 wire \u_cpu.REG_FILE._01692_ ;
 wire \u_cpu.REG_FILE._01693_ ;
 wire \u_cpu.REG_FILE._01694_ ;
 wire \u_cpu.REG_FILE._01695_ ;
 wire \u_cpu.REG_FILE._01696_ ;
 wire \u_cpu.REG_FILE._01697_ ;
 wire \u_cpu.REG_FILE._01698_ ;
 wire \u_cpu.REG_FILE._01699_ ;
 wire \u_cpu.REG_FILE._01700_ ;
 wire \u_cpu.REG_FILE._01701_ ;
 wire \u_cpu.REG_FILE._01702_ ;
 wire \u_cpu.REG_FILE._01703_ ;
 wire \u_cpu.REG_FILE._01704_ ;
 wire \u_cpu.REG_FILE._01705_ ;
 wire \u_cpu.REG_FILE._01706_ ;
 wire \u_cpu.REG_FILE._01707_ ;
 wire \u_cpu.REG_FILE._01708_ ;
 wire \u_cpu.REG_FILE._01709_ ;
 wire \u_cpu.REG_FILE._01710_ ;
 wire \u_cpu.REG_FILE._01711_ ;
 wire \u_cpu.REG_FILE._01712_ ;
 wire \u_cpu.REG_FILE._01713_ ;
 wire \u_cpu.REG_FILE._01714_ ;
 wire \u_cpu.REG_FILE._01715_ ;
 wire \u_cpu.REG_FILE._01716_ ;
 wire \u_cpu.REG_FILE._01717_ ;
 wire \u_cpu.REG_FILE._01718_ ;
 wire \u_cpu.REG_FILE._01719_ ;
 wire \u_cpu.REG_FILE._01720_ ;
 wire \u_cpu.REG_FILE._01721_ ;
 wire \u_cpu.REG_FILE._01722_ ;
 wire \u_cpu.REG_FILE._01723_ ;
 wire \u_cpu.REG_FILE._01724_ ;
 wire \u_cpu.REG_FILE._01725_ ;
 wire \u_cpu.REG_FILE._01726_ ;
 wire \u_cpu.REG_FILE._01727_ ;
 wire \u_cpu.REG_FILE._01728_ ;
 wire \u_cpu.REG_FILE._01729_ ;
 wire \u_cpu.REG_FILE._01730_ ;
 wire \u_cpu.REG_FILE._01731_ ;
 wire \u_cpu.REG_FILE._01732_ ;
 wire \u_cpu.REG_FILE._01733_ ;
 wire \u_cpu.REG_FILE._01734_ ;
 wire \u_cpu.REG_FILE._01735_ ;
 wire \u_cpu.REG_FILE._01736_ ;
 wire \u_cpu.REG_FILE._01737_ ;
 wire \u_cpu.REG_FILE._01738_ ;
 wire \u_cpu.REG_FILE._01739_ ;
 wire \u_cpu.REG_FILE._01740_ ;
 wire \u_cpu.REG_FILE._01741_ ;
 wire \u_cpu.REG_FILE._01742_ ;
 wire \u_cpu.REG_FILE._01743_ ;
 wire \u_cpu.REG_FILE._01744_ ;
 wire \u_cpu.REG_FILE._01745_ ;
 wire \u_cpu.REG_FILE._01746_ ;
 wire \u_cpu.REG_FILE._01747_ ;
 wire \u_cpu.REG_FILE._01748_ ;
 wire \u_cpu.REG_FILE._01749_ ;
 wire \u_cpu.REG_FILE._01750_ ;
 wire \u_cpu.REG_FILE._01751_ ;
 wire \u_cpu.REG_FILE._01752_ ;
 wire \u_cpu.REG_FILE._01753_ ;
 wire \u_cpu.REG_FILE._01754_ ;
 wire \u_cpu.REG_FILE._01755_ ;
 wire \u_cpu.REG_FILE._01756_ ;
 wire \u_cpu.REG_FILE._01757_ ;
 wire \u_cpu.REG_FILE._01758_ ;
 wire \u_cpu.REG_FILE._01759_ ;
 wire \u_cpu.REG_FILE._01760_ ;
 wire \u_cpu.REG_FILE._01761_ ;
 wire \u_cpu.REG_FILE._01762_ ;
 wire \u_cpu.REG_FILE._01763_ ;
 wire \u_cpu.REG_FILE._01764_ ;
 wire \u_cpu.REG_FILE._01765_ ;
 wire \u_cpu.REG_FILE._01766_ ;
 wire \u_cpu.REG_FILE._01767_ ;
 wire \u_cpu.REG_FILE._01768_ ;
 wire \u_cpu.REG_FILE._01769_ ;
 wire \u_cpu.REG_FILE._01770_ ;
 wire \u_cpu.REG_FILE._01771_ ;
 wire \u_cpu.REG_FILE._01772_ ;
 wire \u_cpu.REG_FILE._01773_ ;
 wire \u_cpu.REG_FILE._01774_ ;
 wire \u_cpu.REG_FILE._01775_ ;
 wire \u_cpu.REG_FILE._01776_ ;
 wire \u_cpu.REG_FILE._01777_ ;
 wire \u_cpu.REG_FILE._01778_ ;
 wire \u_cpu.REG_FILE._01779_ ;
 wire \u_cpu.REG_FILE._01780_ ;
 wire \u_cpu.REG_FILE._01781_ ;
 wire \u_cpu.REG_FILE._01782_ ;
 wire \u_cpu.REG_FILE._01783_ ;
 wire \u_cpu.REG_FILE._01784_ ;
 wire \u_cpu.REG_FILE._01785_ ;
 wire \u_cpu.REG_FILE._01786_ ;
 wire \u_cpu.REG_FILE._01787_ ;
 wire \u_cpu.REG_FILE._01788_ ;
 wire \u_cpu.REG_FILE._01789_ ;
 wire \u_cpu.REG_FILE._01790_ ;
 wire \u_cpu.REG_FILE._01791_ ;
 wire \u_cpu.REG_FILE._01792_ ;
 wire \u_cpu.REG_FILE._01793_ ;
 wire \u_cpu.REG_FILE._01794_ ;
 wire \u_cpu.REG_FILE._01795_ ;
 wire \u_cpu.REG_FILE._01796_ ;
 wire \u_cpu.REG_FILE._01797_ ;
 wire \u_cpu.REG_FILE._01798_ ;
 wire \u_cpu.REG_FILE._01799_ ;
 wire \u_cpu.REG_FILE._01800_ ;
 wire \u_cpu.REG_FILE._01801_ ;
 wire \u_cpu.REG_FILE._01802_ ;
 wire \u_cpu.REG_FILE._01803_ ;
 wire \u_cpu.REG_FILE._01804_ ;
 wire \u_cpu.REG_FILE._01805_ ;
 wire \u_cpu.REG_FILE._01806_ ;
 wire \u_cpu.REG_FILE._01807_ ;
 wire \u_cpu.REG_FILE._01808_ ;
 wire \u_cpu.REG_FILE._01809_ ;
 wire \u_cpu.REG_FILE._01810_ ;
 wire \u_cpu.REG_FILE._01811_ ;
 wire \u_cpu.REG_FILE._01812_ ;
 wire \u_cpu.REG_FILE._01813_ ;
 wire \u_cpu.REG_FILE._01814_ ;
 wire \u_cpu.REG_FILE._01815_ ;
 wire \u_cpu.REG_FILE._01816_ ;
 wire \u_cpu.REG_FILE._01817_ ;
 wire \u_cpu.REG_FILE._01818_ ;
 wire \u_cpu.REG_FILE._01819_ ;
 wire \u_cpu.REG_FILE._01820_ ;
 wire \u_cpu.REG_FILE._01821_ ;
 wire \u_cpu.REG_FILE._01822_ ;
 wire \u_cpu.REG_FILE._01823_ ;
 wire \u_cpu.REG_FILE._01824_ ;
 wire \u_cpu.REG_FILE._01825_ ;
 wire \u_cpu.REG_FILE._01826_ ;
 wire \u_cpu.REG_FILE._01827_ ;
 wire \u_cpu.REG_FILE._01828_ ;
 wire \u_cpu.REG_FILE._01829_ ;
 wire \u_cpu.REG_FILE._01830_ ;
 wire \u_cpu.REG_FILE._01831_ ;
 wire \u_cpu.REG_FILE._01832_ ;
 wire \u_cpu.REG_FILE._01833_ ;
 wire \u_cpu.REG_FILE._01834_ ;
 wire \u_cpu.REG_FILE._01835_ ;
 wire \u_cpu.REG_FILE._01836_ ;
 wire \u_cpu.REG_FILE._01837_ ;
 wire \u_cpu.REG_FILE._01838_ ;
 wire \u_cpu.REG_FILE._01839_ ;
 wire \u_cpu.REG_FILE._01840_ ;
 wire \u_cpu.REG_FILE._01841_ ;
 wire \u_cpu.REG_FILE._01842_ ;
 wire \u_cpu.REG_FILE._01843_ ;
 wire \u_cpu.REG_FILE._01844_ ;
 wire \u_cpu.REG_FILE._01845_ ;
 wire \u_cpu.REG_FILE._01846_ ;
 wire \u_cpu.REG_FILE._01847_ ;
 wire \u_cpu.REG_FILE._01848_ ;
 wire \u_cpu.REG_FILE._01849_ ;
 wire \u_cpu.REG_FILE._01850_ ;
 wire \u_cpu.REG_FILE._01851_ ;
 wire \u_cpu.REG_FILE._01852_ ;
 wire \u_cpu.REG_FILE._01853_ ;
 wire \u_cpu.REG_FILE._01854_ ;
 wire \u_cpu.REG_FILE._01855_ ;
 wire \u_cpu.REG_FILE._01856_ ;
 wire \u_cpu.REG_FILE._01857_ ;
 wire \u_cpu.REG_FILE._01858_ ;
 wire \u_cpu.REG_FILE._01859_ ;
 wire \u_cpu.REG_FILE._01860_ ;
 wire \u_cpu.REG_FILE._01861_ ;
 wire \u_cpu.REG_FILE._01862_ ;
 wire \u_cpu.REG_FILE._01863_ ;
 wire \u_cpu.REG_FILE._01864_ ;
 wire \u_cpu.REG_FILE._01865_ ;
 wire \u_cpu.REG_FILE._01866_ ;
 wire \u_cpu.REG_FILE._01867_ ;
 wire \u_cpu.REG_FILE._01868_ ;
 wire \u_cpu.REG_FILE._01869_ ;
 wire \u_cpu.REG_FILE._01870_ ;
 wire \u_cpu.REG_FILE._01871_ ;
 wire \u_cpu.REG_FILE._01872_ ;
 wire \u_cpu.REG_FILE._01873_ ;
 wire \u_cpu.REG_FILE._01874_ ;
 wire \u_cpu.REG_FILE._01875_ ;
 wire \u_cpu.REG_FILE._01876_ ;
 wire \u_cpu.REG_FILE._01877_ ;
 wire \u_cpu.REG_FILE._01878_ ;
 wire \u_cpu.REG_FILE._01879_ ;
 wire \u_cpu.REG_FILE._01880_ ;
 wire \u_cpu.REG_FILE._01881_ ;
 wire \u_cpu.REG_FILE._01882_ ;
 wire \u_cpu.REG_FILE._01883_ ;
 wire \u_cpu.REG_FILE._01884_ ;
 wire \u_cpu.REG_FILE._01885_ ;
 wire \u_cpu.REG_FILE._01886_ ;
 wire \u_cpu.REG_FILE._01887_ ;
 wire \u_cpu.REG_FILE._01888_ ;
 wire \u_cpu.REG_FILE._01889_ ;
 wire \u_cpu.REG_FILE._01890_ ;
 wire \u_cpu.REG_FILE._01891_ ;
 wire \u_cpu.REG_FILE._01892_ ;
 wire \u_cpu.REG_FILE._01893_ ;
 wire \u_cpu.REG_FILE._01894_ ;
 wire \u_cpu.REG_FILE._01895_ ;
 wire \u_cpu.REG_FILE._01896_ ;
 wire \u_cpu.REG_FILE._01897_ ;
 wire \u_cpu.REG_FILE._01898_ ;
 wire \u_cpu.REG_FILE._01899_ ;
 wire \u_cpu.REG_FILE._01900_ ;
 wire \u_cpu.REG_FILE._01901_ ;
 wire \u_cpu.REG_FILE._01902_ ;
 wire \u_cpu.REG_FILE._01903_ ;
 wire \u_cpu.REG_FILE._01904_ ;
 wire \u_cpu.REG_FILE._01905_ ;
 wire \u_cpu.REG_FILE._01906_ ;
 wire \u_cpu.REG_FILE._01907_ ;
 wire \u_cpu.REG_FILE._01908_ ;
 wire \u_cpu.REG_FILE._01909_ ;
 wire \u_cpu.REG_FILE._01910_ ;
 wire \u_cpu.REG_FILE._01911_ ;
 wire \u_cpu.REG_FILE._01912_ ;
 wire \u_cpu.REG_FILE._01913_ ;
 wire \u_cpu.REG_FILE._01914_ ;
 wire \u_cpu.REG_FILE._01915_ ;
 wire \u_cpu.REG_FILE._01916_ ;
 wire \u_cpu.REG_FILE._01917_ ;
 wire \u_cpu.REG_FILE._01918_ ;
 wire \u_cpu.REG_FILE._01919_ ;
 wire \u_cpu.REG_FILE._01920_ ;
 wire \u_cpu.REG_FILE._01921_ ;
 wire \u_cpu.REG_FILE._01922_ ;
 wire \u_cpu.REG_FILE._01923_ ;
 wire \u_cpu.REG_FILE._01924_ ;
 wire \u_cpu.REG_FILE._01925_ ;
 wire \u_cpu.REG_FILE._01926_ ;
 wire \u_cpu.REG_FILE._01927_ ;
 wire \u_cpu.REG_FILE._01928_ ;
 wire \u_cpu.REG_FILE._01929_ ;
 wire \u_cpu.REG_FILE._01930_ ;
 wire \u_cpu.REG_FILE._01931_ ;
 wire \u_cpu.REG_FILE._01932_ ;
 wire \u_cpu.REG_FILE._01933_ ;
 wire \u_cpu.REG_FILE._01934_ ;
 wire \u_cpu.REG_FILE._01935_ ;
 wire \u_cpu.REG_FILE._01936_ ;
 wire \u_cpu.REG_FILE._01937_ ;
 wire \u_cpu.REG_FILE._01938_ ;
 wire \u_cpu.REG_FILE._01939_ ;
 wire \u_cpu.REG_FILE._01940_ ;
 wire \u_cpu.REG_FILE._01941_ ;
 wire \u_cpu.REG_FILE._01942_ ;
 wire \u_cpu.REG_FILE._01943_ ;
 wire \u_cpu.REG_FILE._01944_ ;
 wire \u_cpu.REG_FILE._01945_ ;
 wire \u_cpu.REG_FILE._01946_ ;
 wire \u_cpu.REG_FILE._01947_ ;
 wire \u_cpu.REG_FILE._01948_ ;
 wire \u_cpu.REG_FILE._01949_ ;
 wire \u_cpu.REG_FILE._01950_ ;
 wire \u_cpu.REG_FILE._01951_ ;
 wire \u_cpu.REG_FILE._01952_ ;
 wire \u_cpu.REG_FILE._01953_ ;
 wire \u_cpu.REG_FILE._01954_ ;
 wire \u_cpu.REG_FILE._01955_ ;
 wire \u_cpu.REG_FILE._01956_ ;
 wire \u_cpu.REG_FILE._01957_ ;
 wire \u_cpu.REG_FILE._01958_ ;
 wire \u_cpu.REG_FILE._01959_ ;
 wire \u_cpu.REG_FILE._01960_ ;
 wire \u_cpu.REG_FILE._01961_ ;
 wire \u_cpu.REG_FILE._01962_ ;
 wire \u_cpu.REG_FILE._01963_ ;
 wire \u_cpu.REG_FILE._01964_ ;
 wire \u_cpu.REG_FILE._01965_ ;
 wire \u_cpu.REG_FILE._01966_ ;
 wire \u_cpu.REG_FILE._01967_ ;
 wire \u_cpu.REG_FILE._01968_ ;
 wire \u_cpu.REG_FILE._01969_ ;
 wire \u_cpu.REG_FILE._01970_ ;
 wire \u_cpu.REG_FILE._01971_ ;
 wire \u_cpu.REG_FILE._01972_ ;
 wire \u_cpu.REG_FILE._01973_ ;
 wire \u_cpu.REG_FILE._01974_ ;
 wire \u_cpu.REG_FILE._01975_ ;
 wire \u_cpu.REG_FILE._01976_ ;
 wire \u_cpu.REG_FILE._01977_ ;
 wire \u_cpu.REG_FILE._01978_ ;
 wire \u_cpu.REG_FILE._01979_ ;
 wire \u_cpu.REG_FILE._01980_ ;
 wire \u_cpu.REG_FILE._01981_ ;
 wire \u_cpu.REG_FILE._01982_ ;
 wire \u_cpu.REG_FILE._01983_ ;
 wire \u_cpu.REG_FILE._01984_ ;
 wire \u_cpu.REG_FILE._01985_ ;
 wire \u_cpu.REG_FILE._01986_ ;
 wire \u_cpu.REG_FILE._01987_ ;
 wire \u_cpu.REG_FILE._01988_ ;
 wire \u_cpu.REG_FILE._01989_ ;
 wire \u_cpu.REG_FILE._01990_ ;
 wire \u_cpu.REG_FILE._01991_ ;
 wire \u_cpu.REG_FILE._01992_ ;
 wire \u_cpu.REG_FILE._01993_ ;
 wire \u_cpu.REG_FILE._01994_ ;
 wire \u_cpu.REG_FILE._01995_ ;
 wire \u_cpu.REG_FILE._01996_ ;
 wire \u_cpu.REG_FILE._01997_ ;
 wire \u_cpu.REG_FILE._01998_ ;
 wire \u_cpu.REG_FILE._01999_ ;
 wire \u_cpu.REG_FILE._02000_ ;
 wire \u_cpu.REG_FILE._02001_ ;
 wire \u_cpu.REG_FILE._02002_ ;
 wire \u_cpu.REG_FILE._02003_ ;
 wire \u_cpu.REG_FILE._02004_ ;
 wire \u_cpu.REG_FILE._02005_ ;
 wire \u_cpu.REG_FILE._02006_ ;
 wire \u_cpu.REG_FILE._02007_ ;
 wire \u_cpu.REG_FILE._02008_ ;
 wire \u_cpu.REG_FILE._02009_ ;
 wire \u_cpu.REG_FILE._02010_ ;
 wire \u_cpu.REG_FILE._02011_ ;
 wire \u_cpu.REG_FILE._02012_ ;
 wire \u_cpu.REG_FILE._02013_ ;
 wire \u_cpu.REG_FILE._02014_ ;
 wire \u_cpu.REG_FILE._02015_ ;
 wire \u_cpu.REG_FILE._02016_ ;
 wire \u_cpu.REG_FILE._02017_ ;
 wire \u_cpu.REG_FILE._02018_ ;
 wire \u_cpu.REG_FILE._02019_ ;
 wire \u_cpu.REG_FILE._02020_ ;
 wire \u_cpu.REG_FILE._02021_ ;
 wire \u_cpu.REG_FILE._02022_ ;
 wire \u_cpu.REG_FILE._02023_ ;
 wire \u_cpu.REG_FILE._02024_ ;
 wire \u_cpu.REG_FILE._02025_ ;
 wire \u_cpu.REG_FILE._02026_ ;
 wire \u_cpu.REG_FILE._02027_ ;
 wire \u_cpu.REG_FILE._02028_ ;
 wire \u_cpu.REG_FILE._02029_ ;
 wire \u_cpu.REG_FILE._02030_ ;
 wire \u_cpu.REG_FILE._02031_ ;
 wire \u_cpu.REG_FILE._02032_ ;
 wire \u_cpu.REG_FILE._02033_ ;
 wire \u_cpu.REG_FILE._02034_ ;
 wire \u_cpu.REG_FILE._02035_ ;
 wire \u_cpu.REG_FILE._02036_ ;
 wire \u_cpu.REG_FILE._02037_ ;
 wire \u_cpu.REG_FILE._02038_ ;
 wire \u_cpu.REG_FILE._02039_ ;
 wire \u_cpu.REG_FILE._02040_ ;
 wire \u_cpu.REG_FILE._02041_ ;
 wire \u_cpu.REG_FILE._02042_ ;
 wire \u_cpu.REG_FILE._02043_ ;
 wire \u_cpu.REG_FILE._02044_ ;
 wire \u_cpu.REG_FILE._02045_ ;
 wire \u_cpu.REG_FILE._02046_ ;
 wire \u_cpu.REG_FILE._02047_ ;
 wire \u_cpu.REG_FILE._02048_ ;
 wire \u_cpu.REG_FILE._02049_ ;
 wire \u_cpu.REG_FILE._02050_ ;
 wire \u_cpu.REG_FILE._02051_ ;
 wire \u_cpu.REG_FILE._02052_ ;
 wire \u_cpu.REG_FILE._02053_ ;
 wire \u_cpu.REG_FILE._02054_ ;
 wire \u_cpu.REG_FILE._02055_ ;
 wire \u_cpu.REG_FILE._02056_ ;
 wire \u_cpu.REG_FILE._02057_ ;
 wire \u_cpu.REG_FILE._02058_ ;
 wire \u_cpu.REG_FILE._02059_ ;
 wire \u_cpu.REG_FILE._02060_ ;
 wire \u_cpu.REG_FILE._02061_ ;
 wire \u_cpu.REG_FILE._02062_ ;
 wire \u_cpu.REG_FILE._02063_ ;
 wire \u_cpu.REG_FILE._02064_ ;
 wire \u_cpu.REG_FILE._02065_ ;
 wire \u_cpu.REG_FILE._02066_ ;
 wire \u_cpu.REG_FILE._02067_ ;
 wire \u_cpu.REG_FILE._02068_ ;
 wire \u_cpu.REG_FILE._02069_ ;
 wire \u_cpu.REG_FILE._02070_ ;
 wire \u_cpu.REG_FILE._02071_ ;
 wire \u_cpu.REG_FILE._02072_ ;
 wire \u_cpu.REG_FILE._02073_ ;
 wire \u_cpu.REG_FILE._02074_ ;
 wire \u_cpu.REG_FILE._02075_ ;
 wire \u_cpu.REG_FILE._02076_ ;
 wire \u_cpu.REG_FILE._02077_ ;
 wire \u_cpu.REG_FILE._02078_ ;
 wire \u_cpu.REG_FILE._02079_ ;
 wire \u_cpu.REG_FILE._02080_ ;
 wire \u_cpu.REG_FILE._02081_ ;
 wire \u_cpu.REG_FILE._02082_ ;
 wire \u_cpu.REG_FILE._02083_ ;
 wire \u_cpu.REG_FILE._02084_ ;
 wire \u_cpu.REG_FILE._02085_ ;
 wire \u_cpu.REG_FILE._02086_ ;
 wire \u_cpu.REG_FILE._02087_ ;
 wire \u_cpu.REG_FILE._02088_ ;
 wire \u_cpu.REG_FILE._02089_ ;
 wire \u_cpu.REG_FILE._02090_ ;
 wire \u_cpu.REG_FILE._02091_ ;
 wire \u_cpu.REG_FILE._02092_ ;
 wire \u_cpu.REG_FILE._02093_ ;
 wire \u_cpu.REG_FILE._02094_ ;
 wire \u_cpu.REG_FILE._02095_ ;
 wire \u_cpu.REG_FILE._02096_ ;
 wire \u_cpu.REG_FILE._02097_ ;
 wire \u_cpu.REG_FILE._02098_ ;
 wire \u_cpu.REG_FILE._02099_ ;
 wire \u_cpu.REG_FILE._02100_ ;
 wire \u_cpu.REG_FILE._02101_ ;
 wire \u_cpu.REG_FILE._02102_ ;
 wire \u_cpu.REG_FILE._02103_ ;
 wire \u_cpu.REG_FILE._02104_ ;
 wire \u_cpu.REG_FILE._02105_ ;
 wire \u_cpu.REG_FILE._02106_ ;
 wire \u_cpu.REG_FILE._02107_ ;
 wire \u_cpu.REG_FILE._02108_ ;
 wire \u_cpu.REG_FILE._02109_ ;
 wire \u_cpu.REG_FILE._02110_ ;
 wire \u_cpu.REG_FILE._02111_ ;
 wire \u_cpu.REG_FILE._02112_ ;
 wire \u_cpu.REG_FILE._02113_ ;
 wire \u_cpu.REG_FILE._02114_ ;
 wire \u_cpu.REG_FILE._02115_ ;
 wire \u_cpu.REG_FILE._02116_ ;
 wire \u_cpu.REG_FILE._02117_ ;
 wire \u_cpu.REG_FILE._02118_ ;
 wire \u_cpu.REG_FILE._02119_ ;
 wire \u_cpu.REG_FILE._02120_ ;
 wire \u_cpu.REG_FILE._02121_ ;
 wire \u_cpu.REG_FILE._02122_ ;
 wire \u_cpu.REG_FILE._02123_ ;
 wire \u_cpu.REG_FILE._02124_ ;
 wire \u_cpu.REG_FILE._02125_ ;
 wire \u_cpu.REG_FILE._02126_ ;
 wire \u_cpu.REG_FILE._02127_ ;
 wire \u_cpu.REG_FILE._02128_ ;
 wire \u_cpu.REG_FILE._02129_ ;
 wire \u_cpu.REG_FILE._02130_ ;
 wire \u_cpu.REG_FILE._02131_ ;
 wire \u_cpu.REG_FILE._02132_ ;
 wire \u_cpu.REG_FILE._02133_ ;
 wire \u_cpu.REG_FILE._02134_ ;
 wire \u_cpu.REG_FILE._02135_ ;
 wire \u_cpu.REG_FILE._02136_ ;
 wire \u_cpu.REG_FILE._02137_ ;
 wire \u_cpu.REG_FILE._02138_ ;
 wire \u_cpu.REG_FILE._02139_ ;
 wire \u_cpu.REG_FILE._02140_ ;
 wire \u_cpu.REG_FILE._02141_ ;
 wire \u_cpu.REG_FILE._02142_ ;
 wire \u_cpu.REG_FILE._02143_ ;
 wire \u_cpu.REG_FILE._02144_ ;
 wire \u_cpu.REG_FILE._02145_ ;
 wire \u_cpu.REG_FILE._02146_ ;
 wire \u_cpu.REG_FILE._02147_ ;
 wire \u_cpu.REG_FILE._02148_ ;
 wire \u_cpu.REG_FILE._02149_ ;
 wire \u_cpu.REG_FILE._02150_ ;
 wire \u_cpu.REG_FILE._02151_ ;
 wire \u_cpu.REG_FILE._02152_ ;
 wire \u_cpu.REG_FILE._02153_ ;
 wire \u_cpu.REG_FILE._02154_ ;
 wire \u_cpu.REG_FILE._02155_ ;
 wire \u_cpu.REG_FILE._02156_ ;
 wire \u_cpu.REG_FILE._02157_ ;
 wire \u_cpu.REG_FILE._02158_ ;
 wire \u_cpu.REG_FILE._02159_ ;
 wire \u_cpu.REG_FILE._02160_ ;
 wire \u_cpu.REG_FILE._02161_ ;
 wire \u_cpu.REG_FILE._02162_ ;
 wire \u_cpu.REG_FILE._02163_ ;
 wire \u_cpu.REG_FILE._02164_ ;
 wire \u_cpu.REG_FILE._02165_ ;
 wire \u_cpu.REG_FILE._02166_ ;
 wire \u_cpu.REG_FILE._02167_ ;
 wire \u_cpu.REG_FILE._02168_ ;
 wire \u_cpu.REG_FILE._02169_ ;
 wire \u_cpu.REG_FILE._02170_ ;
 wire \u_cpu.REG_FILE._02171_ ;
 wire \u_cpu.REG_FILE._02172_ ;
 wire \u_cpu.REG_FILE._02173_ ;
 wire \u_cpu.REG_FILE._02174_ ;
 wire \u_cpu.REG_FILE._02175_ ;
 wire \u_cpu.REG_FILE._02176_ ;
 wire \u_cpu.REG_FILE._02177_ ;
 wire \u_cpu.REG_FILE._02178_ ;
 wire \u_cpu.REG_FILE._02179_ ;
 wire \u_cpu.REG_FILE._02180_ ;
 wire \u_cpu.REG_FILE._02181_ ;
 wire \u_cpu.REG_FILE._02182_ ;
 wire \u_cpu.REG_FILE._02183_ ;
 wire \u_cpu.REG_FILE._02184_ ;
 wire \u_cpu.REG_FILE._02185_ ;
 wire \u_cpu.REG_FILE._02186_ ;
 wire \u_cpu.REG_FILE._02187_ ;
 wire \u_cpu.REG_FILE._02188_ ;
 wire \u_cpu.REG_FILE._02189_ ;
 wire \u_cpu.REG_FILE._02190_ ;
 wire \u_cpu.REG_FILE._02191_ ;
 wire \u_cpu.REG_FILE._02192_ ;
 wire \u_cpu.REG_FILE._02193_ ;
 wire \u_cpu.REG_FILE._02194_ ;
 wire \u_cpu.REG_FILE._02195_ ;
 wire \u_cpu.REG_FILE._02196_ ;
 wire \u_cpu.REG_FILE._02197_ ;
 wire \u_cpu.REG_FILE._02198_ ;
 wire \u_cpu.REG_FILE._02199_ ;
 wire \u_cpu.REG_FILE._02200_ ;
 wire \u_cpu.REG_FILE._02201_ ;
 wire \u_cpu.REG_FILE._02202_ ;
 wire \u_cpu.REG_FILE._02203_ ;
 wire \u_cpu.REG_FILE._02204_ ;
 wire \u_cpu.REG_FILE._02205_ ;
 wire \u_cpu.REG_FILE._02206_ ;
 wire \u_cpu.REG_FILE._02207_ ;
 wire \u_cpu.REG_FILE._02208_ ;
 wire \u_cpu.REG_FILE._02209_ ;
 wire \u_cpu.REG_FILE._02210_ ;
 wire \u_cpu.REG_FILE._02211_ ;
 wire \u_cpu.REG_FILE._02212_ ;
 wire \u_cpu.REG_FILE._02213_ ;
 wire \u_cpu.REG_FILE._02214_ ;
 wire \u_cpu.REG_FILE._02215_ ;
 wire \u_cpu.REG_FILE._02216_ ;
 wire \u_cpu.REG_FILE._02217_ ;
 wire \u_cpu.REG_FILE._02218_ ;
 wire \u_cpu.REG_FILE._02219_ ;
 wire \u_cpu.REG_FILE._02220_ ;
 wire \u_cpu.REG_FILE._02221_ ;
 wire \u_cpu.REG_FILE._02222_ ;
 wire \u_cpu.REG_FILE._02223_ ;
 wire \u_cpu.REG_FILE._02224_ ;
 wire \u_cpu.REG_FILE._02225_ ;
 wire \u_cpu.REG_FILE._02226_ ;
 wire \u_cpu.REG_FILE._02227_ ;
 wire \u_cpu.REG_FILE._02228_ ;
 wire \u_cpu.REG_FILE._02229_ ;
 wire \u_cpu.REG_FILE._02230_ ;
 wire \u_cpu.REG_FILE._02231_ ;
 wire \u_cpu.REG_FILE._02232_ ;
 wire \u_cpu.REG_FILE._02233_ ;
 wire \u_cpu.REG_FILE._02234_ ;
 wire \u_cpu.REG_FILE._02235_ ;
 wire \u_cpu.REG_FILE._02236_ ;
 wire \u_cpu.REG_FILE._02237_ ;
 wire \u_cpu.REG_FILE._02238_ ;
 wire \u_cpu.REG_FILE._02239_ ;
 wire \u_cpu.REG_FILE._02240_ ;
 wire \u_cpu.REG_FILE._02241_ ;
 wire \u_cpu.REG_FILE._02242_ ;
 wire \u_cpu.REG_FILE._02243_ ;
 wire \u_cpu.REG_FILE._02244_ ;
 wire \u_cpu.REG_FILE._02245_ ;
 wire \u_cpu.REG_FILE._02246_ ;
 wire \u_cpu.REG_FILE._02247_ ;
 wire \u_cpu.REG_FILE._02248_ ;
 wire \u_cpu.REG_FILE._02249_ ;
 wire \u_cpu.REG_FILE._02250_ ;
 wire \u_cpu.REG_FILE._02251_ ;
 wire \u_cpu.REG_FILE._02252_ ;
 wire \u_cpu.REG_FILE._02253_ ;
 wire \u_cpu.REG_FILE._02254_ ;
 wire \u_cpu.REG_FILE._02255_ ;
 wire \u_cpu.REG_FILE._02256_ ;
 wire \u_cpu.REG_FILE._02257_ ;
 wire \u_cpu.REG_FILE._02258_ ;
 wire \u_cpu.REG_FILE._02259_ ;
 wire \u_cpu.REG_FILE._02260_ ;
 wire \u_cpu.REG_FILE._02261_ ;
 wire \u_cpu.REG_FILE._02262_ ;
 wire \u_cpu.REG_FILE._02263_ ;
 wire \u_cpu.REG_FILE._02264_ ;
 wire \u_cpu.REG_FILE._02265_ ;
 wire \u_cpu.REG_FILE._02266_ ;
 wire \u_cpu.REG_FILE._02267_ ;
 wire \u_cpu.REG_FILE._02268_ ;
 wire \u_cpu.REG_FILE._02269_ ;
 wire \u_cpu.REG_FILE._02270_ ;
 wire \u_cpu.REG_FILE._02271_ ;
 wire \u_cpu.REG_FILE._02272_ ;
 wire \u_cpu.REG_FILE._02273_ ;
 wire \u_cpu.REG_FILE._02274_ ;
 wire \u_cpu.REG_FILE._02275_ ;
 wire \u_cpu.REG_FILE._02276_ ;
 wire \u_cpu.REG_FILE._02277_ ;
 wire \u_cpu.REG_FILE._02278_ ;
 wire \u_cpu.REG_FILE._02279_ ;
 wire \u_cpu.REG_FILE._02280_ ;
 wire \u_cpu.REG_FILE._02281_ ;
 wire \u_cpu.REG_FILE._02282_ ;
 wire \u_cpu.REG_FILE._02283_ ;
 wire \u_cpu.REG_FILE._02284_ ;
 wire \u_cpu.REG_FILE._02285_ ;
 wire \u_cpu.REG_FILE._02286_ ;
 wire \u_cpu.REG_FILE._02287_ ;
 wire \u_cpu.REG_FILE._02288_ ;
 wire \u_cpu.REG_FILE._02289_ ;
 wire \u_cpu.REG_FILE._02290_ ;
 wire \u_cpu.REG_FILE._02291_ ;
 wire \u_cpu.REG_FILE._02292_ ;
 wire \u_cpu.REG_FILE._02293_ ;
 wire \u_cpu.REG_FILE._02294_ ;
 wire \u_cpu.REG_FILE._02295_ ;
 wire \u_cpu.REG_FILE._02296_ ;
 wire \u_cpu.REG_FILE._02297_ ;
 wire \u_cpu.REG_FILE._02298_ ;
 wire \u_cpu.REG_FILE._02299_ ;
 wire \u_cpu.REG_FILE._02300_ ;
 wire \u_cpu.REG_FILE._02301_ ;
 wire \u_cpu.REG_FILE._02302_ ;
 wire \u_cpu.REG_FILE._02303_ ;
 wire \u_cpu.REG_FILE._02304_ ;
 wire \u_cpu.REG_FILE._02305_ ;
 wire \u_cpu.REG_FILE._02306_ ;
 wire \u_cpu.REG_FILE._02307_ ;
 wire \u_cpu.REG_FILE._02308_ ;
 wire \u_cpu.REG_FILE._02309_ ;
 wire \u_cpu.REG_FILE._02310_ ;
 wire \u_cpu.REG_FILE._02311_ ;
 wire \u_cpu.REG_FILE._02312_ ;
 wire \u_cpu.REG_FILE._02313_ ;
 wire \u_cpu.REG_FILE._02314_ ;
 wire \u_cpu.REG_FILE._02315_ ;
 wire \u_cpu.REG_FILE._02316_ ;
 wire \u_cpu.REG_FILE._02317_ ;
 wire \u_cpu.REG_FILE._02318_ ;
 wire \u_cpu.REG_FILE._02319_ ;
 wire \u_cpu.REG_FILE._02320_ ;
 wire \u_cpu.REG_FILE._02321_ ;
 wire \u_cpu.REG_FILE._02322_ ;
 wire \u_cpu.REG_FILE._02323_ ;
 wire \u_cpu.REG_FILE._02324_ ;
 wire \u_cpu.REG_FILE._02325_ ;
 wire \u_cpu.REG_FILE._02326_ ;
 wire \u_cpu.REG_FILE._02327_ ;
 wire \u_cpu.REG_FILE._02328_ ;
 wire \u_cpu.REG_FILE._02329_ ;
 wire \u_cpu.REG_FILE._02330_ ;
 wire \u_cpu.REG_FILE._02331_ ;
 wire \u_cpu.REG_FILE._02332_ ;
 wire \u_cpu.REG_FILE._02333_ ;
 wire \u_cpu.REG_FILE._02334_ ;
 wire \u_cpu.REG_FILE._02335_ ;
 wire \u_cpu.REG_FILE._02336_ ;
 wire \u_cpu.REG_FILE._02337_ ;
 wire \u_cpu.REG_FILE._02338_ ;
 wire \u_cpu.REG_FILE._02339_ ;
 wire \u_cpu.REG_FILE._02340_ ;
 wire \u_cpu.REG_FILE._02341_ ;
 wire \u_cpu.REG_FILE._02342_ ;
 wire \u_cpu.REG_FILE._02343_ ;
 wire \u_cpu.REG_FILE._02344_ ;
 wire \u_cpu.REG_FILE._02345_ ;
 wire \u_cpu.REG_FILE._02346_ ;
 wire \u_cpu.REG_FILE._02347_ ;
 wire \u_cpu.REG_FILE._02348_ ;
 wire \u_cpu.REG_FILE._02349_ ;
 wire \u_cpu.REG_FILE._02350_ ;
 wire \u_cpu.REG_FILE._02351_ ;
 wire \u_cpu.REG_FILE._02352_ ;
 wire \u_cpu.REG_FILE._02353_ ;
 wire \u_cpu.REG_FILE._02354_ ;
 wire \u_cpu.REG_FILE._02355_ ;
 wire \u_cpu.REG_FILE._02356_ ;
 wire \u_cpu.REG_FILE._02357_ ;
 wire \u_cpu.REG_FILE._02358_ ;
 wire \u_cpu.REG_FILE._02359_ ;
 wire \u_cpu.REG_FILE._02360_ ;
 wire \u_cpu.REG_FILE._02361_ ;
 wire \u_cpu.REG_FILE._02362_ ;
 wire \u_cpu.REG_FILE._02363_ ;
 wire \u_cpu.REG_FILE._02364_ ;
 wire \u_cpu.REG_FILE._02365_ ;
 wire \u_cpu.REG_FILE._02366_ ;
 wire \u_cpu.REG_FILE._02367_ ;
 wire \u_cpu.REG_FILE._02368_ ;
 wire \u_cpu.REG_FILE._02369_ ;
 wire \u_cpu.REG_FILE._02370_ ;
 wire \u_cpu.REG_FILE._02371_ ;
 wire \u_cpu.REG_FILE._02372_ ;
 wire \u_cpu.REG_FILE._02373_ ;
 wire \u_cpu.REG_FILE._02374_ ;
 wire \u_cpu.REG_FILE._02375_ ;
 wire \u_cpu.REG_FILE._02376_ ;
 wire \u_cpu.REG_FILE._02377_ ;
 wire \u_cpu.REG_FILE._02378_ ;
 wire \u_cpu.REG_FILE._02379_ ;
 wire \u_cpu.REG_FILE._02380_ ;
 wire \u_cpu.REG_FILE._02381_ ;
 wire \u_cpu.REG_FILE._02382_ ;
 wire \u_cpu.REG_FILE._02383_ ;
 wire \u_cpu.REG_FILE._02384_ ;
 wire \u_cpu.REG_FILE._02385_ ;
 wire \u_cpu.REG_FILE._02386_ ;
 wire \u_cpu.REG_FILE._02387_ ;
 wire \u_cpu.REG_FILE._02388_ ;
 wire \u_cpu.REG_FILE._02389_ ;
 wire \u_cpu.REG_FILE._02390_ ;
 wire \u_cpu.REG_FILE._02391_ ;
 wire \u_cpu.REG_FILE._02392_ ;
 wire \u_cpu.REG_FILE._02393_ ;
 wire \u_cpu.REG_FILE._02394_ ;
 wire \u_cpu.REG_FILE._02395_ ;
 wire \u_cpu.REG_FILE._02396_ ;
 wire \u_cpu.REG_FILE._02397_ ;
 wire \u_cpu.REG_FILE._02398_ ;
 wire \u_cpu.REG_FILE._02399_ ;
 wire \u_cpu.REG_FILE._02400_ ;
 wire \u_cpu.REG_FILE._02401_ ;
 wire \u_cpu.REG_FILE._02402_ ;
 wire \u_cpu.REG_FILE._02403_ ;
 wire \u_cpu.REG_FILE._02404_ ;
 wire \u_cpu.REG_FILE._02405_ ;
 wire \u_cpu.REG_FILE._02406_ ;
 wire \u_cpu.REG_FILE._02407_ ;
 wire \u_cpu.REG_FILE._02408_ ;
 wire \u_cpu.REG_FILE._02409_ ;
 wire \u_cpu.REG_FILE._02410_ ;
 wire \u_cpu.REG_FILE._02411_ ;
 wire \u_cpu.REG_FILE._02412_ ;
 wire \u_cpu.REG_FILE._02413_ ;
 wire \u_cpu.REG_FILE._02414_ ;
 wire \u_cpu.REG_FILE._02415_ ;
 wire \u_cpu.REG_FILE._02416_ ;
 wire \u_cpu.REG_FILE._02417_ ;
 wire \u_cpu.REG_FILE._02418_ ;
 wire \u_cpu.REG_FILE._02419_ ;
 wire \u_cpu.REG_FILE._02420_ ;
 wire \u_cpu.REG_FILE._02421_ ;
 wire \u_cpu.REG_FILE._02422_ ;
 wire \u_cpu.REG_FILE._02423_ ;
 wire \u_cpu.REG_FILE._02424_ ;
 wire \u_cpu.REG_FILE._02425_ ;
 wire \u_cpu.REG_FILE._02426_ ;
 wire \u_cpu.REG_FILE._02427_ ;
 wire \u_cpu.REG_FILE._02428_ ;
 wire \u_cpu.REG_FILE._02429_ ;
 wire \u_cpu.REG_FILE._02430_ ;
 wire \u_cpu.REG_FILE._02431_ ;
 wire \u_cpu.REG_FILE._02432_ ;
 wire \u_cpu.REG_FILE._02433_ ;
 wire \u_cpu.REG_FILE._02434_ ;
 wire \u_cpu.REG_FILE._02435_ ;
 wire \u_cpu.REG_FILE._02436_ ;
 wire \u_cpu.REG_FILE._02437_ ;
 wire \u_cpu.REG_FILE._02438_ ;
 wire \u_cpu.REG_FILE._02439_ ;
 wire \u_cpu.REG_FILE._02440_ ;
 wire \u_cpu.REG_FILE._02441_ ;
 wire \u_cpu.REG_FILE._02442_ ;
 wire \u_cpu.REG_FILE._02443_ ;
 wire \u_cpu.REG_FILE._02444_ ;
 wire \u_cpu.REG_FILE._02445_ ;
 wire \u_cpu.REG_FILE._02446_ ;
 wire \u_cpu.REG_FILE._02447_ ;
 wire \u_cpu.REG_FILE._02448_ ;
 wire \u_cpu.REG_FILE._02449_ ;
 wire \u_cpu.REG_FILE._02450_ ;
 wire \u_cpu.REG_FILE._02451_ ;
 wire \u_cpu.REG_FILE._02452_ ;
 wire \u_cpu.REG_FILE._02453_ ;
 wire \u_cpu.REG_FILE._02454_ ;
 wire \u_cpu.REG_FILE._02455_ ;
 wire \u_cpu.REG_FILE._02456_ ;
 wire \u_cpu.REG_FILE._02457_ ;
 wire \u_cpu.REG_FILE._02458_ ;
 wire \u_cpu.REG_FILE._02459_ ;
 wire \u_cpu.REG_FILE._02460_ ;
 wire \u_cpu.REG_FILE._02461_ ;
 wire \u_cpu.REG_FILE._02462_ ;
 wire \u_cpu.REG_FILE._02463_ ;
 wire \u_cpu.REG_FILE._02464_ ;
 wire \u_cpu.REG_FILE._02465_ ;
 wire \u_cpu.REG_FILE._02466_ ;
 wire \u_cpu.REG_FILE._02467_ ;
 wire \u_cpu.REG_FILE._02468_ ;
 wire \u_cpu.REG_FILE._02469_ ;
 wire \u_cpu.REG_FILE._02470_ ;
 wire \u_cpu.REG_FILE._02471_ ;
 wire \u_cpu.REG_FILE._02472_ ;
 wire \u_cpu.REG_FILE._02473_ ;
 wire \u_cpu.REG_FILE._02474_ ;
 wire \u_cpu.REG_FILE._02475_ ;
 wire \u_cpu.REG_FILE._02476_ ;
 wire \u_cpu.REG_FILE._02477_ ;
 wire \u_cpu.REG_FILE._02478_ ;
 wire \u_cpu.REG_FILE._02479_ ;
 wire \u_cpu.REG_FILE._02480_ ;
 wire \u_cpu.REG_FILE._02481_ ;
 wire \u_cpu.REG_FILE._02482_ ;
 wire \u_cpu.REG_FILE._02483_ ;
 wire \u_cpu.REG_FILE._02484_ ;
 wire \u_cpu.REG_FILE._02485_ ;
 wire \u_cpu.REG_FILE._02486_ ;
 wire \u_cpu.REG_FILE._02487_ ;
 wire \u_cpu.REG_FILE._02488_ ;
 wire \u_cpu.REG_FILE._02489_ ;
 wire \u_cpu.REG_FILE._02490_ ;
 wire \u_cpu.REG_FILE._02491_ ;
 wire \u_cpu.REG_FILE._02492_ ;
 wire \u_cpu.REG_FILE._02493_ ;
 wire \u_cpu.REG_FILE._02494_ ;
 wire \u_cpu.REG_FILE._02495_ ;
 wire \u_cpu.REG_FILE._02496_ ;
 wire \u_cpu.REG_FILE._02497_ ;
 wire \u_cpu.REG_FILE._02498_ ;
 wire \u_cpu.REG_FILE._02499_ ;
 wire \u_cpu.REG_FILE._02500_ ;
 wire \u_cpu.REG_FILE._02501_ ;
 wire \u_cpu.REG_FILE._02502_ ;
 wire \u_cpu.REG_FILE._02503_ ;
 wire \u_cpu.REG_FILE._02504_ ;
 wire \u_cpu.REG_FILE._02505_ ;
 wire \u_cpu.REG_FILE._02506_ ;
 wire \u_cpu.REG_FILE._02507_ ;
 wire \u_cpu.REG_FILE._02508_ ;
 wire \u_cpu.REG_FILE._02509_ ;
 wire \u_cpu.REG_FILE._02510_ ;
 wire \u_cpu.REG_FILE._02511_ ;
 wire \u_cpu.REG_FILE._02512_ ;
 wire \u_cpu.REG_FILE._02513_ ;
 wire \u_cpu.REG_FILE._02514_ ;
 wire \u_cpu.REG_FILE._02515_ ;
 wire \u_cpu.REG_FILE._02516_ ;
 wire \u_cpu.REG_FILE._02517_ ;
 wire \u_cpu.REG_FILE._02518_ ;
 wire \u_cpu.REG_FILE._02519_ ;
 wire \u_cpu.REG_FILE._02520_ ;
 wire \u_cpu.REG_FILE._02521_ ;
 wire \u_cpu.REG_FILE._02522_ ;
 wire \u_cpu.REG_FILE._02523_ ;
 wire \u_cpu.REG_FILE._02524_ ;
 wire \u_cpu.REG_FILE._02525_ ;
 wire \u_cpu.REG_FILE._02526_ ;
 wire \u_cpu.REG_FILE._02527_ ;
 wire \u_cpu.REG_FILE._02528_ ;
 wire \u_cpu.REG_FILE._02529_ ;
 wire \u_cpu.REG_FILE._02530_ ;
 wire \u_cpu.REG_FILE._02531_ ;
 wire \u_cpu.REG_FILE._02532_ ;
 wire \u_cpu.REG_FILE._02533_ ;
 wire \u_cpu.REG_FILE._02534_ ;
 wire \u_cpu.REG_FILE._02535_ ;
 wire \u_cpu.REG_FILE._02536_ ;
 wire \u_cpu.REG_FILE._02537_ ;
 wire \u_cpu.REG_FILE._02538_ ;
 wire \u_cpu.REG_FILE._02539_ ;
 wire \u_cpu.REG_FILE._02540_ ;
 wire \u_cpu.REG_FILE._02541_ ;
 wire \u_cpu.REG_FILE._02542_ ;
 wire \u_cpu.REG_FILE._02543_ ;
 wire \u_cpu.REG_FILE._02544_ ;
 wire \u_cpu.REG_FILE._02545_ ;
 wire \u_cpu.REG_FILE._02546_ ;
 wire \u_cpu.REG_FILE._02547_ ;
 wire \u_cpu.REG_FILE._02548_ ;
 wire \u_cpu.REG_FILE._02549_ ;
 wire \u_cpu.REG_FILE._02550_ ;
 wire \u_cpu.REG_FILE._02551_ ;
 wire \u_cpu.REG_FILE._02552_ ;
 wire \u_cpu.REG_FILE._02553_ ;
 wire \u_cpu.REG_FILE._02554_ ;
 wire \u_cpu.REG_FILE._02555_ ;
 wire \u_cpu.REG_FILE._02556_ ;
 wire \u_cpu.REG_FILE._02557_ ;
 wire \u_cpu.REG_FILE._02558_ ;
 wire \u_cpu.REG_FILE._02559_ ;
 wire \u_cpu.REG_FILE._02560_ ;
 wire \u_cpu.REG_FILE._02561_ ;
 wire \u_cpu.REG_FILE._02562_ ;
 wire \u_cpu.REG_FILE._02563_ ;
 wire \u_cpu.REG_FILE._02564_ ;
 wire \u_cpu.REG_FILE._02565_ ;
 wire \u_cpu.REG_FILE._02566_ ;
 wire \u_cpu.REG_FILE._02567_ ;
 wire \u_cpu.REG_FILE._02568_ ;
 wire \u_cpu.REG_FILE._02569_ ;
 wire \u_cpu.REG_FILE._02570_ ;
 wire \u_cpu.REG_FILE._02571_ ;
 wire \u_cpu.REG_FILE._02572_ ;
 wire \u_cpu.REG_FILE._02573_ ;
 wire \u_cpu.REG_FILE._02574_ ;
 wire \u_cpu.REG_FILE._02575_ ;
 wire \u_cpu.REG_FILE._02576_ ;
 wire \u_cpu.REG_FILE._02577_ ;
 wire \u_cpu.REG_FILE._02578_ ;
 wire \u_cpu.REG_FILE._02579_ ;
 wire \u_cpu.REG_FILE._02580_ ;
 wire \u_cpu.REG_FILE._02581_ ;
 wire \u_cpu.REG_FILE._02582_ ;
 wire \u_cpu.REG_FILE._02583_ ;
 wire \u_cpu.REG_FILE._02584_ ;
 wire \u_cpu.REG_FILE._02585_ ;
 wire \u_cpu.REG_FILE._02586_ ;
 wire \u_cpu.REG_FILE._02587_ ;
 wire \u_cpu.REG_FILE._02588_ ;
 wire \u_cpu.REG_FILE._02589_ ;
 wire \u_cpu.REG_FILE._02590_ ;
 wire \u_cpu.REG_FILE._02591_ ;
 wire \u_cpu.REG_FILE._02592_ ;
 wire \u_cpu.REG_FILE._02593_ ;
 wire \u_cpu.REG_FILE._02594_ ;
 wire \u_cpu.REG_FILE._02595_ ;
 wire \u_cpu.REG_FILE._02596_ ;
 wire \u_cpu.REG_FILE._02597_ ;
 wire \u_cpu.REG_FILE._02598_ ;
 wire \u_cpu.REG_FILE._02599_ ;
 wire \u_cpu.REG_FILE._02600_ ;
 wire \u_cpu.REG_FILE._02601_ ;
 wire \u_cpu.REG_FILE._02602_ ;
 wire \u_cpu.REG_FILE._02603_ ;
 wire \u_cpu.REG_FILE._02604_ ;
 wire \u_cpu.REG_FILE._02605_ ;
 wire \u_cpu.REG_FILE._02606_ ;
 wire \u_cpu.REG_FILE._02607_ ;
 wire \u_cpu.REG_FILE._02608_ ;
 wire \u_cpu.REG_FILE._02609_ ;
 wire \u_cpu.REG_FILE._02610_ ;
 wire \u_cpu.REG_FILE._02611_ ;
 wire \u_cpu.REG_FILE._02612_ ;
 wire \u_cpu.REG_FILE._02613_ ;
 wire \u_cpu.REG_FILE._02614_ ;
 wire \u_cpu.REG_FILE._02615_ ;
 wire \u_cpu.REG_FILE._02616_ ;
 wire \u_cpu.REG_FILE._02617_ ;
 wire \u_cpu.REG_FILE._02618_ ;
 wire \u_cpu.REG_FILE._02619_ ;
 wire \u_cpu.REG_FILE._02620_ ;
 wire \u_cpu.REG_FILE._02621_ ;
 wire \u_cpu.REG_FILE._02622_ ;
 wire \u_cpu.REG_FILE._02623_ ;
 wire \u_cpu.REG_FILE._02624_ ;
 wire \u_cpu.REG_FILE._02625_ ;
 wire \u_cpu.REG_FILE._02626_ ;
 wire \u_cpu.REG_FILE._02627_ ;
 wire \u_cpu.REG_FILE._02628_ ;
 wire \u_cpu.REG_FILE._02629_ ;
 wire \u_cpu.REG_FILE._02630_ ;
 wire \u_cpu.REG_FILE._02631_ ;
 wire \u_cpu.REG_FILE._02632_ ;
 wire \u_cpu.REG_FILE._02633_ ;
 wire \u_cpu.REG_FILE._02634_ ;
 wire \u_cpu.REG_FILE._02635_ ;
 wire \u_cpu.REG_FILE._02636_ ;
 wire \u_cpu.REG_FILE._02637_ ;
 wire \u_cpu.REG_FILE._02638_ ;
 wire \u_cpu.REG_FILE._02639_ ;
 wire \u_cpu.REG_FILE._02640_ ;
 wire \u_cpu.REG_FILE._02641_ ;
 wire \u_cpu.REG_FILE._02642_ ;
 wire \u_cpu.REG_FILE._02643_ ;
 wire \u_cpu.REG_FILE._02644_ ;
 wire \u_cpu.REG_FILE._02645_ ;
 wire \u_cpu.REG_FILE._02646_ ;
 wire \u_cpu.REG_FILE._02647_ ;
 wire \u_cpu.REG_FILE._02648_ ;
 wire \u_cpu.REG_FILE._02649_ ;
 wire \u_cpu.REG_FILE._02650_ ;
 wire \u_cpu.REG_FILE._02651_ ;
 wire \u_cpu.REG_FILE._02652_ ;
 wire \u_cpu.REG_FILE._02653_ ;
 wire \u_cpu.REG_FILE._02654_ ;
 wire \u_cpu.REG_FILE._02655_ ;
 wire \u_cpu.REG_FILE._02656_ ;
 wire \u_cpu.REG_FILE._02657_ ;
 wire \u_cpu.REG_FILE._02658_ ;
 wire \u_cpu.REG_FILE._02659_ ;
 wire \u_cpu.REG_FILE._02660_ ;
 wire \u_cpu.REG_FILE._02661_ ;
 wire \u_cpu.REG_FILE._02662_ ;
 wire \u_cpu.REG_FILE._02663_ ;
 wire \u_cpu.REG_FILE._02664_ ;
 wire \u_cpu.REG_FILE._02665_ ;
 wire \u_cpu.REG_FILE._02666_ ;
 wire \u_cpu.REG_FILE._02667_ ;
 wire \u_cpu.REG_FILE._02668_ ;
 wire \u_cpu.REG_FILE._02669_ ;
 wire \u_cpu.REG_FILE._02670_ ;
 wire \u_cpu.REG_FILE._02671_ ;
 wire \u_cpu.REG_FILE._02672_ ;
 wire \u_cpu.REG_FILE._02673_ ;
 wire \u_cpu.REG_FILE._02674_ ;
 wire \u_cpu.REG_FILE._02675_ ;
 wire \u_cpu.REG_FILE._02676_ ;
 wire \u_cpu.REG_FILE._02677_ ;
 wire \u_cpu.REG_FILE._02678_ ;
 wire \u_cpu.REG_FILE._02679_ ;
 wire \u_cpu.REG_FILE._02680_ ;
 wire \u_cpu.REG_FILE._02681_ ;
 wire \u_cpu.REG_FILE._02682_ ;
 wire \u_cpu.REG_FILE._02683_ ;
 wire \u_cpu.REG_FILE._02684_ ;
 wire \u_cpu.REG_FILE._02685_ ;
 wire \u_cpu.REG_FILE._02686_ ;
 wire \u_cpu.REG_FILE._02687_ ;
 wire \u_cpu.REG_FILE._02688_ ;
 wire \u_cpu.REG_FILE._02689_ ;
 wire \u_cpu.REG_FILE._02690_ ;
 wire \u_cpu.REG_FILE._02691_ ;
 wire \u_cpu.REG_FILE._02692_ ;
 wire \u_cpu.REG_FILE._02693_ ;
 wire \u_cpu.REG_FILE._02694_ ;
 wire \u_cpu.REG_FILE._02695_ ;
 wire \u_cpu.REG_FILE._02696_ ;
 wire \u_cpu.REG_FILE._02697_ ;
 wire \u_cpu.REG_FILE._02698_ ;
 wire \u_cpu.REG_FILE._02699_ ;
 wire \u_cpu.REG_FILE._02700_ ;
 wire \u_cpu.REG_FILE._02701_ ;
 wire \u_cpu.REG_FILE._02702_ ;
 wire \u_cpu.REG_FILE._02703_ ;
 wire \u_cpu.REG_FILE._02704_ ;
 wire \u_cpu.REG_FILE._02705_ ;
 wire \u_cpu.REG_FILE._02706_ ;
 wire \u_cpu.REG_FILE._02707_ ;
 wire \u_cpu.REG_FILE._02708_ ;
 wire \u_cpu.REG_FILE._02709_ ;
 wire \u_cpu.REG_FILE._02710_ ;
 wire \u_cpu.REG_FILE._02711_ ;
 wire \u_cpu.REG_FILE._02712_ ;
 wire \u_cpu.REG_FILE._02713_ ;
 wire \u_cpu.REG_FILE._02714_ ;
 wire \u_cpu.REG_FILE._02715_ ;
 wire \u_cpu.REG_FILE._02716_ ;
 wire \u_cpu.REG_FILE._02717_ ;
 wire \u_cpu.REG_FILE._02718_ ;
 wire \u_cpu.REG_FILE._02719_ ;
 wire \u_cpu.REG_FILE._02720_ ;
 wire \u_cpu.REG_FILE._02721_ ;
 wire \u_cpu.REG_FILE._02722_ ;
 wire \u_cpu.REG_FILE._02723_ ;
 wire \u_cpu.REG_FILE._02724_ ;
 wire \u_cpu.REG_FILE._02725_ ;
 wire \u_cpu.REG_FILE._02726_ ;
 wire \u_cpu.REG_FILE._02727_ ;
 wire \u_cpu.REG_FILE._02728_ ;
 wire \u_cpu.REG_FILE._02729_ ;
 wire \u_cpu.REG_FILE._02730_ ;
 wire \u_cpu.REG_FILE._02731_ ;
 wire \u_cpu.REG_FILE._02732_ ;
 wire \u_cpu.REG_FILE._02733_ ;
 wire \u_cpu.REG_FILE._02734_ ;
 wire \u_cpu.REG_FILE._02735_ ;
 wire \u_cpu.REG_FILE._02736_ ;
 wire \u_cpu.REG_FILE._02737_ ;
 wire \u_cpu.REG_FILE._02738_ ;
 wire \u_cpu.REG_FILE._02739_ ;
 wire \u_cpu.REG_FILE._02740_ ;
 wire \u_cpu.REG_FILE._02741_ ;
 wire \u_cpu.REG_FILE._02742_ ;
 wire \u_cpu.REG_FILE._02743_ ;
 wire \u_cpu.REG_FILE._02744_ ;
 wire \u_cpu.REG_FILE._02745_ ;
 wire \u_cpu.REG_FILE._02746_ ;
 wire \u_cpu.REG_FILE._02747_ ;
 wire \u_cpu.REG_FILE._02748_ ;
 wire \u_cpu.REG_FILE._02749_ ;
 wire \u_cpu.REG_FILE._02750_ ;
 wire \u_cpu.REG_FILE._02751_ ;
 wire \u_cpu.REG_FILE._02752_ ;
 wire \u_cpu.REG_FILE._02753_ ;
 wire \u_cpu.REG_FILE._02754_ ;
 wire \u_cpu.REG_FILE._02755_ ;
 wire \u_cpu.REG_FILE._02756_ ;
 wire \u_cpu.REG_FILE._02757_ ;
 wire \u_cpu.REG_FILE._02758_ ;
 wire \u_cpu.REG_FILE._02759_ ;
 wire \u_cpu.REG_FILE._02760_ ;
 wire \u_cpu.REG_FILE._02761_ ;
 wire \u_cpu.REG_FILE._02762_ ;
 wire \u_cpu.REG_FILE._02763_ ;
 wire \u_cpu.REG_FILE._02764_ ;
 wire \u_cpu.REG_FILE._02765_ ;
 wire \u_cpu.REG_FILE._02766_ ;
 wire \u_cpu.REG_FILE._02767_ ;
 wire \u_cpu.REG_FILE._02768_ ;
 wire \u_cpu.REG_FILE._02769_ ;
 wire \u_cpu.REG_FILE._02770_ ;
 wire \u_cpu.REG_FILE._02771_ ;
 wire \u_cpu.REG_FILE._02772_ ;
 wire \u_cpu.REG_FILE._02773_ ;
 wire \u_cpu.REG_FILE._02774_ ;
 wire \u_cpu.REG_FILE._02775_ ;
 wire \u_cpu.REG_FILE._02776_ ;
 wire \u_cpu.REG_FILE._02777_ ;
 wire \u_cpu.REG_FILE._02778_ ;
 wire \u_cpu.REG_FILE._02779_ ;
 wire \u_cpu.REG_FILE._02780_ ;
 wire \u_cpu.REG_FILE._02781_ ;
 wire \u_cpu.REG_FILE._02782_ ;
 wire \u_cpu.REG_FILE._02783_ ;
 wire \u_cpu.REG_FILE._02784_ ;
 wire \u_cpu.REG_FILE._02785_ ;
 wire \u_cpu.REG_FILE._02786_ ;
 wire \u_cpu.REG_FILE._02787_ ;
 wire \u_cpu.REG_FILE._02788_ ;
 wire \u_cpu.REG_FILE._02789_ ;
 wire \u_cpu.REG_FILE._02790_ ;
 wire \u_cpu.REG_FILE._02791_ ;
 wire \u_cpu.REG_FILE._02792_ ;
 wire \u_cpu.REG_FILE._02793_ ;
 wire \u_cpu.REG_FILE._02794_ ;
 wire \u_cpu.REG_FILE._02795_ ;
 wire \u_cpu.REG_FILE._02796_ ;
 wire \u_cpu.REG_FILE._02797_ ;
 wire \u_cpu.REG_FILE._02798_ ;
 wire \u_cpu.REG_FILE._02799_ ;
 wire \u_cpu.REG_FILE._02800_ ;
 wire \u_cpu.REG_FILE._02801_ ;
 wire \u_cpu.REG_FILE._02802_ ;
 wire \u_cpu.REG_FILE._02803_ ;
 wire \u_cpu.REG_FILE._02804_ ;
 wire \u_cpu.REG_FILE._02805_ ;
 wire \u_cpu.REG_FILE._02806_ ;
 wire \u_cpu.REG_FILE._02807_ ;
 wire \u_cpu.REG_FILE._02808_ ;
 wire \u_cpu.REG_FILE._02809_ ;
 wire \u_cpu.REG_FILE._02810_ ;
 wire \u_cpu.REG_FILE._02811_ ;
 wire \u_cpu.REG_FILE._02812_ ;
 wire \u_cpu.REG_FILE._02813_ ;
 wire \u_cpu.REG_FILE._02814_ ;
 wire \u_cpu.REG_FILE._02815_ ;
 wire \u_cpu.REG_FILE._02816_ ;
 wire \u_cpu.REG_FILE._02817_ ;
 wire \u_cpu.REG_FILE._02818_ ;
 wire \u_cpu.REG_FILE._02819_ ;
 wire \u_cpu.REG_FILE._02820_ ;
 wire \u_cpu.REG_FILE._02821_ ;
 wire \u_cpu.REG_FILE._02822_ ;
 wire \u_cpu.REG_FILE._02823_ ;
 wire \u_cpu.REG_FILE._02824_ ;
 wire \u_cpu.REG_FILE._02825_ ;
 wire \u_cpu.REG_FILE._02826_ ;
 wire \u_cpu.REG_FILE._02827_ ;
 wire \u_cpu.REG_FILE._02828_ ;
 wire \u_cpu.REG_FILE._02829_ ;
 wire \u_cpu.REG_FILE._02830_ ;
 wire \u_cpu.REG_FILE._02831_ ;
 wire \u_cpu.REG_FILE._02832_ ;
 wire \u_cpu.REG_FILE._02833_ ;
 wire \u_cpu.REG_FILE._02834_ ;
 wire \u_cpu.REG_FILE._02835_ ;
 wire \u_cpu.REG_FILE._02836_ ;
 wire \u_cpu.REG_FILE._02837_ ;
 wire \u_cpu.REG_FILE._02838_ ;
 wire \u_cpu.REG_FILE._02839_ ;
 wire \u_cpu.REG_FILE._02840_ ;
 wire \u_cpu.REG_FILE._02841_ ;
 wire \u_cpu.REG_FILE._02842_ ;
 wire \u_cpu.REG_FILE._02843_ ;
 wire \u_cpu.REG_FILE._02844_ ;
 wire \u_cpu.REG_FILE._02845_ ;
 wire \u_cpu.REG_FILE._02846_ ;
 wire \u_cpu.REG_FILE._02847_ ;
 wire \u_cpu.REG_FILE._02848_ ;
 wire \u_cpu.REG_FILE._02849_ ;
 wire \u_cpu.REG_FILE._02850_ ;
 wire \u_cpu.REG_FILE._02851_ ;
 wire \u_cpu.REG_FILE._02852_ ;
 wire \u_cpu.REG_FILE._02853_ ;
 wire \u_cpu.REG_FILE._02854_ ;
 wire \u_cpu.REG_FILE._02855_ ;
 wire \u_cpu.REG_FILE._02856_ ;
 wire \u_cpu.REG_FILE._02857_ ;
 wire \u_cpu.REG_FILE._02858_ ;
 wire \u_cpu.REG_FILE._02859_ ;
 wire \u_cpu.REG_FILE._02860_ ;
 wire \u_cpu.REG_FILE._02861_ ;
 wire \u_cpu.REG_FILE._02862_ ;
 wire \u_cpu.REG_FILE._02863_ ;
 wire \u_cpu.REG_FILE._02864_ ;
 wire \u_cpu.REG_FILE._02865_ ;
 wire \u_cpu.REG_FILE._02866_ ;
 wire \u_cpu.REG_FILE._02867_ ;
 wire \u_cpu.REG_FILE._02868_ ;
 wire \u_cpu.REG_FILE._02869_ ;
 wire \u_cpu.REG_FILE._02870_ ;
 wire \u_cpu.REG_FILE._02871_ ;
 wire \u_cpu.REG_FILE._02872_ ;
 wire \u_cpu.REG_FILE._02873_ ;
 wire \u_cpu.REG_FILE._02874_ ;
 wire \u_cpu.REG_FILE._02875_ ;
 wire \u_cpu.REG_FILE._02876_ ;
 wire \u_cpu.REG_FILE._02877_ ;
 wire \u_cpu.REG_FILE._02878_ ;
 wire \u_cpu.REG_FILE._02879_ ;
 wire \u_cpu.REG_FILE._02880_ ;
 wire \u_cpu.REG_FILE._02881_ ;
 wire \u_cpu.REG_FILE._02882_ ;
 wire \u_cpu.REG_FILE._02883_ ;
 wire \u_cpu.REG_FILE._02884_ ;
 wire \u_cpu.REG_FILE._02885_ ;
 wire \u_cpu.REG_FILE._02886_ ;
 wire \u_cpu.REG_FILE._02887_ ;
 wire \u_cpu.REG_FILE._02888_ ;
 wire \u_cpu.REG_FILE._02889_ ;
 wire \u_cpu.REG_FILE._02890_ ;
 wire \u_cpu.REG_FILE._02891_ ;
 wire \u_cpu.REG_FILE._02892_ ;
 wire \u_cpu.REG_FILE._02893_ ;
 wire \u_cpu.REG_FILE._02894_ ;
 wire \u_cpu.REG_FILE._02895_ ;
 wire \u_cpu.REG_FILE._02896_ ;
 wire \u_cpu.REG_FILE._02897_ ;
 wire \u_cpu.REG_FILE._02898_ ;
 wire \u_cpu.REG_FILE._02899_ ;
 wire \u_cpu.REG_FILE._02900_ ;
 wire \u_cpu.REG_FILE._02901_ ;
 wire \u_cpu.REG_FILE._02902_ ;
 wire \u_cpu.REG_FILE._02903_ ;
 wire \u_cpu.REG_FILE._02904_ ;
 wire \u_cpu.REG_FILE._02905_ ;
 wire \u_cpu.REG_FILE._02906_ ;
 wire \u_cpu.REG_FILE._02907_ ;
 wire \u_cpu.REG_FILE._02908_ ;
 wire \u_cpu.REG_FILE._02909_ ;
 wire \u_cpu.REG_FILE._02910_ ;
 wire \u_cpu.REG_FILE._02911_ ;
 wire \u_cpu.REG_FILE._02912_ ;
 wire \u_cpu.REG_FILE._02913_ ;
 wire \u_cpu.REG_FILE._02914_ ;
 wire \u_cpu.REG_FILE._02915_ ;
 wire \u_cpu.REG_FILE._02916_ ;
 wire \u_cpu.REG_FILE._02917_ ;
 wire \u_cpu.REG_FILE._02918_ ;
 wire \u_cpu.REG_FILE._02919_ ;
 wire \u_cpu.REG_FILE._02920_ ;
 wire \u_cpu.REG_FILE._02921_ ;
 wire \u_cpu.REG_FILE._02922_ ;
 wire \u_cpu.REG_FILE._02923_ ;
 wire \u_cpu.REG_FILE._02924_ ;
 wire \u_cpu.REG_FILE._02925_ ;
 wire \u_cpu.REG_FILE._02926_ ;
 wire \u_cpu.REG_FILE._02927_ ;
 wire \u_cpu.REG_FILE._02928_ ;
 wire \u_cpu.REG_FILE._02929_ ;
 wire \u_cpu.REG_FILE._02930_ ;
 wire \u_cpu.REG_FILE._02931_ ;
 wire \u_cpu.REG_FILE._02932_ ;
 wire \u_cpu.REG_FILE._02933_ ;
 wire \u_cpu.REG_FILE._02934_ ;
 wire \u_cpu.REG_FILE._02935_ ;
 wire \u_cpu.REG_FILE._02936_ ;
 wire \u_cpu.REG_FILE._02937_ ;
 wire \u_cpu.REG_FILE._02938_ ;
 wire \u_cpu.REG_FILE._02939_ ;
 wire \u_cpu.REG_FILE._02940_ ;
 wire \u_cpu.REG_FILE._02941_ ;
 wire \u_cpu.REG_FILE._02942_ ;
 wire \u_cpu.REG_FILE._02943_ ;
 wire \u_cpu.REG_FILE._02944_ ;
 wire \u_cpu.REG_FILE._02945_ ;
 wire \u_cpu.REG_FILE._02946_ ;
 wire \u_cpu.REG_FILE._02947_ ;
 wire \u_cpu.REG_FILE._02948_ ;
 wire \u_cpu.REG_FILE._02949_ ;
 wire \u_cpu.REG_FILE._02950_ ;
 wire \u_cpu.REG_FILE._02951_ ;
 wire \u_cpu.REG_FILE._02952_ ;
 wire \u_cpu.REG_FILE._02953_ ;
 wire \u_cpu.REG_FILE._02954_ ;
 wire \u_cpu.REG_FILE._02955_ ;
 wire \u_cpu.REG_FILE._02956_ ;
 wire \u_cpu.REG_FILE._02957_ ;
 wire \u_cpu.REG_FILE._02958_ ;
 wire \u_cpu.REG_FILE._02959_ ;
 wire \u_cpu.REG_FILE._02960_ ;
 wire \u_cpu.REG_FILE._02961_ ;
 wire \u_cpu.REG_FILE._02962_ ;
 wire \u_cpu.REG_FILE._02963_ ;
 wire \u_cpu.REG_FILE._02964_ ;
 wire \u_cpu.REG_FILE._02965_ ;
 wire \u_cpu.REG_FILE._02966_ ;
 wire \u_cpu.REG_FILE._02967_ ;
 wire \u_cpu.REG_FILE._02968_ ;
 wire \u_cpu.REG_FILE._02969_ ;
 wire \u_cpu.REG_FILE._02970_ ;
 wire \u_cpu.REG_FILE._02971_ ;
 wire \u_cpu.REG_FILE._02972_ ;
 wire \u_cpu.REG_FILE._02973_ ;
 wire \u_cpu.REG_FILE._02974_ ;
 wire \u_cpu.REG_FILE._02975_ ;
 wire \u_cpu.REG_FILE._02976_ ;
 wire \u_cpu.REG_FILE._02977_ ;
 wire \u_cpu.REG_FILE._02978_ ;
 wire \u_cpu.REG_FILE._02979_ ;
 wire \u_cpu.REG_FILE._02980_ ;
 wire \u_cpu.REG_FILE._02981_ ;
 wire \u_cpu.REG_FILE._02982_ ;
 wire \u_cpu.REG_FILE._02983_ ;
 wire \u_cpu.REG_FILE._02984_ ;
 wire \u_cpu.REG_FILE._02985_ ;
 wire \u_cpu.REG_FILE._02986_ ;
 wire \u_cpu.REG_FILE._02987_ ;
 wire \u_cpu.REG_FILE._02988_ ;
 wire \u_cpu.REG_FILE._02989_ ;
 wire \u_cpu.REG_FILE._02990_ ;
 wire \u_cpu.REG_FILE._02991_ ;
 wire \u_cpu.REG_FILE._02992_ ;
 wire \u_cpu.REG_FILE._02993_ ;
 wire \u_cpu.REG_FILE._02994_ ;
 wire \u_cpu.REG_FILE._02995_ ;
 wire \u_cpu.REG_FILE._02996_ ;
 wire \u_cpu.REG_FILE._02997_ ;
 wire \u_cpu.REG_FILE._02998_ ;
 wire \u_cpu.REG_FILE._02999_ ;
 wire \u_cpu.REG_FILE._03000_ ;
 wire \u_cpu.REG_FILE._03001_ ;
 wire \u_cpu.REG_FILE._03002_ ;
 wire \u_cpu.REG_FILE._03003_ ;
 wire \u_cpu.REG_FILE._03004_ ;
 wire \u_cpu.REG_FILE._03005_ ;
 wire \u_cpu.REG_FILE._03006_ ;
 wire \u_cpu.REG_FILE._03007_ ;
 wire \u_cpu.REG_FILE._03008_ ;
 wire \u_cpu.REG_FILE._03009_ ;
 wire \u_cpu.REG_FILE._03010_ ;
 wire \u_cpu.REG_FILE._03011_ ;
 wire \u_cpu.REG_FILE._03012_ ;
 wire \u_cpu.REG_FILE._03013_ ;
 wire \u_cpu.REG_FILE._03014_ ;
 wire \u_cpu.REG_FILE._03015_ ;
 wire \u_cpu.REG_FILE._03016_ ;
 wire \u_cpu.REG_FILE._03017_ ;
 wire \u_cpu.REG_FILE._03018_ ;
 wire \u_cpu.REG_FILE._03019_ ;
 wire \u_cpu.REG_FILE._03020_ ;
 wire \u_cpu.REG_FILE._03021_ ;
 wire \u_cpu.REG_FILE._03022_ ;
 wire \u_cpu.REG_FILE._03023_ ;
 wire \u_cpu.REG_FILE._03024_ ;
 wire \u_cpu.REG_FILE._03025_ ;
 wire \u_cpu.REG_FILE._03026_ ;
 wire \u_cpu.REG_FILE._03027_ ;
 wire \u_cpu.REG_FILE._03028_ ;
 wire \u_cpu.REG_FILE._03029_ ;
 wire \u_cpu.REG_FILE._03030_ ;
 wire \u_cpu.REG_FILE._03031_ ;
 wire \u_cpu.REG_FILE._03032_ ;
 wire \u_cpu.REG_FILE._03033_ ;
 wire \u_cpu.REG_FILE._03034_ ;
 wire \u_cpu.REG_FILE._03035_ ;
 wire \u_cpu.REG_FILE._03036_ ;
 wire \u_cpu.REG_FILE._03037_ ;
 wire \u_cpu.REG_FILE._03038_ ;
 wire \u_cpu.REG_FILE._03039_ ;
 wire \u_cpu.REG_FILE._03040_ ;
 wire \u_cpu.REG_FILE._03041_ ;
 wire \u_cpu.REG_FILE._03042_ ;
 wire \u_cpu.REG_FILE._03043_ ;
 wire \u_cpu.REG_FILE._03044_ ;
 wire \u_cpu.REG_FILE._03045_ ;
 wire \u_cpu.REG_FILE._03046_ ;
 wire \u_cpu.REG_FILE._03047_ ;
 wire \u_cpu.REG_FILE._03048_ ;
 wire \u_cpu.REG_FILE._03049_ ;
 wire \u_cpu.REG_FILE._03050_ ;
 wire \u_cpu.REG_FILE._03051_ ;
 wire \u_cpu.REG_FILE._03052_ ;
 wire \u_cpu.REG_FILE._03053_ ;
 wire \u_cpu.REG_FILE._03054_ ;
 wire \u_cpu.REG_FILE._03055_ ;
 wire \u_cpu.REG_FILE._03056_ ;
 wire \u_cpu.REG_FILE._03057_ ;
 wire \u_cpu.REG_FILE._03058_ ;
 wire \u_cpu.REG_FILE._03059_ ;
 wire \u_cpu.REG_FILE._03060_ ;
 wire \u_cpu.REG_FILE._03061_ ;
 wire \u_cpu.REG_FILE._03062_ ;
 wire \u_cpu.REG_FILE._03063_ ;
 wire \u_cpu.REG_FILE._03064_ ;
 wire \u_cpu.REG_FILE._03065_ ;
 wire \u_cpu.REG_FILE._03066_ ;
 wire \u_cpu.REG_FILE._03067_ ;
 wire \u_cpu.REG_FILE._03068_ ;
 wire \u_cpu.REG_FILE._03069_ ;
 wire \u_cpu.REG_FILE._03070_ ;
 wire \u_cpu.REG_FILE._03071_ ;
 wire \u_cpu.REG_FILE._03072_ ;
 wire \u_cpu.REG_FILE._03073_ ;
 wire \u_cpu.REG_FILE._03074_ ;
 wire \u_cpu.REG_FILE._03075_ ;
 wire \u_cpu.REG_FILE._03076_ ;
 wire \u_cpu.REG_FILE._03077_ ;
 wire \u_cpu.REG_FILE._03078_ ;
 wire \u_cpu.REG_FILE._03079_ ;
 wire \u_cpu.REG_FILE._03080_ ;
 wire \u_cpu.REG_FILE._03081_ ;
 wire \u_cpu.REG_FILE._03082_ ;
 wire \u_cpu.REG_FILE._03083_ ;
 wire \u_cpu.REG_FILE._03084_ ;
 wire \u_cpu.REG_FILE._03085_ ;
 wire \u_cpu.REG_FILE._03086_ ;
 wire \u_cpu.REG_FILE._03087_ ;
 wire \u_cpu.REG_FILE._03088_ ;
 wire \u_cpu.REG_FILE._03089_ ;
 wire \u_cpu.REG_FILE._03090_ ;
 wire \u_cpu.REG_FILE._03091_ ;
 wire \u_cpu.REG_FILE._03092_ ;
 wire \u_cpu.REG_FILE._03093_ ;
 wire \u_cpu.REG_FILE._03094_ ;
 wire \u_cpu.REG_FILE._03095_ ;
 wire \u_cpu.REG_FILE._03096_ ;
 wire \u_cpu.REG_FILE._03097_ ;
 wire \u_cpu.REG_FILE._03098_ ;
 wire \u_cpu.REG_FILE._03099_ ;
 wire \u_cpu.REG_FILE._03100_ ;
 wire \u_cpu.REG_FILE._03101_ ;
 wire \u_cpu.REG_FILE._03102_ ;
 wire \u_cpu.REG_FILE._03103_ ;
 wire \u_cpu.REG_FILE._03104_ ;
 wire \u_cpu.REG_FILE._03105_ ;
 wire \u_cpu.REG_FILE._03106_ ;
 wire \u_cpu.REG_FILE._03107_ ;
 wire \u_cpu.REG_FILE._03108_ ;
 wire \u_cpu.REG_FILE._03109_ ;
 wire \u_cpu.REG_FILE._03110_ ;
 wire \u_cpu.REG_FILE._03111_ ;
 wire \u_cpu.REG_FILE._03112_ ;
 wire \u_cpu.REG_FILE._03113_ ;
 wire \u_cpu.REG_FILE._03114_ ;
 wire \u_cpu.REG_FILE._03115_ ;
 wire \u_cpu.REG_FILE._03116_ ;
 wire \u_cpu.REG_FILE._03117_ ;
 wire \u_cpu.REG_FILE._03118_ ;
 wire \u_cpu.REG_FILE._03119_ ;
 wire \u_cpu.REG_FILE._03120_ ;
 wire \u_cpu.REG_FILE._03121_ ;
 wire \u_cpu.REG_FILE._03122_ ;
 wire \u_cpu.REG_FILE._03123_ ;
 wire \u_cpu.REG_FILE._03124_ ;
 wire \u_cpu.REG_FILE._03125_ ;
 wire \u_cpu.REG_FILE._03126_ ;
 wire \u_cpu.REG_FILE._03127_ ;
 wire \u_cpu.REG_FILE._03128_ ;
 wire \u_cpu.REG_FILE._03129_ ;
 wire \u_cpu.REG_FILE._03130_ ;
 wire \u_cpu.REG_FILE._03131_ ;
 wire \u_cpu.REG_FILE._03132_ ;
 wire \u_cpu.REG_FILE._03133_ ;
 wire \u_cpu.REG_FILE._03134_ ;
 wire \u_cpu.REG_FILE._03135_ ;
 wire \u_cpu.REG_FILE._03136_ ;
 wire \u_cpu.REG_FILE._03137_ ;
 wire \u_cpu.REG_FILE._03138_ ;
 wire \u_cpu.REG_FILE._03139_ ;
 wire \u_cpu.REG_FILE._03140_ ;
 wire \u_cpu.REG_FILE._03141_ ;
 wire \u_cpu.REG_FILE._03142_ ;
 wire \u_cpu.REG_FILE._03143_ ;
 wire \u_cpu.REG_FILE._03144_ ;
 wire \u_cpu.REG_FILE._03145_ ;
 wire \u_cpu.REG_FILE._03146_ ;
 wire \u_cpu.REG_FILE._03147_ ;
 wire \u_cpu.REG_FILE._03148_ ;
 wire \u_cpu.REG_FILE._03149_ ;
 wire \u_cpu.REG_FILE._03150_ ;
 wire \u_cpu.REG_FILE._03151_ ;
 wire \u_cpu.REG_FILE._03152_ ;
 wire \u_cpu.REG_FILE._03153_ ;
 wire \u_cpu.REG_FILE._03154_ ;
 wire \u_cpu.REG_FILE._03155_ ;
 wire \u_cpu.REG_FILE._03156_ ;
 wire \u_cpu.REG_FILE._03157_ ;
 wire \u_cpu.REG_FILE._03158_ ;
 wire \u_cpu.REG_FILE._03159_ ;
 wire \u_cpu.REG_FILE._03160_ ;
 wire \u_cpu.REG_FILE._03161_ ;
 wire \u_cpu.REG_FILE._03162_ ;
 wire \u_cpu.REG_FILE._03163_ ;
 wire \u_cpu.REG_FILE._03164_ ;
 wire \u_cpu.REG_FILE._03165_ ;
 wire \u_cpu.REG_FILE._03166_ ;
 wire \u_cpu.REG_FILE._03167_ ;
 wire \u_cpu.REG_FILE._03168_ ;
 wire \u_cpu.REG_FILE._03169_ ;
 wire \u_cpu.REG_FILE._03170_ ;
 wire \u_cpu.REG_FILE._03171_ ;
 wire \u_cpu.REG_FILE._03172_ ;
 wire \u_cpu.REG_FILE._03173_ ;
 wire \u_cpu.REG_FILE._03174_ ;
 wire \u_cpu.REG_FILE._03175_ ;
 wire \u_cpu.REG_FILE._03176_ ;
 wire \u_cpu.REG_FILE._03177_ ;
 wire \u_cpu.REG_FILE._03178_ ;
 wire \u_cpu.REG_FILE._03179_ ;
 wire \u_cpu.REG_FILE._03180_ ;
 wire \u_cpu.REG_FILE._03181_ ;
 wire \u_cpu.REG_FILE._03182_ ;
 wire \u_cpu.REG_FILE._03183_ ;
 wire \u_cpu.REG_FILE._03184_ ;
 wire \u_cpu.REG_FILE._03185_ ;
 wire \u_cpu.REG_FILE._03186_ ;
 wire \u_cpu.REG_FILE._03187_ ;
 wire \u_cpu.REG_FILE._03188_ ;
 wire \u_cpu.REG_FILE._03189_ ;
 wire \u_cpu.REG_FILE._03190_ ;
 wire \u_cpu.REG_FILE._03191_ ;
 wire \u_cpu.REG_FILE._03192_ ;
 wire \u_cpu.REG_FILE._03193_ ;
 wire \u_cpu.REG_FILE._03194_ ;
 wire \u_cpu.REG_FILE._03195_ ;
 wire \u_cpu.REG_FILE._03196_ ;
 wire \u_cpu.REG_FILE._03197_ ;
 wire \u_cpu.REG_FILE._03198_ ;
 wire \u_cpu.REG_FILE._03199_ ;
 wire \u_cpu.REG_FILE._03200_ ;
 wire \u_cpu.REG_FILE._03201_ ;
 wire \u_cpu.REG_FILE._03202_ ;
 wire \u_cpu.REG_FILE._03203_ ;
 wire \u_cpu.REG_FILE._03204_ ;
 wire \u_cpu.REG_FILE._03205_ ;
 wire \u_cpu.REG_FILE._03206_ ;
 wire \u_cpu.REG_FILE._03207_ ;
 wire \u_cpu.REG_FILE._03208_ ;
 wire \u_cpu.REG_FILE._03209_ ;
 wire \u_cpu.REG_FILE._03210_ ;
 wire \u_cpu.REG_FILE._03211_ ;
 wire \u_cpu.REG_FILE._03212_ ;
 wire \u_cpu.REG_FILE._03213_ ;
 wire \u_cpu.REG_FILE._03214_ ;
 wire \u_cpu.REG_FILE._03215_ ;
 wire \u_cpu.REG_FILE._03216_ ;
 wire \u_cpu.REG_FILE._03217_ ;
 wire \u_cpu.REG_FILE._03218_ ;
 wire \u_cpu.REG_FILE._03219_ ;
 wire \u_cpu.REG_FILE._03220_ ;
 wire \u_cpu.REG_FILE._03221_ ;
 wire \u_cpu.REG_FILE._03222_ ;
 wire \u_cpu.REG_FILE._03223_ ;
 wire \u_cpu.REG_FILE._03224_ ;
 wire \u_cpu.REG_FILE._03225_ ;
 wire \u_cpu.REG_FILE._03226_ ;
 wire \u_cpu.REG_FILE._03227_ ;
 wire \u_cpu.REG_FILE._03228_ ;
 wire \u_cpu.REG_FILE._03229_ ;
 wire \u_cpu.REG_FILE._03230_ ;
 wire \u_cpu.REG_FILE._03231_ ;
 wire \u_cpu.REG_FILE._03232_ ;
 wire \u_cpu.REG_FILE._03233_ ;
 wire \u_cpu.REG_FILE._03234_ ;
 wire \u_cpu.REG_FILE._03235_ ;
 wire \u_cpu.REG_FILE._03236_ ;
 wire \u_cpu.REG_FILE._03237_ ;
 wire \u_cpu.REG_FILE._03238_ ;
 wire \u_cpu.REG_FILE._03239_ ;
 wire \u_cpu.REG_FILE._03240_ ;
 wire \u_cpu.REG_FILE._03241_ ;
 wire \u_cpu.REG_FILE._03242_ ;
 wire \u_cpu.REG_FILE._03243_ ;
 wire \u_cpu.REG_FILE._03244_ ;
 wire \u_cpu.REG_FILE._03245_ ;
 wire \u_cpu.REG_FILE._03246_ ;
 wire \u_cpu.REG_FILE._03247_ ;
 wire \u_cpu.REG_FILE._03248_ ;
 wire \u_cpu.REG_FILE._03249_ ;
 wire \u_cpu.REG_FILE._03250_ ;
 wire \u_cpu.REG_FILE._03251_ ;
 wire \u_cpu.REG_FILE._03252_ ;
 wire \u_cpu.REG_FILE._03253_ ;
 wire \u_cpu.REG_FILE._03254_ ;
 wire \u_cpu.REG_FILE._03255_ ;
 wire \u_cpu.REG_FILE._03256_ ;
 wire \u_cpu.REG_FILE._03257_ ;
 wire \u_cpu.REG_FILE._03258_ ;
 wire \u_cpu.REG_FILE._03259_ ;
 wire \u_cpu.REG_FILE._03260_ ;
 wire \u_cpu.REG_FILE._03261_ ;
 wire \u_cpu.REG_FILE._03262_ ;
 wire \u_cpu.REG_FILE._03263_ ;
 wire \u_cpu.REG_FILE._03264_ ;
 wire \u_cpu.REG_FILE._03265_ ;
 wire \u_cpu.REG_FILE._03266_ ;
 wire \u_cpu.REG_FILE._03267_ ;
 wire \u_cpu.REG_FILE._03268_ ;
 wire \u_cpu.REG_FILE._03269_ ;
 wire \u_cpu.REG_FILE._03270_ ;
 wire \u_cpu.REG_FILE._03271_ ;
 wire \u_cpu.REG_FILE._03272_ ;
 wire \u_cpu.REG_FILE._03273_ ;
 wire \u_cpu.REG_FILE._03274_ ;
 wire \u_cpu.REG_FILE._03275_ ;
 wire \u_cpu.REG_FILE._03276_ ;
 wire \u_cpu.REG_FILE._03277_ ;
 wire \u_cpu.REG_FILE._03278_ ;
 wire \u_cpu.REG_FILE._03279_ ;
 wire \u_cpu.REG_FILE._03280_ ;
 wire \u_cpu.REG_FILE._03281_ ;
 wire \u_cpu.REG_FILE._03282_ ;
 wire \u_cpu.REG_FILE._03283_ ;
 wire \u_cpu.REG_FILE._03284_ ;
 wire \u_cpu.REG_FILE._03285_ ;
 wire \u_cpu.REG_FILE._03286_ ;
 wire \u_cpu.REG_FILE._03287_ ;
 wire \u_cpu.REG_FILE._03288_ ;
 wire \u_cpu.REG_FILE._03289_ ;
 wire \u_cpu.REG_FILE._03290_ ;
 wire \u_cpu.REG_FILE._03291_ ;
 wire \u_cpu.REG_FILE._03292_ ;
 wire \u_cpu.REG_FILE._03293_ ;
 wire \u_cpu.REG_FILE._03294_ ;
 wire \u_cpu.REG_FILE._03295_ ;
 wire \u_cpu.REG_FILE._03296_ ;
 wire \u_cpu.REG_FILE._03297_ ;
 wire \u_cpu.REG_FILE._03298_ ;
 wire \u_cpu.REG_FILE._03299_ ;
 wire \u_cpu.REG_FILE._03300_ ;
 wire \u_cpu.REG_FILE._03301_ ;
 wire \u_cpu.REG_FILE._03302_ ;
 wire \u_cpu.REG_FILE._03303_ ;
 wire \u_cpu.REG_FILE._03304_ ;
 wire \u_cpu.REG_FILE._03305_ ;
 wire \u_cpu.REG_FILE._03306_ ;
 wire \u_cpu.REG_FILE._03307_ ;
 wire \u_cpu.REG_FILE._03308_ ;
 wire \u_cpu.REG_FILE._03309_ ;
 wire \u_cpu.REG_FILE._03310_ ;
 wire \u_cpu.REG_FILE._03311_ ;
 wire \u_cpu.REG_FILE._03312_ ;
 wire \u_cpu.REG_FILE._03313_ ;
 wire \u_cpu.REG_FILE._03314_ ;
 wire \u_cpu.REG_FILE._03315_ ;
 wire \u_cpu.REG_FILE._03316_ ;
 wire \u_cpu.REG_FILE._03317_ ;
 wire \u_cpu.REG_FILE._03318_ ;
 wire \u_cpu.REG_FILE._03319_ ;
 wire \u_cpu.REG_FILE._03320_ ;
 wire \u_cpu.REG_FILE._03321_ ;
 wire \u_cpu.REG_FILE._03322_ ;
 wire \u_cpu.REG_FILE._03323_ ;
 wire \u_cpu.REG_FILE._03324_ ;
 wire \u_cpu.REG_FILE._03325_ ;
 wire \u_cpu.REG_FILE._03326_ ;
 wire \u_cpu.REG_FILE._03327_ ;
 wire \u_cpu.REG_FILE._03328_ ;
 wire \u_cpu.REG_FILE._03329_ ;
 wire \u_cpu.REG_FILE._03330_ ;
 wire \u_cpu.REG_FILE._03331_ ;
 wire \u_cpu.REG_FILE._03332_ ;
 wire \u_cpu.REG_FILE._03333_ ;
 wire \u_cpu.REG_FILE._03334_ ;
 wire \u_cpu.REG_FILE._03335_ ;
 wire \u_cpu.REG_FILE._03336_ ;
 wire \u_cpu.REG_FILE._03337_ ;
 wire \u_cpu.REG_FILE._03338_ ;
 wire \u_cpu.REG_FILE._03339_ ;
 wire \u_cpu.REG_FILE._03340_ ;
 wire \u_cpu.REG_FILE._03341_ ;
 wire \u_cpu.REG_FILE._03342_ ;
 wire \u_cpu.REG_FILE._03343_ ;
 wire \u_cpu.REG_FILE._03344_ ;
 wire \u_cpu.REG_FILE._03345_ ;
 wire \u_cpu.REG_FILE._03346_ ;
 wire \u_cpu.REG_FILE._03347_ ;
 wire \u_cpu.REG_FILE._03348_ ;
 wire \u_cpu.REG_FILE._03349_ ;
 wire \u_cpu.REG_FILE._03350_ ;
 wire \u_cpu.REG_FILE._03351_ ;
 wire \u_cpu.REG_FILE._03352_ ;
 wire \u_cpu.REG_FILE._03353_ ;
 wire \u_cpu.REG_FILE._03354_ ;
 wire \u_cpu.REG_FILE._03355_ ;
 wire \u_cpu.REG_FILE._03356_ ;
 wire \u_cpu.REG_FILE._03357_ ;
 wire \u_cpu.REG_FILE._03358_ ;
 wire \u_cpu.REG_FILE._03359_ ;
 wire \u_cpu.REG_FILE._03360_ ;
 wire \u_cpu.REG_FILE._03361_ ;
 wire \u_cpu.REG_FILE._03362_ ;
 wire \u_cpu.REG_FILE._03363_ ;
 wire \u_cpu.REG_FILE._03364_ ;
 wire \u_cpu.REG_FILE._03365_ ;
 wire \u_cpu.REG_FILE._03366_ ;
 wire \u_cpu.REG_FILE._03367_ ;
 wire \u_cpu.REG_FILE._03368_ ;
 wire \u_cpu.REG_FILE._03369_ ;
 wire \u_cpu.REG_FILE._03370_ ;
 wire \u_cpu.REG_FILE._03371_ ;
 wire \u_cpu.REG_FILE._03372_ ;
 wire \u_cpu.REG_FILE._03373_ ;
 wire \u_cpu.REG_FILE._03374_ ;
 wire \u_cpu.REG_FILE._03375_ ;
 wire \u_cpu.REG_FILE._03376_ ;
 wire \u_cpu.REG_FILE._03377_ ;
 wire \u_cpu.REG_FILE._03378_ ;
 wire \u_cpu.REG_FILE._03379_ ;
 wire \u_cpu.REG_FILE._03380_ ;
 wire \u_cpu.REG_FILE._03381_ ;
 wire \u_cpu.REG_FILE._03382_ ;
 wire \u_cpu.REG_FILE._03383_ ;
 wire \u_cpu.REG_FILE._03384_ ;
 wire \u_cpu.REG_FILE._03385_ ;
 wire \u_cpu.REG_FILE._03386_ ;
 wire \u_cpu.REG_FILE._03387_ ;
 wire \u_cpu.REG_FILE._03388_ ;
 wire \u_cpu.REG_FILE._03389_ ;
 wire \u_cpu.REG_FILE._03390_ ;
 wire \u_cpu.REG_FILE._03391_ ;
 wire \u_cpu.REG_FILE._03392_ ;
 wire \u_cpu.REG_FILE._03393_ ;
 wire \u_cpu.REG_FILE._03394_ ;
 wire \u_cpu.REG_FILE._03395_ ;
 wire \u_cpu.REG_FILE._03396_ ;
 wire \u_cpu.REG_FILE._03397_ ;
 wire \u_cpu.REG_FILE._03398_ ;
 wire \u_cpu.REG_FILE._03399_ ;
 wire \u_cpu.REG_FILE._03400_ ;
 wire \u_cpu.REG_FILE._03401_ ;
 wire \u_cpu.REG_FILE._03402_ ;
 wire \u_cpu.REG_FILE._03403_ ;
 wire \u_cpu.REG_FILE._03404_ ;
 wire \u_cpu.REG_FILE._03405_ ;
 wire \u_cpu.REG_FILE._03406_ ;
 wire \u_cpu.REG_FILE._03407_ ;
 wire \u_cpu.REG_FILE._03408_ ;
 wire \u_cpu.REG_FILE._03409_ ;
 wire \u_cpu.REG_FILE._03410_ ;
 wire \u_cpu.REG_FILE._03411_ ;
 wire \u_cpu.REG_FILE._03412_ ;
 wire \u_cpu.REG_FILE._03413_ ;
 wire \u_cpu.REG_FILE._03414_ ;
 wire \u_cpu.REG_FILE._03415_ ;
 wire \u_cpu.REG_FILE._03416_ ;
 wire \u_cpu.REG_FILE._03417_ ;
 wire \u_cpu.REG_FILE._03418_ ;
 wire \u_cpu.REG_FILE._03419_ ;
 wire \u_cpu.REG_FILE._03420_ ;
 wire \u_cpu.REG_FILE._03421_ ;
 wire \u_cpu.REG_FILE._03422_ ;
 wire \u_cpu.REG_FILE._03423_ ;
 wire \u_cpu.REG_FILE._03424_ ;
 wire \u_cpu.REG_FILE._03425_ ;
 wire \u_cpu.REG_FILE._03426_ ;
 wire \u_cpu.REG_FILE._03427_ ;
 wire \u_cpu.REG_FILE._03428_ ;
 wire \u_cpu.REG_FILE._03429_ ;
 wire \u_cpu.REG_FILE._03430_ ;
 wire \u_cpu.REG_FILE._03431_ ;
 wire \u_cpu.REG_FILE._03432_ ;
 wire \u_cpu.REG_FILE._03433_ ;
 wire \u_cpu.REG_FILE._03434_ ;
 wire \u_cpu.REG_FILE._03435_ ;
 wire \u_cpu.REG_FILE._03436_ ;
 wire \u_cpu.REG_FILE._03437_ ;
 wire \u_cpu.REG_FILE._03438_ ;
 wire \u_cpu.REG_FILE._03439_ ;
 wire \u_cpu.REG_FILE._03440_ ;
 wire \u_cpu.REG_FILE._03441_ ;
 wire \u_cpu.REG_FILE._03442_ ;
 wire \u_cpu.REG_FILE._03443_ ;
 wire \u_cpu.REG_FILE._03444_ ;
 wire \u_cpu.REG_FILE._03445_ ;
 wire \u_cpu.REG_FILE._03446_ ;
 wire \u_cpu.REG_FILE._03447_ ;
 wire \u_cpu.REG_FILE._03448_ ;
 wire \u_cpu.REG_FILE._03449_ ;
 wire \u_cpu.REG_FILE._03450_ ;
 wire \u_cpu.REG_FILE._03451_ ;
 wire \u_cpu.REG_FILE._03452_ ;
 wire \u_cpu.REG_FILE._03453_ ;
 wire \u_cpu.REG_FILE._03454_ ;
 wire \u_cpu.REG_FILE._03455_ ;
 wire \u_cpu.REG_FILE._03456_ ;
 wire \u_cpu.REG_FILE._03457_ ;
 wire \u_cpu.REG_FILE._03458_ ;
 wire \u_cpu.REG_FILE._03459_ ;
 wire \u_cpu.REG_FILE._03460_ ;
 wire \u_cpu.REG_FILE._03461_ ;
 wire \u_cpu.REG_FILE._03462_ ;
 wire \u_cpu.REG_FILE._03463_ ;
 wire \u_cpu.REG_FILE._03464_ ;
 wire \u_cpu.REG_FILE._03465_ ;
 wire \u_cpu.REG_FILE._03466_ ;
 wire \u_cpu.REG_FILE._03467_ ;
 wire \u_cpu.REG_FILE._03468_ ;
 wire \u_cpu.REG_FILE._03469_ ;
 wire \u_cpu.REG_FILE._03470_ ;
 wire \u_cpu.REG_FILE._03471_ ;
 wire \u_cpu.REG_FILE._03472_ ;
 wire \u_cpu.REG_FILE._03473_ ;
 wire \u_cpu.REG_FILE._03474_ ;
 wire \u_cpu.REG_FILE._03475_ ;
 wire \u_cpu.REG_FILE._03476_ ;
 wire \u_cpu.REG_FILE._03477_ ;
 wire \u_cpu.REG_FILE._03478_ ;
 wire \u_cpu.REG_FILE._03479_ ;
 wire \u_cpu.REG_FILE._03480_ ;
 wire \u_cpu.REG_FILE._03481_ ;
 wire \u_cpu.REG_FILE._03482_ ;
 wire \u_cpu.REG_FILE._03483_ ;
 wire \u_cpu.REG_FILE._03484_ ;
 wire \u_cpu.REG_FILE._03485_ ;
 wire \u_cpu.REG_FILE._03486_ ;
 wire \u_cpu.REG_FILE._03487_ ;
 wire \u_cpu.REG_FILE._03488_ ;
 wire \u_cpu.REG_FILE._03489_ ;
 wire \u_cpu.REG_FILE._03490_ ;
 wire \u_cpu.REG_FILE._03491_ ;
 wire \u_cpu.REG_FILE._03492_ ;
 wire \u_cpu.REG_FILE._03493_ ;
 wire \u_cpu.REG_FILE._03494_ ;
 wire \u_cpu.REG_FILE._03495_ ;
 wire \u_cpu.REG_FILE._03496_ ;
 wire \u_cpu.REG_FILE._03497_ ;
 wire \u_cpu.REG_FILE._03498_ ;
 wire \u_cpu.REG_FILE._03499_ ;
 wire \u_cpu.REG_FILE._03500_ ;
 wire \u_cpu.REG_FILE._03501_ ;
 wire \u_cpu.REG_FILE._03502_ ;
 wire \u_cpu.REG_FILE._03503_ ;
 wire \u_cpu.REG_FILE._03504_ ;
 wire \u_cpu.REG_FILE._03505_ ;
 wire \u_cpu.REG_FILE._03506_ ;
 wire \u_cpu.REG_FILE._03507_ ;
 wire \u_cpu.REG_FILE._03508_ ;
 wire \u_cpu.REG_FILE._03509_ ;
 wire \u_cpu.REG_FILE._03510_ ;
 wire \u_cpu.REG_FILE._03511_ ;
 wire \u_cpu.REG_FILE._03512_ ;
 wire \u_cpu.REG_FILE._03513_ ;
 wire \u_cpu.REG_FILE._03514_ ;
 wire \u_cpu.REG_FILE._03515_ ;
 wire \u_cpu.REG_FILE._03516_ ;
 wire \u_cpu.REG_FILE._03517_ ;
 wire \u_cpu.REG_FILE._03518_ ;
 wire \u_cpu.REG_FILE._03519_ ;
 wire \u_cpu.REG_FILE._03520_ ;
 wire \u_cpu.REG_FILE._03521_ ;
 wire \u_cpu.REG_FILE._03522_ ;
 wire \u_cpu.REG_FILE._03523_ ;
 wire \u_cpu.REG_FILE._03524_ ;
 wire \u_cpu.REG_FILE._03525_ ;
 wire \u_cpu.REG_FILE._03526_ ;
 wire \u_cpu.REG_FILE._03527_ ;
 wire \u_cpu.REG_FILE._03528_ ;
 wire \u_cpu.REG_FILE._03529_ ;
 wire \u_cpu.REG_FILE._03530_ ;
 wire \u_cpu.REG_FILE._03531_ ;
 wire \u_cpu.REG_FILE._03532_ ;
 wire \u_cpu.REG_FILE._03533_ ;
 wire \u_cpu.REG_FILE._03534_ ;
 wire \u_cpu.REG_FILE._03535_ ;
 wire \u_cpu.REG_FILE._03536_ ;
 wire \u_cpu.REG_FILE._03537_ ;
 wire \u_cpu.REG_FILE._03538_ ;
 wire \u_cpu.REG_FILE._03539_ ;
 wire \u_cpu.REG_FILE._03540_ ;
 wire \u_cpu.REG_FILE._03541_ ;
 wire \u_cpu.REG_FILE._03542_ ;
 wire \u_cpu.REG_FILE._03543_ ;
 wire \u_cpu.REG_FILE._03544_ ;
 wire \u_cpu.REG_FILE._03545_ ;
 wire \u_cpu.REG_FILE._03546_ ;
 wire \u_cpu.REG_FILE._03547_ ;
 wire \u_cpu.REG_FILE._03548_ ;
 wire \u_cpu.REG_FILE._03549_ ;
 wire \u_cpu.REG_FILE._03550_ ;
 wire \u_cpu.REG_FILE._03551_ ;
 wire \u_cpu.REG_FILE._03552_ ;
 wire \u_cpu.REG_FILE._03553_ ;
 wire \u_cpu.REG_FILE._03554_ ;
 wire \u_cpu.REG_FILE._03555_ ;
 wire \u_cpu.REG_FILE._03556_ ;
 wire \u_cpu.REG_FILE._03557_ ;
 wire \u_cpu.REG_FILE._03558_ ;
 wire \u_cpu.REG_FILE._03559_ ;
 wire \u_cpu.REG_FILE._03560_ ;
 wire \u_cpu.REG_FILE._03561_ ;
 wire \u_cpu.REG_FILE._03562_ ;
 wire \u_cpu.REG_FILE._03563_ ;
 wire \u_cpu.REG_FILE._03564_ ;
 wire \u_cpu.REG_FILE._03565_ ;
 wire \u_cpu.REG_FILE._03566_ ;
 wire \u_cpu.REG_FILE._03567_ ;
 wire \u_cpu.REG_FILE._03568_ ;
 wire \u_cpu.REG_FILE._03569_ ;
 wire \u_cpu.REG_FILE._03570_ ;
 wire \u_cpu.REG_FILE._03571_ ;
 wire \u_cpu.REG_FILE._03572_ ;
 wire \u_cpu.REG_FILE._03573_ ;
 wire \u_cpu.REG_FILE._03574_ ;
 wire \u_cpu.REG_FILE._03575_ ;
 wire \u_cpu.REG_FILE._03576_ ;
 wire \u_cpu.REG_FILE._03577_ ;
 wire \u_cpu.REG_FILE._03578_ ;
 wire \u_cpu.REG_FILE._03579_ ;
 wire \u_cpu.REG_FILE._03580_ ;
 wire \u_cpu.REG_FILE._03581_ ;
 wire \u_cpu.REG_FILE._03582_ ;
 wire \u_cpu.REG_FILE._03583_ ;
 wire \u_cpu.REG_FILE._03584_ ;
 wire \u_cpu.REG_FILE._03585_ ;
 wire \u_cpu.REG_FILE._03586_ ;
 wire \u_cpu.REG_FILE._03587_ ;
 wire \u_cpu.REG_FILE._03588_ ;
 wire \u_cpu.REG_FILE._03589_ ;
 wire \u_cpu.REG_FILE._03590_ ;
 wire \u_cpu.REG_FILE._03591_ ;
 wire \u_cpu.REG_FILE._03592_ ;
 wire \u_cpu.REG_FILE._03593_ ;
 wire \u_cpu.REG_FILE._03594_ ;
 wire \u_cpu.REG_FILE._03595_ ;
 wire \u_cpu.REG_FILE._03596_ ;
 wire \u_cpu.REG_FILE._03597_ ;
 wire \u_cpu.REG_FILE._03598_ ;
 wire \u_cpu.REG_FILE._03599_ ;
 wire \u_cpu.REG_FILE._03600_ ;
 wire \u_cpu.REG_FILE._03601_ ;
 wire \u_cpu.REG_FILE._03602_ ;
 wire \u_cpu.REG_FILE._03603_ ;
 wire \u_cpu.REG_FILE._03604_ ;
 wire \u_cpu.REG_FILE._03605_ ;
 wire \u_cpu.REG_FILE._03606_ ;
 wire \u_cpu.REG_FILE._03607_ ;
 wire \u_cpu.REG_FILE._03608_ ;
 wire \u_cpu.REG_FILE._03609_ ;
 wire \u_cpu.REG_FILE._03610_ ;
 wire \u_cpu.REG_FILE._03611_ ;
 wire \u_cpu.REG_FILE._03612_ ;
 wire \u_cpu.REG_FILE._03613_ ;
 wire \u_cpu.REG_FILE._03614_ ;
 wire \u_cpu.REG_FILE._03615_ ;
 wire \u_cpu.REG_FILE._03616_ ;
 wire \u_cpu.REG_FILE._03617_ ;
 wire \u_cpu.REG_FILE._03618_ ;
 wire \u_cpu.REG_FILE._03619_ ;
 wire \u_cpu.REG_FILE._03620_ ;
 wire \u_cpu.REG_FILE._03621_ ;
 wire \u_cpu.REG_FILE._03622_ ;
 wire \u_cpu.REG_FILE._03623_ ;
 wire \u_cpu.REG_FILE._03624_ ;
 wire \u_cpu.REG_FILE._03625_ ;
 wire \u_cpu.REG_FILE._03626_ ;
 wire \u_cpu.REG_FILE._03627_ ;
 wire \u_cpu.REG_FILE._03628_ ;
 wire \u_cpu.REG_FILE._03629_ ;
 wire \u_cpu.REG_FILE._03630_ ;
 wire \u_cpu.REG_FILE._03631_ ;
 wire \u_cpu.REG_FILE._03632_ ;
 wire \u_cpu.REG_FILE._03633_ ;
 wire \u_cpu.REG_FILE._03634_ ;
 wire \u_cpu.REG_FILE._03635_ ;
 wire \u_cpu.REG_FILE._03636_ ;
 wire \u_cpu.REG_FILE._03637_ ;
 wire \u_cpu.REG_FILE._03638_ ;
 wire \u_cpu.REG_FILE._03639_ ;
 wire \u_cpu.REG_FILE._03640_ ;
 wire \u_cpu.REG_FILE._03641_ ;
 wire \u_cpu.REG_FILE._03642_ ;
 wire \u_cpu.REG_FILE._03643_ ;
 wire \u_cpu.REG_FILE._03644_ ;
 wire \u_cpu.REG_FILE._03645_ ;
 wire \u_cpu.REG_FILE._03646_ ;
 wire \u_cpu.REG_FILE._03647_ ;
 wire \u_cpu.REG_FILE._03648_ ;
 wire \u_cpu.REG_FILE._03649_ ;
 wire \u_cpu.REG_FILE._03650_ ;
 wire \u_cpu.REG_FILE._03651_ ;
 wire \u_cpu.REG_FILE._03652_ ;
 wire \u_cpu.REG_FILE._03653_ ;
 wire \u_cpu.REG_FILE._03654_ ;
 wire \u_cpu.REG_FILE._03655_ ;
 wire \u_cpu.REG_FILE._03656_ ;
 wire \u_cpu.REG_FILE._03657_ ;
 wire \u_cpu.REG_FILE._03658_ ;
 wire \u_cpu.REG_FILE._03659_ ;
 wire \u_cpu.REG_FILE._03660_ ;
 wire \u_cpu.REG_FILE._03661_ ;
 wire \u_cpu.REG_FILE._03662_ ;
 wire \u_cpu.REG_FILE._03663_ ;
 wire \u_cpu.REG_FILE._03664_ ;
 wire \u_cpu.REG_FILE._03665_ ;
 wire \u_cpu.REG_FILE._03666_ ;
 wire \u_cpu.REG_FILE._03667_ ;
 wire \u_cpu.REG_FILE._03668_ ;
 wire \u_cpu.REG_FILE._03669_ ;
 wire \u_cpu.REG_FILE._03670_ ;
 wire \u_cpu.REG_FILE._03671_ ;
 wire \u_cpu.REG_FILE._03672_ ;
 wire \u_cpu.REG_FILE._03673_ ;
 wire \u_cpu.REG_FILE._03674_ ;
 wire \u_cpu.REG_FILE._03675_ ;
 wire \u_cpu.REG_FILE._03676_ ;
 wire \u_cpu.REG_FILE._03677_ ;
 wire \u_cpu.REG_FILE._03678_ ;
 wire \u_cpu.REG_FILE._03679_ ;
 wire \u_cpu.REG_FILE._03680_ ;
 wire \u_cpu.REG_FILE._03681_ ;
 wire \u_cpu.REG_FILE._03682_ ;
 wire \u_cpu.REG_FILE._03683_ ;
 wire \u_cpu.REG_FILE._03684_ ;
 wire \u_cpu.REG_FILE._03685_ ;
 wire \u_cpu.REG_FILE._03686_ ;
 wire \u_cpu.REG_FILE._03687_ ;
 wire \u_cpu.REG_FILE._03688_ ;
 wire \u_cpu.REG_FILE._03689_ ;
 wire \u_cpu.REG_FILE._03690_ ;
 wire \u_cpu.REG_FILE._03691_ ;
 wire \u_cpu.REG_FILE._03692_ ;
 wire \u_cpu.REG_FILE._03693_ ;
 wire \u_cpu.REG_FILE._03694_ ;
 wire \u_cpu.REG_FILE._03695_ ;
 wire \u_cpu.REG_FILE._03696_ ;
 wire \u_cpu.REG_FILE._03697_ ;
 wire \u_cpu.REG_FILE._03698_ ;
 wire \u_cpu.REG_FILE._03699_ ;
 wire \u_cpu.REG_FILE._03700_ ;
 wire \u_cpu.REG_FILE._03701_ ;
 wire \u_cpu.REG_FILE._03702_ ;
 wire \u_cpu.REG_FILE._03703_ ;
 wire \u_cpu.REG_FILE._03704_ ;
 wire \u_cpu.REG_FILE._03705_ ;
 wire \u_cpu.REG_FILE._03706_ ;
 wire \u_cpu.REG_FILE._03707_ ;
 wire \u_cpu.REG_FILE._03708_ ;
 wire \u_cpu.REG_FILE._03709_ ;
 wire \u_cpu.REG_FILE._03710_ ;
 wire \u_cpu.REG_FILE._03711_ ;
 wire \u_cpu.REG_FILE._03712_ ;
 wire \u_cpu.REG_FILE._03713_ ;
 wire \u_cpu.REG_FILE._03714_ ;
 wire \u_cpu.REG_FILE._03715_ ;
 wire \u_cpu.REG_FILE._03716_ ;
 wire \u_cpu.REG_FILE._03717_ ;
 wire \u_cpu.REG_FILE._03718_ ;
 wire \u_cpu.REG_FILE._03719_ ;
 wire \u_cpu.REG_FILE._03720_ ;
 wire \u_cpu.REG_FILE._03721_ ;
 wire \u_cpu.REG_FILE._03722_ ;
 wire \u_cpu.REG_FILE._03723_ ;
 wire \u_cpu.REG_FILE._03724_ ;
 wire \u_cpu.REG_FILE._03725_ ;
 wire \u_cpu.REG_FILE._03726_ ;
 wire \u_cpu.REG_FILE._03727_ ;
 wire \u_cpu.REG_FILE._03728_ ;
 wire \u_cpu.REG_FILE._03729_ ;
 wire \u_cpu.REG_FILE._03730_ ;
 wire \u_cpu.REG_FILE._03731_ ;
 wire \u_cpu.REG_FILE._03732_ ;
 wire \u_cpu.REG_FILE._03733_ ;
 wire \u_cpu.REG_FILE._03734_ ;
 wire \u_cpu.REG_FILE._03735_ ;
 wire \u_cpu.REG_FILE._03736_ ;
 wire \u_cpu.REG_FILE._03737_ ;
 wire \u_cpu.REG_FILE._03738_ ;
 wire \u_cpu.REG_FILE._03739_ ;
 wire \u_cpu.REG_FILE._03740_ ;
 wire \u_cpu.REG_FILE._03741_ ;
 wire \u_cpu.REG_FILE._03742_ ;
 wire \u_cpu.REG_FILE._03743_ ;
 wire \u_cpu.REG_FILE._03744_ ;
 wire \u_cpu.REG_FILE._03745_ ;
 wire \u_cpu.REG_FILE._03746_ ;
 wire \u_cpu.REG_FILE._03747_ ;
 wire \u_cpu.REG_FILE._03748_ ;
 wire \u_cpu.REG_FILE._03749_ ;
 wire \u_cpu.REG_FILE._03750_ ;
 wire \u_cpu.REG_FILE._03751_ ;
 wire \u_cpu.REG_FILE._03752_ ;
 wire \u_cpu.REG_FILE._03753_ ;
 wire \u_cpu.REG_FILE._03754_ ;
 wire \u_cpu.REG_FILE._03755_ ;
 wire \u_cpu.REG_FILE._03756_ ;
 wire \u_cpu.REG_FILE._03757_ ;
 wire \u_cpu.REG_FILE._03758_ ;
 wire \u_cpu.REG_FILE._03759_ ;
 wire \u_cpu.REG_FILE._03760_ ;
 wire \u_cpu.REG_FILE._03761_ ;
 wire \u_cpu.REG_FILE._03762_ ;
 wire \u_cpu.REG_FILE._03763_ ;
 wire \u_cpu.REG_FILE._03764_ ;
 wire \u_cpu.REG_FILE._03765_ ;
 wire \u_cpu.REG_FILE._03766_ ;
 wire \u_cpu.REG_FILE._03767_ ;
 wire \u_cpu.REG_FILE._03768_ ;
 wire \u_cpu.REG_FILE._03769_ ;
 wire \u_cpu.REG_FILE._03770_ ;
 wire \u_cpu.REG_FILE._03771_ ;
 wire \u_cpu.REG_FILE._03772_ ;
 wire \u_cpu.REG_FILE._03773_ ;
 wire \u_cpu.REG_FILE._03774_ ;
 wire \u_cpu.REG_FILE._03775_ ;
 wire \u_cpu.REG_FILE._03776_ ;
 wire \u_cpu.REG_FILE._03777_ ;
 wire \u_cpu.REG_FILE._03778_ ;
 wire \u_cpu.REG_FILE._03779_ ;
 wire \u_cpu.REG_FILE._03780_ ;
 wire \u_cpu.REG_FILE._03781_ ;
 wire \u_cpu.REG_FILE._03782_ ;
 wire \u_cpu.REG_FILE._03783_ ;
 wire \u_cpu.REG_FILE._03784_ ;
 wire \u_cpu.REG_FILE._03785_ ;
 wire \u_cpu.REG_FILE._03786_ ;
 wire \u_cpu.REG_FILE._03787_ ;
 wire \u_cpu.REG_FILE._03788_ ;
 wire \u_cpu.REG_FILE._03789_ ;
 wire \u_cpu.REG_FILE._03790_ ;
 wire \u_cpu.REG_FILE._03791_ ;
 wire \u_cpu.REG_FILE._03792_ ;
 wire \u_cpu.REG_FILE._03793_ ;
 wire \u_cpu.REG_FILE._03794_ ;
 wire \u_cpu.REG_FILE._03795_ ;
 wire \u_cpu.REG_FILE._03796_ ;
 wire \u_cpu.REG_FILE._03797_ ;
 wire \u_cpu.REG_FILE._03798_ ;
 wire \u_cpu.REG_FILE._03799_ ;
 wire \u_cpu.REG_FILE._03800_ ;
 wire \u_cpu.REG_FILE._03801_ ;
 wire \u_cpu.REG_FILE._03802_ ;
 wire \u_cpu.REG_FILE._03803_ ;
 wire \u_cpu.REG_FILE._03804_ ;
 wire \u_cpu.REG_FILE._03805_ ;
 wire \u_cpu.REG_FILE._03806_ ;
 wire \u_cpu.REG_FILE._03807_ ;
 wire \u_cpu.REG_FILE._03808_ ;
 wire \u_cpu.REG_FILE._03809_ ;
 wire \u_cpu.REG_FILE._03810_ ;
 wire \u_cpu.REG_FILE._03811_ ;
 wire \u_cpu.REG_FILE._03812_ ;
 wire \u_cpu.REG_FILE._03813_ ;
 wire \u_cpu.REG_FILE._03814_ ;
 wire \u_cpu.REG_FILE._03815_ ;
 wire \u_cpu.REG_FILE._03816_ ;
 wire \u_cpu.REG_FILE._03817_ ;
 wire \u_cpu.REG_FILE._03818_ ;
 wire \u_cpu.REG_FILE._03819_ ;
 wire \u_cpu.REG_FILE._03820_ ;
 wire \u_cpu.REG_FILE._03821_ ;
 wire \u_cpu.REG_FILE._03822_ ;
 wire \u_cpu.REG_FILE._03823_ ;
 wire \u_cpu.REG_FILE._03824_ ;
 wire \u_cpu.REG_FILE._03825_ ;
 wire \u_cpu.REG_FILE._03826_ ;
 wire \u_cpu.REG_FILE._03827_ ;
 wire \u_cpu.REG_FILE._03828_ ;
 wire \u_cpu.REG_FILE._03829_ ;
 wire \u_cpu.REG_FILE._03830_ ;
 wire \u_cpu.REG_FILE._03831_ ;
 wire \u_cpu.REG_FILE._03832_ ;
 wire \u_cpu.REG_FILE._03833_ ;
 wire \u_cpu.REG_FILE._03834_ ;
 wire \u_cpu.REG_FILE._03835_ ;
 wire \u_cpu.REG_FILE._03836_ ;
 wire \u_cpu.REG_FILE._03837_ ;
 wire \u_cpu.REG_FILE._03838_ ;
 wire \u_cpu.REG_FILE._03839_ ;
 wire \u_cpu.REG_FILE._03840_ ;
 wire \u_cpu.REG_FILE._03841_ ;
 wire \u_cpu.REG_FILE._03842_ ;
 wire \u_cpu.REG_FILE._03843_ ;
 wire \u_cpu.REG_FILE._03844_ ;
 wire \u_cpu.REG_FILE._03845_ ;
 wire \u_cpu.REG_FILE._03846_ ;
 wire \u_cpu.REG_FILE._03847_ ;
 wire \u_cpu.REG_FILE._03848_ ;
 wire \u_cpu.REG_FILE._03849_ ;
 wire \u_cpu.REG_FILE._03850_ ;
 wire \u_cpu.REG_FILE._03851_ ;
 wire \u_cpu.REG_FILE._03852_ ;
 wire \u_cpu.REG_FILE._03853_ ;
 wire \u_cpu.REG_FILE._03854_ ;
 wire \u_cpu.REG_FILE._03855_ ;
 wire \u_cpu.REG_FILE._03856_ ;
 wire \u_cpu.REG_FILE._03857_ ;
 wire \u_cpu.REG_FILE._03858_ ;
 wire \u_cpu.REG_FILE._03859_ ;
 wire \u_cpu.REG_FILE._03860_ ;
 wire \u_cpu.REG_FILE._03861_ ;
 wire \u_cpu.REG_FILE._03862_ ;
 wire \u_cpu.REG_FILE._03863_ ;
 wire \u_cpu.REG_FILE._03864_ ;
 wire \u_cpu.REG_FILE._03865_ ;
 wire \u_cpu.REG_FILE._03866_ ;
 wire \u_cpu.REG_FILE._03867_ ;
 wire \u_cpu.REG_FILE._03868_ ;
 wire \u_cpu.REG_FILE._03869_ ;
 wire \u_cpu.REG_FILE._03870_ ;
 wire \u_cpu.REG_FILE._03871_ ;
 wire \u_cpu.REG_FILE._03872_ ;
 wire \u_cpu.REG_FILE._03873_ ;
 wire \u_cpu.REG_FILE._03874_ ;
 wire \u_cpu.REG_FILE._03875_ ;
 wire \u_cpu.REG_FILE._03876_ ;
 wire \u_cpu.REG_FILE._03877_ ;
 wire \u_cpu.REG_FILE._03878_ ;
 wire \u_cpu.REG_FILE._03879_ ;
 wire \u_cpu.REG_FILE._03880_ ;
 wire \u_cpu.REG_FILE._03881_ ;
 wire \u_cpu.REG_FILE._03882_ ;
 wire \u_cpu.REG_FILE._03883_ ;
 wire \u_cpu.REG_FILE._03884_ ;
 wire \u_cpu.REG_FILE._03885_ ;
 wire \u_cpu.REG_FILE._03886_ ;
 wire \u_cpu.REG_FILE._03887_ ;
 wire \u_cpu.REG_FILE._03888_ ;
 wire \u_cpu.REG_FILE._03889_ ;
 wire \u_cpu.REG_FILE._03890_ ;
 wire \u_cpu.REG_FILE._03891_ ;
 wire \u_cpu.REG_FILE._03892_ ;
 wire \u_cpu.REG_FILE._03893_ ;
 wire \u_cpu.REG_FILE._03894_ ;
 wire \u_cpu.REG_FILE._03895_ ;
 wire \u_cpu.REG_FILE._03896_ ;
 wire \u_cpu.REG_FILE._03897_ ;
 wire \u_cpu.REG_FILE._03898_ ;
 wire \u_cpu.REG_FILE._03899_ ;
 wire \u_cpu.REG_FILE._03900_ ;
 wire \u_cpu.REG_FILE._03901_ ;
 wire \u_cpu.REG_FILE._03902_ ;
 wire \u_cpu.REG_FILE._03903_ ;
 wire \u_cpu.REG_FILE._03904_ ;
 wire \u_cpu.REG_FILE._03905_ ;
 wire \u_cpu.REG_FILE._03906_ ;
 wire \u_cpu.REG_FILE._03907_ ;
 wire \u_cpu.REG_FILE._03908_ ;
 wire \u_cpu.REG_FILE._03909_ ;
 wire \u_cpu.REG_FILE._03910_ ;
 wire \u_cpu.REG_FILE._03911_ ;
 wire \u_cpu.REG_FILE._03912_ ;
 wire \u_cpu.REG_FILE._03913_ ;
 wire \u_cpu.REG_FILE._03914_ ;
 wire \u_cpu.REG_FILE._03915_ ;
 wire \u_cpu.REG_FILE._03916_ ;
 wire \u_cpu.REG_FILE._03917_ ;
 wire \u_cpu.REG_FILE._03918_ ;
 wire \u_cpu.REG_FILE._03919_ ;
 wire \u_cpu.REG_FILE._03920_ ;
 wire \u_cpu.REG_FILE._03921_ ;
 wire \u_cpu.REG_FILE._03922_ ;
 wire \u_cpu.REG_FILE._03923_ ;
 wire \u_cpu.REG_FILE._03924_ ;
 wire \u_cpu.REG_FILE._03925_ ;
 wire \u_cpu.REG_FILE._03926_ ;
 wire \u_cpu.REG_FILE._03927_ ;
 wire \u_cpu.REG_FILE._03928_ ;
 wire \u_cpu.REG_FILE._03929_ ;
 wire \u_cpu.REG_FILE._03930_ ;
 wire \u_cpu.REG_FILE._03931_ ;
 wire \u_cpu.REG_FILE._03932_ ;
 wire \u_cpu.REG_FILE._03933_ ;
 wire \u_cpu.REG_FILE._03934_ ;
 wire \u_cpu.REG_FILE._03935_ ;
 wire \u_cpu.REG_FILE._03936_ ;
 wire \u_cpu.REG_FILE._03937_ ;
 wire \u_cpu.REG_FILE._03938_ ;
 wire \u_cpu.REG_FILE._03939_ ;
 wire \u_cpu.REG_FILE._03940_ ;
 wire \u_cpu.REG_FILE._03941_ ;
 wire \u_cpu.REG_FILE._03942_ ;
 wire \u_cpu.REG_FILE._03943_ ;
 wire \u_cpu.REG_FILE._03944_ ;
 wire \u_cpu.REG_FILE._03945_ ;
 wire \u_cpu.REG_FILE._03946_ ;
 wire \u_cpu.REG_FILE._03947_ ;
 wire \u_cpu.REG_FILE._03948_ ;
 wire \u_cpu.REG_FILE._03949_ ;
 wire \u_cpu.REG_FILE._03950_ ;
 wire \u_cpu.REG_FILE._03951_ ;
 wire \u_cpu.REG_FILE._03952_ ;
 wire \u_cpu.REG_FILE._03953_ ;
 wire \u_cpu.REG_FILE._03954_ ;
 wire \u_cpu.REG_FILE._03955_ ;
 wire \u_cpu.REG_FILE._03956_ ;
 wire \u_cpu.REG_FILE._03957_ ;
 wire \u_cpu.REG_FILE._03958_ ;
 wire \u_cpu.REG_FILE._03959_ ;
 wire \u_cpu.REG_FILE._03960_ ;
 wire \u_cpu.REG_FILE._03961_ ;
 wire \u_cpu.REG_FILE._03962_ ;
 wire \u_cpu.REG_FILE._03963_ ;
 wire \u_cpu.REG_FILE._03964_ ;
 wire \u_cpu.REG_FILE._03965_ ;
 wire \u_cpu.REG_FILE._03966_ ;
 wire \u_cpu.REG_FILE._03967_ ;
 wire \u_cpu.REG_FILE._03968_ ;
 wire \u_cpu.REG_FILE._03969_ ;
 wire \u_cpu.REG_FILE._03970_ ;
 wire \u_cpu.REG_FILE._03971_ ;
 wire \u_cpu.REG_FILE._03972_ ;
 wire \u_cpu.REG_FILE._03973_ ;
 wire \u_cpu.REG_FILE._03974_ ;
 wire \u_cpu.REG_FILE._03975_ ;
 wire \u_cpu.REG_FILE._03976_ ;
 wire \u_cpu.REG_FILE._03977_ ;
 wire \u_cpu.REG_FILE._03978_ ;
 wire \u_cpu.REG_FILE._03979_ ;
 wire \u_cpu.REG_FILE._03980_ ;
 wire \u_cpu.REG_FILE._03981_ ;
 wire \u_cpu.REG_FILE._03982_ ;
 wire \u_cpu.REG_FILE._03983_ ;
 wire \u_cpu.REG_FILE._03984_ ;
 wire \u_cpu.REG_FILE._03985_ ;
 wire \u_cpu.REG_FILE._03986_ ;
 wire \u_cpu.REG_FILE._03987_ ;
 wire \u_cpu.REG_FILE._03988_ ;
 wire \u_cpu.REG_FILE._03989_ ;
 wire \u_cpu.REG_FILE._03990_ ;
 wire \u_cpu.REG_FILE._03991_ ;
 wire \u_cpu.REG_FILE._03992_ ;
 wire \u_cpu.REG_FILE._03993_ ;
 wire \u_cpu.REG_FILE._03994_ ;
 wire \u_cpu.REG_FILE._03995_ ;
 wire \u_cpu.REG_FILE._03996_ ;
 wire \u_cpu.REG_FILE._03997_ ;
 wire \u_cpu.REG_FILE._03998_ ;
 wire \u_cpu.REG_FILE._03999_ ;
 wire \u_cpu.REG_FILE._04000_ ;
 wire \u_cpu.REG_FILE._04001_ ;
 wire \u_cpu.REG_FILE._04002_ ;
 wire \u_cpu.REG_FILE._04003_ ;
 wire \u_cpu.REG_FILE._04004_ ;
 wire \u_cpu.REG_FILE._04005_ ;
 wire \u_cpu.REG_FILE._04006_ ;
 wire \u_cpu.REG_FILE._04007_ ;
 wire \u_cpu.REG_FILE._04008_ ;
 wire \u_cpu.REG_FILE._04009_ ;
 wire \u_cpu.REG_FILE._04010_ ;
 wire \u_cpu.REG_FILE._04011_ ;
 wire \u_cpu.REG_FILE._04012_ ;
 wire \u_cpu.REG_FILE._04013_ ;
 wire \u_cpu.REG_FILE._04014_ ;
 wire \u_cpu.REG_FILE._04015_ ;
 wire \u_cpu.REG_FILE._04016_ ;
 wire \u_cpu.REG_FILE._04017_ ;
 wire \u_cpu.REG_FILE._04018_ ;
 wire \u_cpu.REG_FILE._04019_ ;
 wire \u_cpu.REG_FILE._04020_ ;
 wire \u_cpu.REG_FILE._04021_ ;
 wire \u_cpu.REG_FILE._04022_ ;
 wire \u_cpu.REG_FILE._04023_ ;
 wire \u_cpu.REG_FILE._04024_ ;
 wire \u_cpu.REG_FILE._04025_ ;
 wire \u_cpu.REG_FILE._04026_ ;
 wire \u_cpu.REG_FILE._04027_ ;
 wire \u_cpu.REG_FILE._04028_ ;
 wire \u_cpu.REG_FILE._04029_ ;
 wire \u_cpu.REG_FILE._04030_ ;
 wire \u_cpu.REG_FILE._04031_ ;
 wire \u_cpu.REG_FILE._04032_ ;
 wire \u_cpu.REG_FILE._04033_ ;
 wire \u_cpu.REG_FILE._04034_ ;
 wire \u_cpu.REG_FILE._04035_ ;
 wire \u_cpu.REG_FILE._04036_ ;
 wire \u_cpu.REG_FILE._04037_ ;
 wire \u_cpu.REG_FILE._04038_ ;
 wire \u_cpu.REG_FILE._04039_ ;
 wire \u_cpu.REG_FILE._04040_ ;
 wire \u_cpu.REG_FILE._04041_ ;
 wire \u_cpu.REG_FILE._04042_ ;
 wire \u_cpu.REG_FILE._04043_ ;
 wire \u_cpu.REG_FILE._04044_ ;
 wire \u_cpu.REG_FILE._04045_ ;
 wire \u_cpu.REG_FILE._04046_ ;
 wire \u_cpu.REG_FILE._04047_ ;
 wire \u_cpu.REG_FILE._04048_ ;
 wire \u_cpu.REG_FILE._04049_ ;
 wire \u_cpu.REG_FILE._04050_ ;
 wire \u_cpu.REG_FILE._04051_ ;
 wire \u_cpu.REG_FILE._04052_ ;
 wire \u_cpu.REG_FILE._04053_ ;
 wire \u_cpu.REG_FILE._04054_ ;
 wire \u_cpu.REG_FILE._04055_ ;
 wire \u_cpu.REG_FILE._04056_ ;
 wire \u_cpu.REG_FILE._04057_ ;
 wire \u_cpu.REG_FILE._04058_ ;
 wire \u_cpu.REG_FILE._04059_ ;
 wire \u_cpu.REG_FILE._04060_ ;
 wire \u_cpu.REG_FILE._04061_ ;
 wire \u_cpu.REG_FILE._04062_ ;
 wire \u_cpu.REG_FILE._04063_ ;
 wire \u_cpu.REG_FILE._04064_ ;
 wire \u_cpu.REG_FILE._04065_ ;
 wire \u_cpu.REG_FILE._04066_ ;
 wire \u_cpu.REG_FILE._04067_ ;
 wire \u_cpu.REG_FILE._04068_ ;
 wire \u_cpu.REG_FILE._04069_ ;
 wire \u_cpu.REG_FILE._04070_ ;
 wire \u_cpu.REG_FILE._04071_ ;
 wire \u_cpu.REG_FILE._04072_ ;
 wire \u_cpu.REG_FILE._04073_ ;
 wire \u_cpu.REG_FILE._04074_ ;
 wire \u_cpu.REG_FILE._04075_ ;
 wire \u_cpu.REG_FILE._04076_ ;
 wire \u_cpu.REG_FILE._04077_ ;
 wire \u_cpu.REG_FILE._04078_ ;
 wire \u_cpu.REG_FILE._04079_ ;
 wire \u_cpu.REG_FILE._04080_ ;
 wire \u_cpu.REG_FILE._04081_ ;
 wire \u_cpu.REG_FILE._04082_ ;
 wire \u_cpu.REG_FILE._04083_ ;
 wire \u_cpu.REG_FILE._04084_ ;
 wire \u_cpu.REG_FILE._04085_ ;
 wire \u_cpu.REG_FILE._04086_ ;
 wire \u_cpu.REG_FILE._04087_ ;
 wire \u_cpu.REG_FILE._04088_ ;
 wire \u_cpu.REG_FILE._04089_ ;
 wire \u_cpu.REG_FILE._04090_ ;
 wire \u_cpu.REG_FILE._04091_ ;
 wire \u_cpu.REG_FILE._04092_ ;
 wire \u_cpu.REG_FILE._04093_ ;
 wire \u_cpu.REG_FILE._04094_ ;
 wire \u_cpu.REG_FILE._04095_ ;
 wire \u_cpu.REG_FILE._04096_ ;
 wire \u_cpu.REG_FILE._04097_ ;
 wire \u_cpu.REG_FILE._04098_ ;
 wire \u_cpu.REG_FILE._04099_ ;
 wire \u_cpu.REG_FILE._04100_ ;
 wire \u_cpu.REG_FILE._04101_ ;
 wire \u_cpu.REG_FILE._04102_ ;
 wire \u_cpu.REG_FILE._04103_ ;
 wire \u_cpu.REG_FILE._04104_ ;
 wire \u_cpu.REG_FILE._04105_ ;
 wire \u_cpu.REG_FILE._04106_ ;
 wire \u_cpu.REG_FILE._04107_ ;
 wire \u_cpu.REG_FILE._04108_ ;
 wire \u_cpu.REG_FILE._04109_ ;
 wire \u_cpu.REG_FILE._04110_ ;
 wire \u_cpu.REG_FILE._04111_ ;
 wire \u_cpu.REG_FILE._04112_ ;
 wire \u_cpu.REG_FILE._04113_ ;
 wire \u_cpu.REG_FILE._04114_ ;
 wire \u_cpu.REG_FILE._04115_ ;
 wire \u_cpu.REG_FILE._04116_ ;
 wire \u_cpu.REG_FILE._04117_ ;
 wire \u_cpu.REG_FILE._04118_ ;
 wire \u_cpu.REG_FILE._04119_ ;
 wire \u_cpu.REG_FILE._04120_ ;
 wire \u_cpu.REG_FILE._04121_ ;
 wire \u_cpu.REG_FILE._04122_ ;
 wire \u_cpu.REG_FILE._04123_ ;
 wire \u_cpu.REG_FILE._04124_ ;
 wire \u_cpu.REG_FILE._04125_ ;
 wire \u_cpu.REG_FILE._04126_ ;
 wire \u_cpu.REG_FILE._04127_ ;
 wire \u_cpu.REG_FILE._04128_ ;
 wire \u_cpu.REG_FILE._04129_ ;
 wire \u_cpu.REG_FILE._04130_ ;
 wire \u_cpu.REG_FILE._04131_ ;
 wire \u_cpu.REG_FILE._04132_ ;
 wire \u_cpu.REG_FILE._04133_ ;
 wire \u_cpu.REG_FILE._04134_ ;
 wire \u_cpu.REG_FILE._04135_ ;
 wire \u_cpu.REG_FILE._04136_ ;
 wire \u_cpu.REG_FILE._04137_ ;
 wire \u_cpu.REG_FILE._04138_ ;
 wire \u_cpu.REG_FILE._04139_ ;
 wire \u_cpu.REG_FILE._04140_ ;
 wire \u_cpu.REG_FILE._04141_ ;
 wire \u_cpu.REG_FILE._04142_ ;
 wire \u_cpu.REG_FILE._04143_ ;
 wire \u_cpu.REG_FILE._04144_ ;
 wire \u_cpu.REG_FILE._04145_ ;
 wire \u_cpu.REG_FILE._04146_ ;
 wire \u_cpu.REG_FILE._04147_ ;
 wire \u_cpu.REG_FILE._04148_ ;
 wire \u_cpu.REG_FILE._04149_ ;
 wire \u_cpu.REG_FILE._04150_ ;
 wire \u_cpu.REG_FILE._04151_ ;
 wire \u_cpu.REG_FILE._04152_ ;
 wire \u_cpu.REG_FILE._04153_ ;
 wire \u_cpu.REG_FILE._04154_ ;
 wire \u_cpu.REG_FILE._04155_ ;
 wire \u_cpu.REG_FILE._04156_ ;
 wire \u_cpu.REG_FILE._04157_ ;
 wire \u_cpu.REG_FILE._04158_ ;
 wire \u_cpu.REG_FILE._04159_ ;
 wire \u_cpu.REG_FILE._04160_ ;
 wire \u_cpu.REG_FILE._04161_ ;
 wire \u_cpu.REG_FILE._04162_ ;
 wire \u_cpu.REG_FILE._04163_ ;
 wire \u_cpu.REG_FILE._04164_ ;
 wire \u_cpu.REG_FILE._04165_ ;
 wire \u_cpu.REG_FILE._04166_ ;
 wire \u_cpu.REG_FILE._04167_ ;
 wire \u_cpu.REG_FILE._04168_ ;
 wire \u_cpu.REG_FILE._04169_ ;
 wire \u_cpu.REG_FILE._04170_ ;
 wire \u_cpu.REG_FILE._04171_ ;
 wire \u_cpu.REG_FILE._04172_ ;
 wire \u_cpu.REG_FILE._04173_ ;
 wire \u_cpu.REG_FILE._04174_ ;
 wire \u_cpu.REG_FILE._04175_ ;
 wire \u_cpu.REG_FILE._04176_ ;
 wire \u_cpu.REG_FILE._04177_ ;
 wire \u_cpu.REG_FILE._04178_ ;
 wire \u_cpu.REG_FILE._04179_ ;
 wire \u_cpu.REG_FILE._04180_ ;
 wire \u_cpu.REG_FILE._04181_ ;
 wire \u_cpu.REG_FILE._04182_ ;
 wire \u_cpu.REG_FILE._04183_ ;
 wire \u_cpu.REG_FILE._04184_ ;
 wire \u_cpu.REG_FILE._04185_ ;
 wire \u_cpu.REG_FILE._04186_ ;
 wire \u_cpu.REG_FILE._04187_ ;
 wire \u_cpu.REG_FILE._04188_ ;
 wire \u_cpu.REG_FILE._04189_ ;
 wire \u_cpu.REG_FILE._04190_ ;
 wire \u_cpu.REG_FILE._04191_ ;
 wire \u_cpu.REG_FILE._04192_ ;
 wire \u_cpu.REG_FILE._04193_ ;
 wire \u_cpu.REG_FILE._04194_ ;
 wire \u_cpu.REG_FILE._04195_ ;
 wire \u_cpu.REG_FILE._04196_ ;
 wire \u_cpu.REG_FILE._04197_ ;
 wire \u_cpu.REG_FILE._04198_ ;
 wire \u_cpu.REG_FILE._04199_ ;
 wire \u_cpu.REG_FILE._04200_ ;
 wire \u_cpu.REG_FILE._04201_ ;
 wire \u_cpu.REG_FILE._04202_ ;
 wire \u_cpu.REG_FILE._04203_ ;
 wire \u_cpu.REG_FILE._04204_ ;
 wire \u_cpu.REG_FILE._04205_ ;
 wire \u_cpu.REG_FILE._04206_ ;
 wire \u_cpu.REG_FILE._04207_ ;
 wire \u_cpu.REG_FILE._04208_ ;
 wire \u_cpu.REG_FILE._04209_ ;
 wire \u_cpu.REG_FILE._04210_ ;
 wire \u_cpu.REG_FILE._04211_ ;
 wire \u_cpu.REG_FILE._04212_ ;
 wire \u_cpu.REG_FILE._04213_ ;
 wire \u_cpu.REG_FILE._04214_ ;
 wire \u_cpu.REG_FILE._04215_ ;
 wire \u_cpu.REG_FILE._04216_ ;
 wire \u_cpu.REG_FILE._04217_ ;
 wire \u_cpu.REG_FILE._04218_ ;
 wire \u_cpu.REG_FILE._04219_ ;
 wire \u_cpu.REG_FILE._04220_ ;
 wire \u_cpu.REG_FILE._04221_ ;
 wire \u_cpu.REG_FILE._04222_ ;
 wire \u_cpu.REG_FILE._04223_ ;
 wire \u_cpu.REG_FILE._04224_ ;
 wire \u_cpu.REG_FILE._04225_ ;
 wire \u_cpu.REG_FILE._04226_ ;
 wire \u_cpu.REG_FILE._04227_ ;
 wire \u_cpu.REG_FILE._04228_ ;
 wire \u_cpu.REG_FILE._04229_ ;
 wire \u_cpu.REG_FILE._04230_ ;
 wire \u_cpu.REG_FILE._04231_ ;
 wire \u_cpu.REG_FILE._04232_ ;
 wire \u_cpu.REG_FILE._04233_ ;
 wire \u_cpu.REG_FILE._04234_ ;
 wire \u_cpu.REG_FILE._04235_ ;
 wire \u_cpu.REG_FILE._04236_ ;
 wire \u_cpu.REG_FILE._04237_ ;
 wire \u_cpu.REG_FILE._04238_ ;
 wire \u_cpu.REG_FILE._04239_ ;
 wire \u_cpu.REG_FILE._04240_ ;
 wire \u_cpu.REG_FILE._04241_ ;
 wire \u_cpu.REG_FILE._04242_ ;
 wire \u_cpu.REG_FILE._04243_ ;
 wire \u_cpu.REG_FILE._04244_ ;
 wire \u_cpu.REG_FILE._04245_ ;
 wire \u_cpu.REG_FILE._04246_ ;
 wire \u_cpu.REG_FILE._04247_ ;
 wire \u_cpu.REG_FILE._04248_ ;
 wire \u_cpu.REG_FILE._04249_ ;
 wire \u_cpu.REG_FILE._04250_ ;
 wire \u_cpu.REG_FILE._04251_ ;
 wire \u_cpu.REG_FILE._04252_ ;
 wire \u_cpu.REG_FILE._04253_ ;
 wire \u_cpu.REG_FILE._04254_ ;
 wire \u_cpu.REG_FILE._04255_ ;
 wire \u_cpu.REG_FILE._04256_ ;
 wire \u_cpu.REG_FILE._04257_ ;
 wire \u_cpu.REG_FILE._04258_ ;
 wire \u_cpu.REG_FILE._04259_ ;
 wire \u_cpu.REG_FILE._04260_ ;
 wire \u_cpu.REG_FILE._04261_ ;
 wire \u_cpu.REG_FILE._04262_ ;
 wire \u_cpu.REG_FILE._04263_ ;
 wire \u_cpu.REG_FILE._04264_ ;
 wire \u_cpu.REG_FILE._04265_ ;
 wire \u_cpu.REG_FILE._04266_ ;
 wire \u_cpu.REG_FILE._04267_ ;
 wire \u_cpu.REG_FILE._04268_ ;
 wire \u_cpu.REG_FILE._04269_ ;
 wire \u_cpu.REG_FILE._04270_ ;
 wire \u_cpu.REG_FILE._04271_ ;
 wire \u_cpu.REG_FILE._04272_ ;
 wire \u_cpu.REG_FILE._04273_ ;
 wire \u_cpu.REG_FILE._04274_ ;
 wire \u_cpu.REG_FILE._04275_ ;
 wire \u_cpu.REG_FILE._04276_ ;
 wire \u_cpu.REG_FILE._04277_ ;
 wire \u_cpu.REG_FILE._04278_ ;
 wire \u_cpu.REG_FILE._04279_ ;
 wire \u_cpu.REG_FILE._04280_ ;
 wire \u_cpu.REG_FILE._04281_ ;
 wire \u_cpu.REG_FILE._04282_ ;
 wire \u_cpu.REG_FILE._04283_ ;
 wire \u_cpu.REG_FILE._04284_ ;
 wire \u_cpu.REG_FILE._04285_ ;
 wire \u_cpu.REG_FILE._04286_ ;
 wire \u_cpu.REG_FILE._04287_ ;
 wire \u_cpu.REG_FILE._04288_ ;
 wire \u_cpu.REG_FILE._04289_ ;
 wire \u_cpu.REG_FILE._04290_ ;
 wire \u_cpu.REG_FILE._04291_ ;
 wire \u_cpu.REG_FILE._04292_ ;
 wire \u_cpu.REG_FILE._04293_ ;
 wire \u_cpu.REG_FILE._04294_ ;
 wire \u_cpu.REG_FILE._04295_ ;
 wire \u_cpu.REG_FILE._04296_ ;
 wire \u_cpu.REG_FILE._04297_ ;
 wire \u_cpu.REG_FILE._04298_ ;
 wire \u_cpu.REG_FILE._04299_ ;
 wire \u_cpu.REG_FILE._04300_ ;
 wire \u_cpu.REG_FILE._04301_ ;
 wire \u_cpu.REG_FILE._04302_ ;
 wire \u_cpu.REG_FILE._04303_ ;
 wire \u_cpu.REG_FILE._04304_ ;
 wire \u_cpu.REG_FILE._04305_ ;
 wire \u_cpu.REG_FILE._04306_ ;
 wire \u_cpu.REG_FILE._04307_ ;
 wire \u_cpu.REG_FILE._04308_ ;
 wire \u_cpu.REG_FILE._04309_ ;
 wire \u_cpu.REG_FILE._04310_ ;
 wire \u_cpu.REG_FILE._04311_ ;
 wire \u_cpu.REG_FILE._04312_ ;
 wire \u_cpu.REG_FILE._04313_ ;
 wire \u_cpu.REG_FILE._04314_ ;
 wire \u_cpu.REG_FILE._04315_ ;
 wire \u_cpu.REG_FILE._04316_ ;
 wire \u_cpu.REG_FILE._04317_ ;
 wire \u_cpu.REG_FILE._04318_ ;
 wire \u_cpu.REG_FILE._04319_ ;
 wire \u_cpu.REG_FILE._04320_ ;
 wire \u_cpu.REG_FILE._04321_ ;
 wire \u_cpu.REG_FILE._04322_ ;
 wire \u_cpu.REG_FILE._04323_ ;
 wire \u_cpu.REG_FILE._04324_ ;
 wire \u_cpu.REG_FILE._04325_ ;
 wire \u_cpu.REG_FILE._04326_ ;
 wire \u_cpu.REG_FILE._04327_ ;
 wire \u_cpu.REG_FILE._04328_ ;
 wire \u_cpu.REG_FILE._04329_ ;
 wire \u_cpu.REG_FILE._04330_ ;
 wire \u_cpu.REG_FILE._04331_ ;
 wire \u_cpu.REG_FILE._04332_ ;
 wire \u_cpu.REG_FILE._04333_ ;
 wire \u_cpu.REG_FILE._04334_ ;
 wire \u_cpu.REG_FILE._04335_ ;
 wire \u_cpu.REG_FILE._04336_ ;
 wire \u_cpu.REG_FILE._04337_ ;
 wire \u_cpu.REG_FILE._04338_ ;
 wire \u_cpu.REG_FILE._04339_ ;
 wire \u_cpu.REG_FILE._04340_ ;
 wire \u_cpu.REG_FILE._04341_ ;
 wire \u_cpu.REG_FILE._04342_ ;
 wire \u_cpu.REG_FILE._04343_ ;
 wire \u_cpu.REG_FILE._04344_ ;
 wire \u_cpu.REG_FILE._04345_ ;
 wire \u_cpu.REG_FILE._04346_ ;
 wire \u_cpu.REG_FILE._04347_ ;
 wire \u_cpu.REG_FILE._04348_ ;
 wire \u_cpu.REG_FILE._04349_ ;
 wire \u_cpu.REG_FILE._04350_ ;
 wire \u_cpu.REG_FILE._04351_ ;
 wire \u_cpu.REG_FILE._04352_ ;
 wire \u_cpu.REG_FILE._04353_ ;
 wire \u_cpu.REG_FILE._04354_ ;
 wire \u_cpu.REG_FILE._04355_ ;
 wire \u_cpu.REG_FILE._04356_ ;
 wire \u_cpu.REG_FILE._04357_ ;
 wire \u_cpu.REG_FILE._04358_ ;
 wire \u_cpu.REG_FILE._04359_ ;
 wire \u_cpu.REG_FILE._04360_ ;
 wire \u_cpu.REG_FILE._04361_ ;
 wire \u_cpu.REG_FILE._04362_ ;
 wire \u_cpu.REG_FILE._04363_ ;
 wire \u_cpu.REG_FILE._04364_ ;
 wire \u_cpu.REG_FILE._04365_ ;
 wire \u_cpu.REG_FILE._04366_ ;
 wire \u_cpu.REG_FILE._04367_ ;
 wire \u_cpu.REG_FILE._04368_ ;
 wire \u_cpu.REG_FILE._04369_ ;
 wire \u_cpu.REG_FILE._04370_ ;
 wire \u_cpu.REG_FILE._04371_ ;
 wire \u_cpu.REG_FILE._04372_ ;
 wire \u_cpu.REG_FILE._04373_ ;
 wire \u_cpu.REG_FILE._04374_ ;
 wire \u_cpu.REG_FILE._04375_ ;
 wire \u_cpu.REG_FILE._04376_ ;
 wire \u_cpu.REG_FILE._04377_ ;
 wire \u_cpu.REG_FILE._04378_ ;
 wire \u_cpu.REG_FILE._04379_ ;
 wire \u_cpu.REG_FILE._04380_ ;
 wire \u_cpu.REG_FILE._04381_ ;
 wire \u_cpu.REG_FILE._04382_ ;
 wire \u_cpu.REG_FILE._04383_ ;
 wire \u_cpu.REG_FILE._04384_ ;
 wire \u_cpu.REG_FILE._04385_ ;
 wire \u_cpu.REG_FILE._04386_ ;
 wire \u_cpu.REG_FILE._04387_ ;
 wire \u_cpu.REG_FILE._04388_ ;
 wire \u_cpu.REG_FILE._04389_ ;
 wire \u_cpu.REG_FILE._04390_ ;
 wire \u_cpu.REG_FILE._04391_ ;
 wire \u_cpu.REG_FILE._04392_ ;
 wire \u_cpu.REG_FILE._04393_ ;
 wire \u_cpu.REG_FILE._04394_ ;
 wire \u_cpu.REG_FILE._04395_ ;
 wire \u_cpu.REG_FILE._04396_ ;
 wire \u_cpu.REG_FILE._04397_ ;
 wire \u_cpu.REG_FILE._04398_ ;
 wire \u_cpu.REG_FILE._04399_ ;
 wire \u_cpu.REG_FILE._04400_ ;
 wire \u_cpu.REG_FILE._04401_ ;
 wire \u_cpu.REG_FILE._04402_ ;
 wire \u_cpu.REG_FILE._04403_ ;
 wire \u_cpu.REG_FILE._04404_ ;
 wire \u_cpu.REG_FILE._04405_ ;
 wire \u_cpu.REG_FILE._04406_ ;
 wire \u_cpu.REG_FILE._04407_ ;
 wire \u_cpu.REG_FILE._04408_ ;
 wire \u_cpu.REG_FILE._04409_ ;
 wire \u_cpu.REG_FILE._04410_ ;
 wire \u_cpu.REG_FILE._04411_ ;
 wire \u_cpu.REG_FILE._04412_ ;
 wire \u_cpu.REG_FILE._04413_ ;
 wire \u_cpu.REG_FILE._04414_ ;
 wire \u_cpu.REG_FILE._04415_ ;
 wire \u_cpu.REG_FILE._04416_ ;
 wire \u_cpu.REG_FILE._04417_ ;
 wire \u_cpu.REG_FILE._04418_ ;
 wire \u_cpu.REG_FILE._04419_ ;
 wire \u_cpu.REG_FILE._04420_ ;
 wire \u_cpu.REG_FILE._04421_ ;
 wire \u_cpu.REG_FILE._04422_ ;
 wire \u_cpu.REG_FILE._04423_ ;
 wire \u_cpu.REG_FILE._04424_ ;
 wire \u_cpu.REG_FILE._04425_ ;
 wire \u_cpu.REG_FILE._04426_ ;
 wire \u_cpu.REG_FILE._04427_ ;
 wire \u_cpu.REG_FILE._04428_ ;
 wire \u_cpu.REG_FILE._04429_ ;
 wire \u_cpu.REG_FILE._04430_ ;
 wire \u_cpu.REG_FILE._04431_ ;
 wire \u_cpu.REG_FILE._04432_ ;
 wire \u_cpu.REG_FILE._04433_ ;
 wire \u_cpu.REG_FILE._04434_ ;
 wire \u_cpu.REG_FILE._04435_ ;
 wire \u_cpu.REG_FILE._04436_ ;
 wire \u_cpu.REG_FILE._04437_ ;
 wire \u_cpu.REG_FILE._04438_ ;
 wire \u_cpu.REG_FILE._04439_ ;
 wire \u_cpu.REG_FILE._04440_ ;
 wire \u_cpu.REG_FILE._04441_ ;
 wire \u_cpu.REG_FILE._04442_ ;
 wire \u_cpu.REG_FILE._04443_ ;
 wire \u_cpu.REG_FILE._04444_ ;
 wire \u_cpu.REG_FILE._04445_ ;
 wire \u_cpu.REG_FILE._04446_ ;
 wire \u_cpu.REG_FILE._04447_ ;
 wire \u_cpu.REG_FILE._04448_ ;
 wire \u_cpu.REG_FILE._04449_ ;
 wire \u_cpu.REG_FILE._04450_ ;
 wire \u_cpu.REG_FILE._04451_ ;
 wire \u_cpu.REG_FILE._04452_ ;
 wire \u_cpu.REG_FILE._04453_ ;
 wire \u_cpu.REG_FILE._04454_ ;
 wire \u_cpu.REG_FILE._04455_ ;
 wire \u_cpu.REG_FILE._04456_ ;
 wire \u_cpu.REG_FILE._04457_ ;
 wire \u_cpu.REG_FILE._04458_ ;
 wire \u_cpu.REG_FILE._04459_ ;
 wire \u_cpu.REG_FILE._04460_ ;
 wire \u_cpu.REG_FILE._04461_ ;
 wire \u_cpu.REG_FILE._04462_ ;
 wire \u_cpu.REG_FILE._04463_ ;
 wire \u_cpu.REG_FILE._04464_ ;
 wire \u_cpu.REG_FILE._04465_ ;
 wire \u_cpu.REG_FILE._04466_ ;
 wire \u_cpu.REG_FILE._04467_ ;
 wire \u_cpu.REG_FILE._04468_ ;
 wire \u_cpu.REG_FILE._04469_ ;
 wire \u_cpu.REG_FILE._04470_ ;
 wire \u_cpu.REG_FILE._04471_ ;
 wire \u_cpu.REG_FILE._04472_ ;
 wire \u_cpu.REG_FILE._04473_ ;
 wire \u_cpu.REG_FILE._04474_ ;
 wire \u_cpu.REG_FILE._04475_ ;
 wire \u_cpu.REG_FILE._04476_ ;
 wire \u_cpu.REG_FILE._04477_ ;
 wire \u_cpu.REG_FILE._04478_ ;
 wire \u_cpu.REG_FILE._04479_ ;
 wire \u_cpu.REG_FILE._04480_ ;
 wire \u_cpu.REG_FILE._04481_ ;
 wire \u_cpu.REG_FILE._04482_ ;
 wire \u_cpu.REG_FILE._04483_ ;
 wire \u_cpu.REG_FILE._04484_ ;
 wire \u_cpu.REG_FILE._04485_ ;
 wire \u_cpu.REG_FILE._04486_ ;
 wire \u_cpu.REG_FILE._04487_ ;
 wire \u_cpu.REG_FILE._04488_ ;
 wire \u_cpu.REG_FILE._04489_ ;
 wire \u_cpu.REG_FILE._04490_ ;
 wire \u_cpu.REG_FILE._04491_ ;
 wire \u_cpu.REG_FILE._04492_ ;
 wire \u_cpu.REG_FILE._04493_ ;
 wire \u_cpu.REG_FILE._04494_ ;
 wire \u_cpu.REG_FILE._04495_ ;
 wire \u_cpu.REG_FILE._04496_ ;
 wire \u_cpu.REG_FILE._04497_ ;
 wire \u_cpu.REG_FILE._04498_ ;
 wire \u_cpu.REG_FILE._04499_ ;
 wire \u_cpu.REG_FILE._04500_ ;
 wire \u_cpu.REG_FILE._04501_ ;
 wire \u_cpu.REG_FILE._04502_ ;
 wire \u_cpu.REG_FILE._04503_ ;
 wire \u_cpu.REG_FILE._04504_ ;
 wire \u_cpu.REG_FILE._04505_ ;
 wire \u_cpu.REG_FILE._04506_ ;
 wire \u_cpu.REG_FILE._04507_ ;
 wire \u_cpu.REG_FILE._04508_ ;
 wire \u_cpu.REG_FILE._04509_ ;
 wire \u_cpu.REG_FILE._04510_ ;
 wire \u_cpu.REG_FILE._04511_ ;
 wire \u_cpu.REG_FILE._04512_ ;
 wire \u_cpu.REG_FILE._04513_ ;
 wire \u_cpu.REG_FILE._04514_ ;
 wire \u_cpu.REG_FILE._04515_ ;
 wire \u_cpu.REG_FILE._04516_ ;
 wire \u_cpu.REG_FILE._04517_ ;
 wire \u_cpu.REG_FILE._04518_ ;
 wire \u_cpu.REG_FILE._04519_ ;
 wire \u_cpu.REG_FILE._04520_ ;
 wire \u_cpu.REG_FILE._04521_ ;
 wire \u_cpu.REG_FILE._04522_ ;
 wire \u_cpu.REG_FILE._04523_ ;
 wire \u_cpu.REG_FILE._04524_ ;
 wire \u_cpu.REG_FILE._04525_ ;
 wire \u_cpu.REG_FILE._04526_ ;
 wire \u_cpu.REG_FILE._04527_ ;
 wire \u_cpu.REG_FILE._04528_ ;
 wire \u_cpu.REG_FILE._04529_ ;
 wire \u_cpu.REG_FILE._04530_ ;
 wire \u_cpu.REG_FILE._04531_ ;
 wire \u_cpu.REG_FILE._04532_ ;
 wire \u_cpu.REG_FILE._04533_ ;
 wire \u_cpu.REG_FILE._04534_ ;
 wire \u_cpu.REG_FILE._04535_ ;
 wire \u_cpu.REG_FILE._04536_ ;
 wire \u_cpu.REG_FILE._04537_ ;
 wire \u_cpu.REG_FILE._04538_ ;
 wire \u_cpu.REG_FILE._04539_ ;
 wire \u_cpu.REG_FILE._04540_ ;
 wire \u_cpu.REG_FILE._04541_ ;
 wire \u_cpu.REG_FILE._04542_ ;
 wire \u_cpu.REG_FILE._04543_ ;
 wire \u_cpu.REG_FILE._04544_ ;
 wire \u_cpu.REG_FILE._04545_ ;
 wire \u_cpu.REG_FILE._04546_ ;
 wire \u_cpu.REG_FILE._04547_ ;
 wire \u_cpu.REG_FILE._04548_ ;
 wire \u_cpu.REG_FILE._04549_ ;
 wire \u_cpu.REG_FILE._04550_ ;
 wire \u_cpu.REG_FILE._04551_ ;
 wire \u_cpu.REG_FILE._04552_ ;
 wire \u_cpu.REG_FILE._04553_ ;
 wire \u_cpu.REG_FILE._04554_ ;
 wire \u_cpu.REG_FILE._04555_ ;
 wire \u_cpu.REG_FILE._04556_ ;
 wire \u_cpu.REG_FILE._04557_ ;
 wire \u_cpu.REG_FILE._04558_ ;
 wire \u_cpu.REG_FILE._04559_ ;
 wire \u_cpu.REG_FILE._04560_ ;
 wire \u_cpu.REG_FILE._04561_ ;
 wire \u_cpu.REG_FILE._04562_ ;
 wire \u_cpu.REG_FILE._04563_ ;
 wire \u_cpu.REG_FILE._04564_ ;
 wire \u_cpu.REG_FILE._04565_ ;
 wire \u_cpu.REG_FILE._04566_ ;
 wire \u_cpu.REG_FILE._04567_ ;
 wire \u_cpu.REG_FILE._04568_ ;
 wire \u_cpu.REG_FILE._04569_ ;
 wire \u_cpu.REG_FILE._04570_ ;
 wire \u_cpu.REG_FILE._04571_ ;
 wire \u_cpu.REG_FILE._04572_ ;
 wire \u_cpu.REG_FILE._04573_ ;
 wire \u_cpu.REG_FILE._04574_ ;
 wire \u_cpu.REG_FILE._04575_ ;
 wire \u_cpu.REG_FILE._04576_ ;
 wire \u_cpu.REG_FILE._04577_ ;
 wire \u_cpu.REG_FILE._04578_ ;
 wire \u_cpu.REG_FILE._04579_ ;
 wire \u_cpu.REG_FILE._04580_ ;
 wire \u_cpu.REG_FILE._04581_ ;
 wire \u_cpu.REG_FILE._04582_ ;
 wire \u_cpu.REG_FILE._04583_ ;
 wire \u_cpu.REG_FILE._04584_ ;
 wire \u_cpu.REG_FILE._04585_ ;
 wire \u_cpu.REG_FILE._04586_ ;
 wire \u_cpu.REG_FILE._04587_ ;
 wire \u_cpu.REG_FILE._04588_ ;
 wire \u_cpu.REG_FILE._04589_ ;
 wire \u_cpu.REG_FILE._04590_ ;
 wire \u_cpu.REG_FILE._04591_ ;
 wire \u_cpu.REG_FILE._04592_ ;
 wire \u_cpu.REG_FILE._04593_ ;
 wire \u_cpu.REG_FILE._04594_ ;
 wire \u_cpu.REG_FILE._04595_ ;
 wire \u_cpu.REG_FILE._04596_ ;
 wire \u_cpu.REG_FILE._04597_ ;
 wire \u_cpu.REG_FILE._04598_ ;
 wire \u_cpu.REG_FILE._04599_ ;
 wire \u_cpu.REG_FILE._04600_ ;
 wire \u_cpu.REG_FILE._04601_ ;
 wire \u_cpu.REG_FILE._04602_ ;
 wire \u_cpu.REG_FILE._04603_ ;
 wire \u_cpu.REG_FILE._04604_ ;
 wire \u_cpu.REG_FILE._04605_ ;
 wire \u_cpu.REG_FILE._04606_ ;
 wire \u_cpu.REG_FILE._04607_ ;
 wire \u_cpu.REG_FILE._04608_ ;
 wire \u_cpu.REG_FILE._04609_ ;
 wire \u_cpu.REG_FILE._04610_ ;
 wire \u_cpu.REG_FILE._04611_ ;
 wire \u_cpu.REG_FILE._04612_ ;
 wire \u_cpu.REG_FILE._04613_ ;
 wire \u_cpu.REG_FILE._04614_ ;
 wire \u_cpu.REG_FILE._04615_ ;
 wire \u_cpu.REG_FILE._04616_ ;
 wire \u_cpu.REG_FILE._04617_ ;
 wire \u_cpu.REG_FILE._04618_ ;
 wire \u_cpu.REG_FILE._04619_ ;
 wire \u_cpu.REG_FILE._04620_ ;
 wire \u_cpu.REG_FILE._04621_ ;
 wire \u_cpu.REG_FILE._04622_ ;
 wire \u_cpu.REG_FILE._04623_ ;
 wire \u_cpu.REG_FILE._04624_ ;
 wire \u_cpu.REG_FILE._04625_ ;
 wire \u_cpu.REG_FILE._04626_ ;
 wire \u_cpu.REG_FILE._04627_ ;
 wire \u_cpu.REG_FILE._04628_ ;
 wire \u_cpu.REG_FILE._04629_ ;
 wire \u_cpu.REG_FILE._04630_ ;
 wire \u_cpu.REG_FILE._04631_ ;
 wire \u_cpu.REG_FILE._04632_ ;
 wire \u_cpu.REG_FILE._04633_ ;
 wire \u_cpu.REG_FILE._04634_ ;
 wire \u_cpu.REG_FILE._04635_ ;
 wire \u_cpu.REG_FILE._04636_ ;
 wire \u_cpu.REG_FILE._04637_ ;
 wire \u_cpu.REG_FILE._04638_ ;
 wire \u_cpu.REG_FILE._04639_ ;
 wire \u_cpu.REG_FILE._04640_ ;
 wire \u_cpu.REG_FILE._04641_ ;
 wire \u_cpu.REG_FILE._04642_ ;
 wire \u_cpu.REG_FILE._04643_ ;
 wire \u_cpu.REG_FILE._04644_ ;
 wire \u_cpu.REG_FILE._04645_ ;
 wire \u_cpu.REG_FILE._04646_ ;
 wire \u_cpu.REG_FILE._04647_ ;
 wire \u_cpu.REG_FILE._04648_ ;
 wire \u_cpu.REG_FILE._04649_ ;
 wire \u_cpu.REG_FILE._04650_ ;
 wire \u_cpu.REG_FILE._04651_ ;
 wire \u_cpu.REG_FILE._04652_ ;
 wire \u_cpu.REG_FILE._04653_ ;
 wire \u_cpu.REG_FILE._04654_ ;
 wire \u_cpu.REG_FILE._04655_ ;
 wire \u_cpu.REG_FILE._04656_ ;
 wire \u_cpu.REG_FILE._04657_ ;
 wire \u_cpu.REG_FILE._04658_ ;
 wire \u_cpu.REG_FILE._04659_ ;
 wire \u_cpu.REG_FILE._04660_ ;
 wire \u_cpu.REG_FILE._04661_ ;
 wire \u_cpu.REG_FILE._04662_ ;
 wire \u_cpu.REG_FILE._04663_ ;
 wire \u_cpu.REG_FILE._04664_ ;
 wire \u_cpu.REG_FILE._04665_ ;
 wire \u_cpu.REG_FILE._04666_ ;
 wire \u_cpu.REG_FILE._04667_ ;
 wire \u_cpu.REG_FILE._04668_ ;
 wire \u_cpu.REG_FILE._04669_ ;
 wire \u_cpu.REG_FILE._04670_ ;
 wire \u_cpu.REG_FILE._04671_ ;
 wire \u_cpu.REG_FILE._04672_ ;
 wire \u_cpu.REG_FILE._04673_ ;
 wire \u_cpu.REG_FILE._04674_ ;
 wire \u_cpu.REG_FILE._04675_ ;
 wire \u_cpu.REG_FILE._04676_ ;
 wire \u_cpu.REG_FILE._04677_ ;
 wire \u_cpu.REG_FILE._04678_ ;
 wire \u_cpu.REG_FILE._04679_ ;
 wire \u_cpu.REG_FILE._04680_ ;
 wire \u_cpu.REG_FILE._04681_ ;
 wire \u_cpu.REG_FILE._04682_ ;
 wire \u_cpu.REG_FILE._04683_ ;
 wire \u_cpu.REG_FILE._04684_ ;
 wire \u_cpu.REG_FILE._04685_ ;
 wire \u_cpu.REG_FILE._04686_ ;
 wire \u_cpu.REG_FILE._04687_ ;
 wire \u_cpu.REG_FILE._04688_ ;
 wire \u_cpu.REG_FILE._04689_ ;
 wire \u_cpu.REG_FILE._04690_ ;
 wire \u_cpu.REG_FILE._04691_ ;
 wire \u_cpu.REG_FILE._04692_ ;
 wire \u_cpu.REG_FILE._04693_ ;
 wire \u_cpu.REG_FILE._04694_ ;
 wire \u_cpu.REG_FILE._04695_ ;
 wire \u_cpu.REG_FILE._04696_ ;
 wire \u_cpu.REG_FILE._04697_ ;
 wire \u_cpu.REG_FILE._04698_ ;
 wire \u_cpu.REG_FILE._04699_ ;
 wire \u_cpu.REG_FILE._04700_ ;
 wire \u_cpu.REG_FILE._04701_ ;
 wire \u_cpu.REG_FILE._04702_ ;
 wire \u_cpu.REG_FILE._04703_ ;
 wire \u_cpu.REG_FILE._04704_ ;
 wire \u_cpu.REG_FILE._04705_ ;
 wire \u_cpu.REG_FILE._04706_ ;
 wire \u_cpu.REG_FILE._04707_ ;
 wire \u_cpu.REG_FILE._04708_ ;
 wire \u_cpu.REG_FILE._04709_ ;
 wire \u_cpu.REG_FILE._04710_ ;
 wire \u_cpu.REG_FILE._04711_ ;
 wire \u_cpu.REG_FILE._04712_ ;
 wire \u_cpu.REG_FILE._04713_ ;
 wire \u_cpu.REG_FILE._04714_ ;
 wire \u_cpu.REG_FILE._04715_ ;
 wire \u_cpu.REG_FILE._04716_ ;
 wire \u_cpu.REG_FILE._04717_ ;
 wire \u_cpu.REG_FILE._04718_ ;
 wire \u_cpu.REG_FILE._04719_ ;
 wire \u_cpu.REG_FILE._04720_ ;
 wire \u_cpu.REG_FILE._04721_ ;
 wire \u_cpu.REG_FILE._04722_ ;
 wire \u_cpu.REG_FILE._04723_ ;
 wire \u_cpu.REG_FILE._04724_ ;
 wire \u_cpu.REG_FILE._04725_ ;
 wire \u_cpu.REG_FILE._04726_ ;
 wire \u_cpu.REG_FILE._04727_ ;
 wire \u_cpu.REG_FILE._04728_ ;
 wire \u_cpu.REG_FILE._04729_ ;
 wire \u_cpu.REG_FILE._04730_ ;
 wire \u_cpu.REG_FILE._04731_ ;
 wire \u_cpu.REG_FILE._04732_ ;
 wire \u_cpu.REG_FILE._04733_ ;
 wire \u_cpu.REG_FILE._04734_ ;
 wire \u_cpu.REG_FILE._04735_ ;
 wire \u_cpu.REG_FILE._04736_ ;
 wire \u_cpu.REG_FILE._04737_ ;
 wire \u_cpu.REG_FILE._04738_ ;
 wire \u_cpu.REG_FILE._04739_ ;
 wire \u_cpu.REG_FILE._04740_ ;
 wire \u_cpu.REG_FILE._04741_ ;
 wire \u_cpu.REG_FILE._04742_ ;
 wire \u_cpu.REG_FILE._04743_ ;
 wire \u_cpu.REG_FILE._04744_ ;
 wire \u_cpu.REG_FILE._04745_ ;
 wire \u_cpu.REG_FILE._04746_ ;
 wire \u_cpu.REG_FILE._04747_ ;
 wire \u_cpu.REG_FILE._04748_ ;
 wire \u_cpu.REG_FILE._04749_ ;
 wire \u_cpu.REG_FILE._04750_ ;
 wire \u_cpu.REG_FILE._04751_ ;
 wire \u_cpu.REG_FILE._04752_ ;
 wire \u_cpu.REG_FILE._04753_ ;
 wire \u_cpu.REG_FILE._04754_ ;
 wire \u_cpu.REG_FILE._04755_ ;
 wire \u_cpu.REG_FILE._04756_ ;
 wire \u_cpu.REG_FILE._04757_ ;
 wire \u_cpu.REG_FILE._04758_ ;
 wire \u_cpu.REG_FILE._04759_ ;
 wire \u_cpu.REG_FILE._04760_ ;
 wire \u_cpu.REG_FILE._04761_ ;
 wire \u_cpu.REG_FILE._04762_ ;
 wire \u_cpu.REG_FILE._04763_ ;
 wire \u_cpu.REG_FILE._04764_ ;
 wire \u_cpu.REG_FILE._04765_ ;
 wire \u_cpu.REG_FILE._04766_ ;
 wire \u_cpu.REG_FILE._04767_ ;
 wire \u_cpu.REG_FILE._04768_ ;
 wire \u_cpu.REG_FILE._04769_ ;
 wire \u_cpu.REG_FILE._04770_ ;
 wire \u_cpu.REG_FILE._04771_ ;
 wire \u_cpu.REG_FILE._04772_ ;
 wire \u_cpu.REG_FILE._04773_ ;
 wire \u_cpu.REG_FILE._04774_ ;
 wire \u_cpu.REG_FILE._04775_ ;
 wire \u_cpu.REG_FILE._04776_ ;
 wire \u_cpu.REG_FILE._04777_ ;
 wire \u_cpu.REG_FILE._04778_ ;
 wire \u_cpu.REG_FILE._04779_ ;
 wire \u_cpu.REG_FILE._04780_ ;
 wire \u_cpu.REG_FILE._04781_ ;
 wire \u_cpu.REG_FILE._04782_ ;
 wire \u_cpu.REG_FILE._04783_ ;
 wire \u_cpu.REG_FILE._04784_ ;
 wire \u_cpu.REG_FILE._04785_ ;
 wire \u_cpu.REG_FILE._04786_ ;
 wire \u_cpu.REG_FILE._04787_ ;
 wire \u_cpu.REG_FILE._04788_ ;
 wire \u_cpu.REG_FILE._04789_ ;
 wire \u_cpu.REG_FILE._04790_ ;
 wire \u_cpu.REG_FILE._04791_ ;
 wire \u_cpu.REG_FILE._04792_ ;
 wire \u_cpu.REG_FILE._04793_ ;
 wire \u_cpu.REG_FILE._04794_ ;
 wire \u_cpu.REG_FILE._04795_ ;
 wire \u_cpu.REG_FILE._04796_ ;
 wire \u_cpu.REG_FILE._04797_ ;
 wire \u_cpu.REG_FILE._04798_ ;
 wire \u_cpu.REG_FILE._04799_ ;
 wire \u_cpu.REG_FILE._04800_ ;
 wire \u_cpu.REG_FILE._04801_ ;
 wire \u_cpu.REG_FILE._04802_ ;
 wire \u_cpu.REG_FILE._04803_ ;
 wire \u_cpu.REG_FILE._04804_ ;
 wire \u_cpu.REG_FILE._04805_ ;
 wire \u_cpu.REG_FILE._04806_ ;
 wire \u_cpu.REG_FILE._04807_ ;
 wire \u_cpu.REG_FILE._04808_ ;
 wire \u_cpu.REG_FILE._04809_ ;
 wire \u_cpu.REG_FILE._04810_ ;
 wire \u_cpu.REG_FILE._04811_ ;
 wire \u_cpu.REG_FILE._04812_ ;
 wire \u_cpu.REG_FILE._04813_ ;
 wire \u_cpu.REG_FILE._04814_ ;
 wire \u_cpu.REG_FILE._04815_ ;
 wire \u_cpu.REG_FILE._04816_ ;
 wire \u_cpu.REG_FILE._04817_ ;
 wire \u_cpu.REG_FILE._04818_ ;
 wire \u_cpu.REG_FILE._04819_ ;
 wire \u_cpu.REG_FILE._04820_ ;
 wire \u_cpu.REG_FILE._04821_ ;
 wire \u_cpu.REG_FILE._04822_ ;
 wire \u_cpu.REG_FILE._04823_ ;
 wire \u_cpu.REG_FILE._04824_ ;
 wire \u_cpu.REG_FILE._04825_ ;
 wire \u_cpu.REG_FILE._04826_ ;
 wire \u_cpu.REG_FILE._04827_ ;
 wire \u_cpu.REG_FILE._04828_ ;
 wire \u_cpu.REG_FILE._04829_ ;
 wire \u_cpu.REG_FILE._04830_ ;
 wire \u_cpu.REG_FILE._04831_ ;
 wire \u_cpu.REG_FILE._04832_ ;
 wire \u_cpu.REG_FILE._04833_ ;
 wire \u_cpu.REG_FILE._04834_ ;
 wire \u_cpu.REG_FILE._04835_ ;
 wire \u_cpu.REG_FILE._04836_ ;
 wire \u_cpu.REG_FILE._04837_ ;
 wire \u_cpu.REG_FILE._04838_ ;
 wire \u_cpu.REG_FILE._04839_ ;
 wire \u_cpu.REG_FILE._04840_ ;
 wire \u_cpu.REG_FILE._04841_ ;
 wire \u_cpu.REG_FILE._04842_ ;
 wire \u_cpu.REG_FILE._04843_ ;
 wire \u_cpu.REG_FILE._04844_ ;
 wire \u_cpu.REG_FILE._04845_ ;
 wire \u_cpu.REG_FILE._04846_ ;
 wire \u_cpu.REG_FILE._04847_ ;
 wire \u_cpu.REG_FILE._04848_ ;
 wire \u_cpu.REG_FILE._04849_ ;
 wire \u_cpu.REG_FILE._04850_ ;
 wire \u_cpu.REG_FILE._04851_ ;
 wire \u_cpu.REG_FILE._04852_ ;
 wire \u_cpu.REG_FILE._04853_ ;
 wire \u_cpu.REG_FILE._04854_ ;
 wire \u_cpu.REG_FILE._04855_ ;
 wire \u_cpu.REG_FILE._04856_ ;
 wire \u_cpu.REG_FILE._04857_ ;
 wire \u_cpu.REG_FILE._04858_ ;
 wire \u_cpu.REG_FILE._04859_ ;
 wire \u_cpu.REG_FILE._04860_ ;
 wire \u_cpu.REG_FILE._04861_ ;
 wire \u_cpu.REG_FILE._04862_ ;
 wire \u_cpu.REG_FILE._04863_ ;
 wire \u_cpu.REG_FILE._04864_ ;
 wire \u_cpu.REG_FILE._04865_ ;
 wire \u_cpu.REG_FILE._04866_ ;
 wire \u_cpu.REG_FILE._04867_ ;
 wire \u_cpu.REG_FILE._04868_ ;
 wire \u_cpu.REG_FILE._04869_ ;
 wire \u_cpu.REG_FILE._04870_ ;
 wire \u_cpu.REG_FILE._04871_ ;
 wire \u_cpu.REG_FILE._04872_ ;
 wire \u_cpu.REG_FILE._04873_ ;
 wire \u_cpu.REG_FILE._04874_ ;
 wire \u_cpu.REG_FILE._04875_ ;
 wire \u_cpu.REG_FILE._04876_ ;
 wire \u_cpu.REG_FILE._04877_ ;
 wire \u_cpu.REG_FILE._04878_ ;
 wire \u_cpu.REG_FILE._04879_ ;
 wire \u_cpu.REG_FILE._04880_ ;
 wire \u_cpu.REG_FILE._04881_ ;
 wire \u_cpu.REG_FILE._04882_ ;
 wire \u_cpu.REG_FILE._04883_ ;
 wire \u_cpu.REG_FILE._04884_ ;
 wire \u_cpu.REG_FILE._04885_ ;
 wire \u_cpu.REG_FILE._04886_ ;
 wire \u_cpu.REG_FILE._04887_ ;
 wire \u_cpu.REG_FILE._04888_ ;
 wire \u_cpu.REG_FILE._04889_ ;
 wire \u_cpu.REG_FILE._04890_ ;
 wire \u_cpu.REG_FILE._04891_ ;
 wire \u_cpu.REG_FILE._04892_ ;
 wire \u_cpu.REG_FILE._04893_ ;
 wire \u_cpu.REG_FILE._04894_ ;
 wire \u_cpu.REG_FILE._04895_ ;
 wire \u_cpu.REG_FILE._04896_ ;
 wire \u_cpu.REG_FILE._04897_ ;
 wire \u_cpu.REG_FILE._04898_ ;
 wire \u_cpu.REG_FILE._04899_ ;
 wire \u_cpu.REG_FILE._04900_ ;
 wire \u_cpu.REG_FILE._04901_ ;
 wire \u_cpu.REG_FILE._04902_ ;
 wire \u_cpu.REG_FILE._04903_ ;
 wire \u_cpu.REG_FILE._04904_ ;
 wire \u_cpu.REG_FILE._04905_ ;
 wire \u_cpu.REG_FILE._04906_ ;
 wire \u_cpu.REG_FILE._04907_ ;
 wire \u_cpu.REG_FILE._04908_ ;
 wire \u_cpu.REG_FILE._04909_ ;
 wire \u_cpu.REG_FILE._04910_ ;
 wire \u_cpu.REG_FILE._04911_ ;
 wire \u_cpu.REG_FILE._04912_ ;
 wire \u_cpu.REG_FILE._04913_ ;
 wire \u_cpu.REG_FILE._04914_ ;
 wire \u_cpu.REG_FILE._04915_ ;
 wire \u_cpu.REG_FILE._04916_ ;
 wire \u_cpu.REG_FILE._04917_ ;
 wire \u_cpu.REG_FILE._04918_ ;
 wire \u_cpu.REG_FILE._04919_ ;
 wire \u_cpu.REG_FILE._04920_ ;
 wire \u_cpu.REG_FILE._04921_ ;
 wire \u_cpu.REG_FILE._04922_ ;
 wire \u_cpu.REG_FILE._04923_ ;
 wire \u_cpu.REG_FILE._04924_ ;
 wire \u_cpu.REG_FILE._04925_ ;
 wire \u_cpu.REG_FILE._04926_ ;
 wire \u_cpu.REG_FILE._04927_ ;
 wire \u_cpu.REG_FILE._04928_ ;
 wire \u_cpu.REG_FILE._04929_ ;
 wire \u_cpu.REG_FILE._04930_ ;
 wire \u_cpu.REG_FILE._04931_ ;
 wire \u_cpu.REG_FILE._04932_ ;
 wire \u_cpu.REG_FILE._04933_ ;
 wire \u_cpu.REG_FILE._04934_ ;
 wire \u_cpu.REG_FILE._04935_ ;
 wire \u_cpu.REG_FILE._04936_ ;
 wire \u_cpu.REG_FILE._04937_ ;
 wire \u_cpu.REG_FILE._04938_ ;
 wire \u_cpu.REG_FILE._04939_ ;
 wire \u_cpu.REG_FILE._04940_ ;
 wire \u_cpu.REG_FILE._04941_ ;
 wire \u_cpu.REG_FILE._04942_ ;
 wire \u_cpu.REG_FILE._04943_ ;
 wire \u_cpu.REG_FILE._04944_ ;
 wire \u_cpu.REG_FILE._04945_ ;
 wire \u_cpu.REG_FILE._04946_ ;
 wire \u_cpu.REG_FILE._04947_ ;
 wire \u_cpu.REG_FILE._04948_ ;
 wire \u_cpu.REG_FILE._04949_ ;
 wire \u_cpu.REG_FILE._04950_ ;
 wire \u_cpu.REG_FILE._04951_ ;
 wire \u_cpu.REG_FILE._04952_ ;
 wire \u_cpu.REG_FILE._04953_ ;
 wire \u_cpu.REG_FILE._04954_ ;
 wire \u_cpu.REG_FILE._04955_ ;
 wire \u_cpu.REG_FILE._04956_ ;
 wire \u_cpu.REG_FILE._04957_ ;
 wire \u_cpu.REG_FILE._04958_ ;
 wire \u_cpu.REG_FILE._04959_ ;
 wire \u_cpu.REG_FILE._04960_ ;
 wire \u_cpu.REG_FILE._04961_ ;
 wire \u_cpu.REG_FILE._04962_ ;
 wire \u_cpu.REG_FILE._04963_ ;
 wire \u_cpu.REG_FILE._04964_ ;
 wire \u_cpu.REG_FILE._04965_ ;
 wire \u_cpu.REG_FILE._04966_ ;
 wire \u_cpu.REG_FILE._04967_ ;
 wire \u_cpu.REG_FILE._04968_ ;
 wire \u_cpu.REG_FILE._04969_ ;
 wire \u_cpu.REG_FILE._04970_ ;
 wire \u_cpu.REG_FILE._04971_ ;
 wire \u_cpu.REG_FILE._04972_ ;
 wire \u_cpu.REG_FILE._04973_ ;
 wire \u_cpu.REG_FILE._04974_ ;
 wire \u_cpu.REG_FILE._04975_ ;
 wire \u_cpu.REG_FILE._04976_ ;
 wire \u_cpu.REG_FILE._04977_ ;
 wire \u_cpu.REG_FILE._04978_ ;
 wire \u_cpu.REG_FILE._04979_ ;
 wire \u_cpu.REG_FILE._04980_ ;
 wire \u_cpu.REG_FILE._04981_ ;
 wire \u_cpu.REG_FILE._04982_ ;
 wire \u_cpu.REG_FILE._04983_ ;
 wire \u_cpu.REG_FILE._04984_ ;
 wire \u_cpu.REG_FILE._04985_ ;
 wire \u_cpu.REG_FILE._04986_ ;
 wire \u_cpu.REG_FILE._04987_ ;
 wire \u_cpu.REG_FILE._04988_ ;
 wire \u_cpu.REG_FILE._04989_ ;
 wire \u_cpu.REG_FILE._04990_ ;
 wire \u_cpu.REG_FILE._04991_ ;
 wire \u_cpu.REG_FILE._04992_ ;
 wire \u_cpu.REG_FILE._04993_ ;
 wire \u_cpu.REG_FILE._04994_ ;
 wire \u_cpu.REG_FILE._04995_ ;
 wire \u_cpu.REG_FILE._04996_ ;
 wire \u_cpu.REG_FILE._04997_ ;
 wire \u_cpu.REG_FILE._04998_ ;
 wire \u_cpu.REG_FILE._04999_ ;
 wire \u_cpu.REG_FILE._05000_ ;
 wire \u_cpu.REG_FILE._05001_ ;
 wire \u_cpu.REG_FILE._05002_ ;
 wire \u_cpu.REG_FILE._05003_ ;
 wire \u_cpu.REG_FILE._05004_ ;
 wire \u_cpu.REG_FILE._05005_ ;
 wire \u_cpu.REG_FILE._05006_ ;
 wire \u_cpu.REG_FILE._05007_ ;
 wire \u_cpu.REG_FILE._05008_ ;
 wire \u_cpu.REG_FILE._05009_ ;
 wire \u_cpu.REG_FILE._05010_ ;
 wire \u_cpu.REG_FILE._05011_ ;
 wire \u_cpu.REG_FILE._05012_ ;
 wire \u_cpu.REG_FILE._05013_ ;
 wire \u_cpu.REG_FILE._05014_ ;
 wire \u_cpu.REG_FILE._05015_ ;
 wire \u_cpu.REG_FILE._05016_ ;
 wire \u_cpu.REG_FILE._05017_ ;
 wire \u_cpu.REG_FILE._05018_ ;
 wire \u_cpu.REG_FILE._05019_ ;
 wire \u_cpu.REG_FILE._05020_ ;
 wire \u_cpu.REG_FILE._05021_ ;
 wire \u_cpu.REG_FILE._05022_ ;
 wire \u_cpu.REG_FILE._05023_ ;
 wire \u_cpu.REG_FILE._05024_ ;
 wire \u_cpu.REG_FILE._05025_ ;
 wire \u_cpu.REG_FILE._05026_ ;
 wire \u_cpu.REG_FILE._05027_ ;
 wire \u_cpu.REG_FILE._05028_ ;
 wire \u_cpu.REG_FILE._05029_ ;
 wire \u_cpu.REG_FILE._05030_ ;
 wire \u_cpu.REG_FILE._05031_ ;
 wire \u_cpu.REG_FILE._05032_ ;
 wire \u_cpu.REG_FILE._05033_ ;
 wire \u_cpu.REG_FILE._05034_ ;
 wire \u_cpu.REG_FILE._05035_ ;
 wire \u_cpu.REG_FILE._05036_ ;
 wire \u_cpu.REG_FILE._05037_ ;
 wire \u_cpu.REG_FILE._05038_ ;
 wire \u_cpu.REG_FILE._05039_ ;
 wire \u_cpu.REG_FILE._05040_ ;
 wire \u_cpu.REG_FILE._05041_ ;
 wire \u_cpu.REG_FILE._05042_ ;
 wire \u_cpu.REG_FILE._05043_ ;
 wire \u_cpu.REG_FILE._05044_ ;
 wire \u_cpu.REG_FILE._05045_ ;
 wire \u_cpu.REG_FILE._05046_ ;
 wire \u_cpu.REG_FILE._05047_ ;
 wire \u_cpu.REG_FILE._05048_ ;
 wire \u_cpu.REG_FILE._05049_ ;
 wire \u_cpu.REG_FILE._05050_ ;
 wire \u_cpu.REG_FILE._05051_ ;
 wire \u_cpu.REG_FILE._05052_ ;
 wire \u_cpu.REG_FILE._05053_ ;
 wire \u_cpu.REG_FILE._05054_ ;
 wire \u_cpu.REG_FILE._05055_ ;
 wire \u_cpu.REG_FILE._05056_ ;
 wire \u_cpu.REG_FILE._05057_ ;
 wire \u_cpu.REG_FILE._05058_ ;
 wire \u_cpu.REG_FILE._05059_ ;
 wire \u_cpu.REG_FILE._05060_ ;
 wire \u_cpu.REG_FILE._05061_ ;
 wire \u_cpu.REG_FILE._05062_ ;
 wire \u_cpu.REG_FILE._05063_ ;
 wire \u_cpu.REG_FILE._05064_ ;
 wire \u_cpu.REG_FILE._05065_ ;
 wire \u_cpu.REG_FILE._05066_ ;
 wire \u_cpu.REG_FILE._05067_ ;
 wire \u_cpu.REG_FILE._05068_ ;
 wire \u_cpu.REG_FILE._05069_ ;
 wire \u_cpu.REG_FILE._05070_ ;
 wire \u_cpu.REG_FILE._05071_ ;
 wire \u_cpu.REG_FILE._05072_ ;
 wire \u_cpu.REG_FILE._05073_ ;
 wire \u_cpu.REG_FILE._05074_ ;
 wire \u_cpu.REG_FILE._05075_ ;
 wire \u_cpu.REG_FILE._05076_ ;
 wire \u_cpu.REG_FILE._05077_ ;
 wire \u_cpu.REG_FILE._05078_ ;
 wire \u_cpu.REG_FILE._05079_ ;
 wire \u_cpu.REG_FILE._05080_ ;
 wire \u_cpu.REG_FILE._05081_ ;
 wire \u_cpu.REG_FILE._05082_ ;
 wire \u_cpu.REG_FILE._05083_ ;
 wire \u_cpu.REG_FILE._05084_ ;
 wire \u_cpu.REG_FILE._05085_ ;
 wire \u_cpu.REG_FILE._05086_ ;
 wire \u_cpu.REG_FILE._05087_ ;
 wire \u_cpu.REG_FILE._05088_ ;
 wire \u_cpu.REG_FILE._05089_ ;
 wire \u_cpu.REG_FILE._05090_ ;
 wire \u_cpu.REG_FILE._05091_ ;
 wire \u_cpu.REG_FILE._05092_ ;
 wire \u_cpu.REG_FILE._05093_ ;
 wire \u_cpu.REG_FILE._05094_ ;
 wire \u_cpu.REG_FILE._05095_ ;
 wire \u_cpu.REG_FILE._05096_ ;
 wire \u_cpu.REG_FILE._05097_ ;
 wire \u_cpu.REG_FILE._05098_ ;
 wire \u_cpu.REG_FILE._05099_ ;
 wire \u_cpu.REG_FILE._05100_ ;
 wire \u_cpu.REG_FILE._05101_ ;
 wire \u_cpu.REG_FILE._05102_ ;
 wire \u_cpu.REG_FILE._05103_ ;
 wire \u_cpu.REG_FILE._05104_ ;
 wire \u_cpu.REG_FILE._05105_ ;
 wire \u_cpu.REG_FILE._05106_ ;
 wire \u_cpu.REG_FILE._05107_ ;
 wire \u_cpu.REG_FILE._05108_ ;
 wire \u_cpu.REG_FILE._05109_ ;
 wire \u_cpu.REG_FILE._05110_ ;
 wire \u_cpu.REG_FILE._05111_ ;
 wire \u_cpu.REG_FILE._05112_ ;
 wire \u_cpu.REG_FILE._05113_ ;
 wire \u_cpu.REG_FILE._05114_ ;
 wire \u_cpu.REG_FILE._05115_ ;
 wire \u_cpu.REG_FILE._05116_ ;
 wire \u_cpu.REG_FILE._05117_ ;
 wire \u_cpu.REG_FILE._05118_ ;
 wire \u_cpu.REG_FILE._05119_ ;
 wire \u_cpu.REG_FILE._05120_ ;
 wire \u_cpu.REG_FILE._05121_ ;
 wire \u_cpu.REG_FILE._05122_ ;
 wire \u_cpu.REG_FILE._05123_ ;
 wire \u_cpu.REG_FILE._05124_ ;
 wire \u_cpu.REG_FILE._05125_ ;
 wire \u_cpu.REG_FILE._05126_ ;
 wire \u_cpu.REG_FILE._05127_ ;
 wire \u_cpu.REG_FILE._05128_ ;
 wire \u_cpu.REG_FILE._05129_ ;
 wire \u_cpu.REG_FILE._05130_ ;
 wire \u_cpu.REG_FILE._05131_ ;
 wire \u_cpu.REG_FILE._05132_ ;
 wire \u_cpu.REG_FILE._05133_ ;
 wire \u_cpu.REG_FILE._05134_ ;
 wire \u_cpu.REG_FILE._05135_ ;
 wire \u_cpu.REG_FILE._05136_ ;
 wire \u_cpu.REG_FILE._05137_ ;
 wire \u_cpu.REG_FILE._05138_ ;
 wire \u_cpu.REG_FILE._05139_ ;
 wire \u_cpu.REG_FILE._05140_ ;
 wire \u_cpu.REG_FILE._05141_ ;
 wire \u_cpu.REG_FILE._05142_ ;
 wire \u_cpu.REG_FILE._05143_ ;
 wire \u_cpu.REG_FILE._05144_ ;
 wire \u_cpu.REG_FILE._05145_ ;
 wire \u_cpu.REG_FILE._05146_ ;
 wire \u_cpu.REG_FILE._05147_ ;
 wire \u_cpu.REG_FILE._05148_ ;
 wire \u_cpu.REG_FILE._05149_ ;
 wire \u_cpu.REG_FILE._05150_ ;
 wire \u_cpu.REG_FILE._05151_ ;
 wire \u_cpu.REG_FILE._05152_ ;
 wire \u_cpu.REG_FILE._05153_ ;
 wire \u_cpu.REG_FILE._05154_ ;
 wire \u_cpu.REG_FILE._05155_ ;
 wire \u_cpu.REG_FILE._05156_ ;
 wire \u_cpu.REG_FILE._05157_ ;
 wire \u_cpu.REG_FILE._05158_ ;
 wire \u_cpu.REG_FILE._05159_ ;
 wire \u_cpu.REG_FILE._05160_ ;
 wire \u_cpu.REG_FILE._05161_ ;
 wire \u_cpu.REG_FILE._05162_ ;
 wire \u_cpu.REG_FILE._05163_ ;
 wire \u_cpu.REG_FILE._05164_ ;
 wire \u_cpu.REG_FILE._05165_ ;
 wire \u_cpu.REG_FILE._05166_ ;
 wire \u_cpu.REG_FILE._05167_ ;
 wire \u_cpu.REG_FILE._05168_ ;
 wire \u_cpu.REG_FILE._05169_ ;
 wire \u_cpu.REG_FILE._05170_ ;
 wire \u_cpu.REG_FILE._05171_ ;
 wire \u_cpu.REG_FILE._05172_ ;
 wire \u_cpu.REG_FILE._05173_ ;
 wire \u_cpu.REG_FILE._05174_ ;
 wire \u_cpu.REG_FILE._05175_ ;
 wire \u_cpu.REG_FILE._05176_ ;
 wire \u_cpu.REG_FILE._05177_ ;
 wire \u_cpu.REG_FILE._05178_ ;
 wire \u_cpu.REG_FILE._05179_ ;
 wire \u_cpu.REG_FILE._05180_ ;
 wire \u_cpu.REG_FILE._05181_ ;
 wire \u_cpu.REG_FILE._05182_ ;
 wire \u_cpu.REG_FILE._05183_ ;
 wire \u_cpu.REG_FILE._05184_ ;
 wire \u_cpu.REG_FILE._05185_ ;
 wire \u_cpu.REG_FILE._05186_ ;
 wire \u_cpu.REG_FILE._05187_ ;
 wire \u_cpu.REG_FILE._05188_ ;
 wire \u_cpu.REG_FILE._05189_ ;
 wire \u_cpu.REG_FILE._05190_ ;
 wire \u_cpu.REG_FILE._05191_ ;
 wire \u_cpu.REG_FILE._05192_ ;
 wire \u_cpu.REG_FILE._05193_ ;
 wire \u_cpu.REG_FILE._05194_ ;
 wire \u_cpu.REG_FILE._05195_ ;
 wire \u_cpu.REG_FILE._05196_ ;
 wire \u_cpu.REG_FILE._05197_ ;
 wire \u_cpu.REG_FILE._05198_ ;
 wire \u_cpu.REG_FILE._05199_ ;
 wire \u_cpu.REG_FILE._05200_ ;
 wire \u_cpu.REG_FILE._05201_ ;
 wire \u_cpu.REG_FILE._05202_ ;
 wire \u_cpu.REG_FILE._05203_ ;
 wire \u_cpu.REG_FILE._05204_ ;
 wire \u_cpu.REG_FILE._05205_ ;
 wire \u_cpu.REG_FILE._05206_ ;
 wire \u_cpu.REG_FILE._05207_ ;
 wire \u_cpu.REG_FILE._05208_ ;
 wire \u_cpu.REG_FILE._05209_ ;
 wire \u_cpu.REG_FILE._05210_ ;
 wire \u_cpu.REG_FILE._05211_ ;
 wire \u_cpu.REG_FILE._05212_ ;
 wire \u_cpu.REG_FILE._05213_ ;
 wire \u_cpu.REG_FILE._05214_ ;
 wire \u_cpu.REG_FILE._05215_ ;
 wire \u_cpu.REG_FILE._05216_ ;
 wire \u_cpu.REG_FILE._05217_ ;
 wire \u_cpu.REG_FILE._05218_ ;
 wire \u_cpu.REG_FILE._05219_ ;
 wire \u_cpu.REG_FILE._05220_ ;
 wire \u_cpu.REG_FILE._05221_ ;
 wire \u_cpu.REG_FILE._05222_ ;
 wire \u_cpu.REG_FILE._05223_ ;
 wire \u_cpu.REG_FILE._05224_ ;
 wire \u_cpu.REG_FILE._05225_ ;
 wire \u_cpu.REG_FILE._05226_ ;
 wire \u_cpu.REG_FILE._05227_ ;
 wire \u_cpu.REG_FILE._05228_ ;
 wire \u_cpu.REG_FILE._05229_ ;
 wire \u_cpu.REG_FILE._05230_ ;
 wire \u_cpu.REG_FILE._05231_ ;
 wire \u_cpu.REG_FILE._05232_ ;
 wire \u_cpu.REG_FILE._05233_ ;
 wire \u_cpu.REG_FILE._05234_ ;
 wire \u_cpu.REG_FILE._05235_ ;
 wire \u_cpu.REG_FILE._05236_ ;
 wire \u_cpu.REG_FILE._05237_ ;
 wire \u_cpu.REG_FILE._05238_ ;
 wire \u_cpu.REG_FILE._05239_ ;
 wire \u_cpu.REG_FILE._05240_ ;
 wire \u_cpu.REG_FILE._05241_ ;
 wire \u_cpu.REG_FILE._05242_ ;
 wire \u_cpu.REG_FILE._05243_ ;
 wire \u_cpu.REG_FILE._05244_ ;
 wire \u_cpu.REG_FILE._05245_ ;
 wire \u_cpu.REG_FILE._05246_ ;
 wire \u_cpu.REG_FILE._05247_ ;
 wire \u_cpu.REG_FILE._05248_ ;
 wire \u_cpu.REG_FILE._05249_ ;
 wire \u_cpu.REG_FILE._05250_ ;
 wire \u_cpu.REG_FILE._05251_ ;
 wire \u_cpu.REG_FILE._05252_ ;
 wire \u_cpu.REG_FILE._05253_ ;
 wire \u_cpu.REG_FILE._05254_ ;
 wire \u_cpu.REG_FILE._05255_ ;
 wire \u_cpu.REG_FILE._05256_ ;
 wire \u_cpu.REG_FILE._05257_ ;
 wire \u_cpu.REG_FILE._05258_ ;
 wire \u_cpu.REG_FILE._05259_ ;
 wire \u_cpu.REG_FILE._05260_ ;
 wire \u_cpu.REG_FILE._05261_ ;
 wire \u_cpu.REG_FILE._05262_ ;
 wire \u_cpu.REG_FILE._05263_ ;
 wire \u_cpu.REG_FILE._05264_ ;
 wire \u_cpu.REG_FILE._05265_ ;
 wire \u_cpu.REG_FILE._05266_ ;
 wire \u_cpu.REG_FILE._05267_ ;
 wire \u_cpu.REG_FILE._05268_ ;
 wire \u_cpu.REG_FILE._05269_ ;
 wire \u_cpu.REG_FILE._05270_ ;
 wire \u_cpu.REG_FILE._05271_ ;
 wire \u_cpu.REG_FILE._05272_ ;
 wire \u_cpu.REG_FILE._05273_ ;
 wire \u_cpu.REG_FILE._05274_ ;
 wire \u_cpu.REG_FILE._05275_ ;
 wire \u_cpu.REG_FILE._05276_ ;
 wire \u_cpu.REG_FILE._05277_ ;
 wire \u_cpu.REG_FILE._05278_ ;
 wire \u_cpu.REG_FILE._05279_ ;
 wire \u_cpu.REG_FILE._05280_ ;
 wire \u_cpu.REG_FILE._05281_ ;
 wire \u_cpu.REG_FILE._05282_ ;
 wire \u_cpu.REG_FILE._05283_ ;
 wire \u_cpu.REG_FILE._05284_ ;
 wire \u_cpu.REG_FILE._05285_ ;
 wire \u_cpu.REG_FILE._05286_ ;
 wire \u_cpu.REG_FILE._05287_ ;
 wire \u_cpu.REG_FILE._05288_ ;
 wire \u_cpu.REG_FILE._05289_ ;
 wire \u_cpu.REG_FILE._05290_ ;
 wire \u_cpu.REG_FILE._05291_ ;
 wire \u_cpu.REG_FILE._05292_ ;
 wire \u_cpu.REG_FILE._05293_ ;
 wire \u_cpu.REG_FILE._05294_ ;
 wire \u_cpu.REG_FILE._05295_ ;
 wire \u_cpu.REG_FILE._05296_ ;
 wire \u_cpu.REG_FILE._05297_ ;
 wire \u_cpu.REG_FILE._05298_ ;
 wire \u_cpu.REG_FILE._05299_ ;
 wire \u_cpu.REG_FILE._05300_ ;
 wire \u_cpu.REG_FILE._05301_ ;
 wire \u_cpu.REG_FILE._05302_ ;
 wire \u_cpu.REG_FILE._05303_ ;
 wire \u_cpu.REG_FILE._05304_ ;
 wire \u_cpu.REG_FILE._05305_ ;
 wire \u_cpu.REG_FILE._05306_ ;
 wire \u_cpu.REG_FILE._05307_ ;
 wire \u_cpu.REG_FILE._05308_ ;
 wire \u_cpu.REG_FILE._05309_ ;
 wire \u_cpu.REG_FILE._05310_ ;
 wire \u_cpu.REG_FILE._05311_ ;
 wire \u_cpu.REG_FILE._05312_ ;
 wire \u_cpu.REG_FILE._05313_ ;
 wire \u_cpu.REG_FILE._05314_ ;
 wire \u_cpu.REG_FILE._05315_ ;
 wire \u_cpu.REG_FILE._05316_ ;
 wire \u_cpu.REG_FILE._05317_ ;
 wire \u_cpu.REG_FILE._05318_ ;
 wire \u_cpu.REG_FILE._05319_ ;
 wire \u_cpu.REG_FILE._05320_ ;
 wire \u_cpu.REG_FILE._05321_ ;
 wire \u_cpu.REG_FILE._05322_ ;
 wire \u_cpu.REG_FILE._05323_ ;
 wire \u_cpu.REG_FILE._05324_ ;
 wire \u_cpu.REG_FILE._05325_ ;
 wire \u_cpu.REG_FILE._05326_ ;
 wire \u_cpu.REG_FILE._05327_ ;
 wire \u_cpu.REG_FILE._05328_ ;
 wire \u_cpu.REG_FILE._05329_ ;
 wire \u_cpu.REG_FILE._05330_ ;
 wire \u_cpu.REG_FILE._05331_ ;
 wire \u_cpu.REG_FILE._05332_ ;
 wire \u_cpu.REG_FILE._05333_ ;
 wire \u_cpu.REG_FILE._05334_ ;
 wire \u_cpu.REG_FILE._05335_ ;
 wire \u_cpu.REG_FILE._05336_ ;
 wire \u_cpu.REG_FILE._05337_ ;
 wire \u_cpu.REG_FILE._05338_ ;
 wire \u_cpu.REG_FILE._05339_ ;
 wire \u_cpu.REG_FILE._05340_ ;
 wire \u_cpu.REG_FILE._05341_ ;
 wire \u_cpu.REG_FILE._05342_ ;
 wire \u_cpu.REG_FILE._05343_ ;
 wire \u_cpu.REG_FILE._05344_ ;
 wire \u_cpu.REG_FILE._05345_ ;
 wire \u_cpu.REG_FILE._05346_ ;
 wire \u_cpu.REG_FILE._05347_ ;
 wire \u_cpu.REG_FILE._05348_ ;
 wire \u_cpu.REG_FILE._05349_ ;
 wire \u_cpu.REG_FILE._05350_ ;
 wire \u_cpu.REG_FILE._05351_ ;
 wire \u_cpu.REG_FILE._05352_ ;
 wire \u_cpu.REG_FILE._05353_ ;
 wire \u_cpu.REG_FILE._05354_ ;
 wire \u_cpu.REG_FILE._05355_ ;
 wire \u_cpu.REG_FILE._05356_ ;
 wire \u_cpu.REG_FILE._05357_ ;
 wire \u_cpu.REG_FILE._05358_ ;
 wire \u_cpu.REG_FILE._05359_ ;
 wire \u_cpu.REG_FILE._05360_ ;
 wire \u_cpu.REG_FILE._05361_ ;
 wire \u_cpu.REG_FILE._05362_ ;
 wire \u_cpu.REG_FILE._05363_ ;
 wire \u_cpu.REG_FILE._05364_ ;
 wire \u_cpu.REG_FILE._05365_ ;
 wire \u_cpu.REG_FILE._05366_ ;
 wire \u_cpu.REG_FILE._05367_ ;
 wire \u_cpu.REG_FILE._05368_ ;
 wire \u_cpu.REG_FILE._05369_ ;
 wire \u_cpu.REG_FILE._05370_ ;
 wire \u_cpu.REG_FILE._05371_ ;
 wire \u_cpu.REG_FILE._05372_ ;
 wire \u_cpu.REG_FILE._05373_ ;
 wire \u_cpu.REG_FILE._05374_ ;
 wire \u_cpu.REG_FILE._05375_ ;
 wire \u_cpu.REG_FILE._05376_ ;
 wire \u_cpu.REG_FILE._05377_ ;
 wire \u_cpu.REG_FILE._05378_ ;
 wire \u_cpu.REG_FILE._05379_ ;
 wire \u_cpu.REG_FILE._05380_ ;
 wire \u_cpu.REG_FILE._05381_ ;
 wire \u_cpu.REG_FILE._05382_ ;
 wire \u_cpu.REG_FILE._05383_ ;
 wire \u_cpu.REG_FILE._05384_ ;
 wire \u_cpu.REG_FILE._05385_ ;
 wire \u_cpu.REG_FILE._05386_ ;
 wire \u_cpu.REG_FILE._05387_ ;
 wire \u_cpu.REG_FILE._05388_ ;
 wire \u_cpu.REG_FILE._05389_ ;
 wire \u_cpu.REG_FILE._05390_ ;
 wire \u_cpu.REG_FILE._05391_ ;
 wire \u_cpu.REG_FILE._05392_ ;
 wire \u_cpu.REG_FILE._05393_ ;
 wire \u_cpu.REG_FILE._05394_ ;
 wire \u_cpu.REG_FILE._05395_ ;
 wire \u_cpu.REG_FILE._05396_ ;
 wire \u_cpu.REG_FILE._05397_ ;
 wire \u_cpu.REG_FILE._05398_ ;
 wire \u_cpu.REG_FILE._05399_ ;
 wire \u_cpu.REG_FILE._05400_ ;
 wire \u_cpu.REG_FILE._05401_ ;
 wire \u_cpu.REG_FILE._05402_ ;
 wire \u_cpu.REG_FILE._05403_ ;
 wire \u_cpu.REG_FILE._05404_ ;
 wire \u_cpu.REG_FILE._05405_ ;
 wire \u_cpu.REG_FILE._05406_ ;
 wire \u_cpu.REG_FILE._05407_ ;
 wire \u_cpu.REG_FILE._05408_ ;
 wire \u_cpu.REG_FILE._05409_ ;
 wire \u_cpu.REG_FILE._05410_ ;
 wire \u_cpu.REG_FILE._05411_ ;
 wire \u_cpu.REG_FILE._05412_ ;
 wire \u_cpu.REG_FILE._05413_ ;
 wire \u_cpu.REG_FILE._05414_ ;
 wire \u_cpu.REG_FILE._05415_ ;
 wire \u_cpu.REG_FILE._05416_ ;
 wire \u_cpu.REG_FILE._05417_ ;
 wire \u_cpu.REG_FILE._05418_ ;
 wire \u_cpu.REG_FILE._05419_ ;
 wire \u_cpu.REG_FILE._05420_ ;
 wire \u_cpu.REG_FILE._05421_ ;
 wire \u_cpu.REG_FILE._05422_ ;
 wire \u_cpu.REG_FILE._05423_ ;
 wire \u_cpu.REG_FILE._05424_ ;
 wire \u_cpu.REG_FILE._05425_ ;
 wire \u_cpu.REG_FILE._05426_ ;
 wire \u_cpu.REG_FILE._05427_ ;
 wire \u_cpu.REG_FILE._05428_ ;
 wire \u_cpu.REG_FILE._05429_ ;
 wire \u_cpu.REG_FILE._05430_ ;
 wire \u_cpu.REG_FILE._05431_ ;
 wire \u_cpu.REG_FILE._05432_ ;
 wire \u_cpu.REG_FILE._05433_ ;
 wire \u_cpu.REG_FILE._05434_ ;
 wire \u_cpu.REG_FILE._05435_ ;
 wire \u_cpu.REG_FILE._05436_ ;
 wire \u_cpu.REG_FILE._05437_ ;
 wire \u_cpu.REG_FILE._05438_ ;
 wire \u_cpu.REG_FILE._05439_ ;
 wire \u_cpu.REG_FILE._05440_ ;
 wire \u_cpu.REG_FILE._05441_ ;
 wire \u_cpu.REG_FILE._05442_ ;
 wire \u_cpu.REG_FILE._05443_ ;
 wire \u_cpu.REG_FILE._05444_ ;
 wire \u_cpu.REG_FILE._05445_ ;
 wire \u_cpu.REG_FILE._05446_ ;
 wire \u_cpu.REG_FILE._05447_ ;
 wire \u_cpu.REG_FILE._05448_ ;
 wire \u_cpu.REG_FILE._05449_ ;
 wire \u_cpu.REG_FILE._05450_ ;
 wire \u_cpu.REG_FILE._05451_ ;
 wire \u_cpu.REG_FILE._05452_ ;
 wire \u_cpu.REG_FILE._05453_ ;
 wire \u_cpu.REG_FILE._05454_ ;
 wire \u_cpu.REG_FILE._05455_ ;
 wire \u_cpu.REG_FILE._05456_ ;
 wire \u_cpu.REG_FILE._05457_ ;
 wire \u_cpu.REG_FILE._05458_ ;
 wire \u_cpu.REG_FILE._05459_ ;
 wire \u_cpu.REG_FILE._05460_ ;
 wire \u_cpu.REG_FILE._05461_ ;
 wire \u_cpu.REG_FILE._05462_ ;
 wire \u_cpu.REG_FILE._05463_ ;
 wire \u_cpu.REG_FILE._05464_ ;
 wire \u_cpu.REG_FILE._05465_ ;
 wire \u_cpu.REG_FILE._05466_ ;
 wire \u_cpu.REG_FILE._05467_ ;
 wire \u_cpu.REG_FILE._05468_ ;
 wire \u_cpu.REG_FILE._05469_ ;
 wire \u_cpu.REG_FILE._05470_ ;
 wire \u_cpu.REG_FILE._05471_ ;
 wire \u_cpu.REG_FILE._05472_ ;
 wire \u_cpu.REG_FILE._05473_ ;
 wire \u_cpu.REG_FILE._05474_ ;
 wire \u_cpu.REG_FILE._05475_ ;
 wire \u_cpu.REG_FILE._05476_ ;
 wire \u_cpu.REG_FILE._05477_ ;
 wire \u_cpu.REG_FILE._05478_ ;
 wire \u_cpu.REG_FILE._05479_ ;
 wire \u_cpu.REG_FILE._05480_ ;
 wire \u_cpu.REG_FILE._05481_ ;
 wire \u_cpu.REG_FILE._05482_ ;
 wire \u_cpu.REG_FILE._05483_ ;
 wire \u_cpu.REG_FILE._05484_ ;
 wire \u_cpu.REG_FILE._05485_ ;
 wire \u_cpu.REG_FILE._05486_ ;
 wire \u_cpu.REG_FILE._05487_ ;
 wire \u_cpu.REG_FILE._05488_ ;
 wire \u_cpu.REG_FILE._05489_ ;
 wire \u_cpu.REG_FILE._05490_ ;
 wire \u_cpu.REG_FILE._05491_ ;
 wire \u_cpu.REG_FILE._05492_ ;
 wire \u_cpu.REG_FILE._05493_ ;
 wire \u_cpu.REG_FILE._05494_ ;
 wire \u_cpu.REG_FILE._05495_ ;
 wire \u_cpu.REG_FILE._05496_ ;
 wire \u_cpu.REG_FILE._05497_ ;
 wire \u_cpu.REG_FILE._05498_ ;
 wire \u_cpu.REG_FILE._05499_ ;
 wire \u_cpu.REG_FILE._05500_ ;
 wire \u_cpu.REG_FILE._05501_ ;
 wire \u_cpu.REG_FILE._05502_ ;
 wire \u_cpu.REG_FILE._05503_ ;
 wire \u_cpu.REG_FILE._05504_ ;
 wire \u_cpu.REG_FILE._05505_ ;
 wire \u_cpu.REG_FILE._05506_ ;
 wire \u_cpu.REG_FILE._05507_ ;
 wire \u_cpu.REG_FILE._05508_ ;
 wire \u_cpu.REG_FILE._05509_ ;
 wire \u_cpu.REG_FILE._05510_ ;
 wire \u_cpu.REG_FILE._05511_ ;
 wire \u_cpu.REG_FILE._05512_ ;
 wire \u_cpu.REG_FILE._05513_ ;
 wire \u_cpu.REG_FILE._05514_ ;
 wire \u_cpu.REG_FILE._05515_ ;
 wire \u_cpu.REG_FILE._05516_ ;
 wire \u_cpu.REG_FILE._05517_ ;
 wire \u_cpu.REG_FILE._05518_ ;
 wire \u_cpu.REG_FILE._05519_ ;
 wire \u_cpu.REG_FILE._05520_ ;
 wire \u_cpu.REG_FILE._05521_ ;
 wire \u_cpu.REG_FILE._05522_ ;
 wire \u_cpu.REG_FILE._05523_ ;
 wire \u_cpu.REG_FILE._05524_ ;
 wire \u_cpu.REG_FILE._05525_ ;
 wire \u_cpu.REG_FILE._05526_ ;
 wire \u_cpu.REG_FILE._05527_ ;
 wire \u_cpu.REG_FILE._05528_ ;
 wire \u_cpu.REG_FILE._05529_ ;
 wire \u_cpu.REG_FILE._05530_ ;
 wire \u_cpu.REG_FILE._05531_ ;
 wire \u_cpu.REG_FILE._05532_ ;
 wire \u_cpu.REG_FILE._05533_ ;
 wire \u_cpu.REG_FILE._05534_ ;
 wire \u_cpu.REG_FILE._05535_ ;
 wire \u_cpu.REG_FILE._05536_ ;
 wire \u_cpu.REG_FILE._05537_ ;
 wire \u_cpu.REG_FILE._05538_ ;
 wire \u_cpu.REG_FILE._05539_ ;
 wire \u_cpu.REG_FILE._05540_ ;
 wire \u_cpu.REG_FILE._05541_ ;
 wire \u_cpu.REG_FILE._05542_ ;
 wire \u_cpu.REG_FILE._05543_ ;
 wire \u_cpu.REG_FILE._05544_ ;
 wire \u_cpu.REG_FILE._05545_ ;
 wire \u_cpu.REG_FILE._05546_ ;
 wire \u_cpu.REG_FILE._05547_ ;
 wire \u_cpu.REG_FILE._05548_ ;
 wire \u_cpu.REG_FILE._05549_ ;
 wire \u_cpu.REG_FILE._05550_ ;
 wire \u_cpu.REG_FILE._05551_ ;
 wire \u_cpu.REG_FILE._05552_ ;
 wire \u_cpu.REG_FILE._05553_ ;
 wire \u_cpu.REG_FILE._05554_ ;
 wire \u_cpu.REG_FILE._05555_ ;
 wire \u_cpu.REG_FILE._05556_ ;
 wire \u_cpu.REG_FILE._05557_ ;
 wire \u_cpu.REG_FILE._05558_ ;
 wire \u_cpu.REG_FILE._05559_ ;
 wire \u_cpu.REG_FILE._05560_ ;
 wire \u_cpu.REG_FILE._05561_ ;
 wire \u_cpu.REG_FILE._05562_ ;
 wire \u_cpu.REG_FILE._05563_ ;
 wire \u_cpu.REG_FILE._05564_ ;
 wire \u_cpu.REG_FILE._05565_ ;
 wire \u_cpu.REG_FILE._05566_ ;
 wire \u_cpu.REG_FILE._05567_ ;
 wire \u_cpu.REG_FILE._05568_ ;
 wire \u_cpu.REG_FILE._05569_ ;
 wire \u_cpu.REG_FILE._05570_ ;
 wire \u_cpu.REG_FILE._05571_ ;
 wire \u_cpu.REG_FILE._05572_ ;
 wire \u_cpu.REG_FILE._05573_ ;
 wire \u_cpu.REG_FILE._05574_ ;
 wire \u_cpu.REG_FILE._05575_ ;
 wire \u_cpu.REG_FILE._05576_ ;
 wire \u_cpu.REG_FILE._05577_ ;
 wire \u_cpu.REG_FILE._05578_ ;
 wire \u_cpu.REG_FILE._05579_ ;
 wire \u_cpu.REG_FILE._05580_ ;
 wire \u_cpu.REG_FILE._05581_ ;
 wire \u_cpu.REG_FILE._05582_ ;
 wire \u_cpu.REG_FILE._05583_ ;
 wire \u_cpu.REG_FILE._05584_ ;
 wire \u_cpu.REG_FILE._05585_ ;
 wire \u_cpu.REG_FILE._05586_ ;
 wire \u_cpu.REG_FILE._05587_ ;
 wire \u_cpu.REG_FILE._05588_ ;
 wire \u_cpu.REG_FILE._05589_ ;
 wire \u_cpu.REG_FILE._05590_ ;
 wire \u_cpu.REG_FILE._05591_ ;
 wire \u_cpu.REG_FILE._05592_ ;
 wire \u_cpu.REG_FILE._05593_ ;
 wire \u_cpu.REG_FILE._05594_ ;
 wire \u_cpu.REG_FILE._05595_ ;
 wire \u_cpu.REG_FILE._05596_ ;
 wire \u_cpu.REG_FILE._05597_ ;
 wire \u_cpu.REG_FILE._05598_ ;
 wire \u_cpu.REG_FILE._05599_ ;
 wire \u_cpu.REG_FILE._05600_ ;
 wire \u_cpu.REG_FILE._05601_ ;
 wire \u_cpu.REG_FILE._05602_ ;
 wire \u_cpu.REG_FILE._05603_ ;
 wire \u_cpu.REG_FILE._05604_ ;
 wire \u_cpu.REG_FILE._05605_ ;
 wire \u_cpu.REG_FILE._05606_ ;
 wire \u_cpu.REG_FILE._05607_ ;
 wire \u_cpu.REG_FILE._05608_ ;
 wire \u_cpu.REG_FILE._05609_ ;
 wire \u_cpu.REG_FILE._05610_ ;
 wire \u_cpu.REG_FILE._05611_ ;
 wire \u_cpu.REG_FILE._05612_ ;
 wire \u_cpu.REG_FILE._05613_ ;
 wire \u_cpu.REG_FILE._05614_ ;
 wire \u_cpu.REG_FILE._05615_ ;
 wire \u_cpu.REG_FILE._05616_ ;
 wire \u_cpu.REG_FILE._05617_ ;
 wire \u_cpu.REG_FILE._05618_ ;
 wire \u_cpu.REG_FILE._05619_ ;
 wire \u_cpu.REG_FILE._05620_ ;
 wire \u_cpu.REG_FILE._05621_ ;
 wire \u_cpu.REG_FILE._05622_ ;
 wire \u_cpu.REG_FILE._05623_ ;
 wire \u_cpu.REG_FILE._05624_ ;
 wire \u_cpu.REG_FILE._05625_ ;
 wire \u_cpu.REG_FILE._05626_ ;
 wire \u_cpu.REG_FILE._05627_ ;
 wire \u_cpu.REG_FILE._05628_ ;
 wire \u_cpu.REG_FILE._05629_ ;
 wire \u_cpu.REG_FILE._05630_ ;
 wire \u_cpu.REG_FILE._05631_ ;
 wire \u_cpu.REG_FILE._05632_ ;
 wire \u_cpu.REG_FILE._05633_ ;
 wire \u_cpu.REG_FILE._05634_ ;
 wire \u_cpu.REG_FILE._05635_ ;
 wire \u_cpu.REG_FILE._05636_ ;
 wire \u_cpu.REG_FILE._05637_ ;
 wire \u_cpu.REG_FILE._05638_ ;
 wire \u_cpu.REG_FILE._05639_ ;
 wire \u_cpu.REG_FILE._05640_ ;
 wire \u_cpu.REG_FILE._05641_ ;
 wire \u_cpu.REG_FILE._05642_ ;
 wire \u_cpu.REG_FILE._05643_ ;
 wire \u_cpu.REG_FILE._05644_ ;
 wire \u_cpu.REG_FILE._05645_ ;
 wire \u_cpu.REG_FILE._05646_ ;
 wire \u_cpu.REG_FILE._05647_ ;
 wire \u_cpu.REG_FILE._05648_ ;
 wire \u_cpu.REG_FILE._05649_ ;
 wire \u_cpu.REG_FILE._05650_ ;
 wire \u_cpu.REG_FILE._05651_ ;
 wire \u_cpu.REG_FILE._05652_ ;
 wire \u_cpu.REG_FILE._05653_ ;
 wire \u_cpu.REG_FILE._05654_ ;
 wire \u_cpu.REG_FILE._05655_ ;
 wire \u_cpu.REG_FILE._05656_ ;
 wire \u_cpu.REG_FILE._05657_ ;
 wire \u_cpu.REG_FILE._05658_ ;
 wire \u_cpu.REG_FILE._05659_ ;
 wire \u_cpu.REG_FILE._05660_ ;
 wire \u_cpu.REG_FILE._05661_ ;
 wire \u_cpu.REG_FILE._05662_ ;
 wire \u_cpu.REG_FILE._05663_ ;
 wire \u_cpu.REG_FILE._05664_ ;
 wire \u_cpu.REG_FILE._05665_ ;
 wire \u_cpu.REG_FILE._05666_ ;
 wire \u_cpu.REG_FILE._05667_ ;
 wire \u_cpu.REG_FILE._05668_ ;
 wire \u_cpu.REG_FILE._05669_ ;
 wire \u_cpu.REG_FILE._05670_ ;
 wire \u_cpu.REG_FILE._05671_ ;
 wire \u_cpu.REG_FILE._05672_ ;
 wire \u_cpu.REG_FILE._05673_ ;
 wire \u_cpu.REG_FILE._05674_ ;
 wire \u_cpu.REG_FILE._05675_ ;
 wire \u_cpu.REG_FILE._05676_ ;
 wire \u_cpu.REG_FILE._05677_ ;
 wire \u_cpu.REG_FILE._05678_ ;
 wire \u_cpu.REG_FILE._05679_ ;
 wire \u_cpu.REG_FILE._05680_ ;
 wire \u_cpu.REG_FILE._05681_ ;
 wire \u_cpu.REG_FILE._05682_ ;
 wire \u_cpu.REG_FILE._05683_ ;
 wire \u_cpu.REG_FILE._05684_ ;
 wire \u_cpu.REG_FILE._05685_ ;
 wire \u_cpu.REG_FILE._05686_ ;
 wire \u_cpu.REG_FILE._05687_ ;
 wire \u_cpu.REG_FILE._05688_ ;
 wire \u_cpu.REG_FILE._05689_ ;
 wire \u_cpu.REG_FILE.a3[0] ;
 wire \u_cpu.REG_FILE.a3[1] ;
 wire \u_cpu.REG_FILE.a3[2] ;
 wire \u_cpu.REG_FILE.a3[3] ;
 wire \u_cpu.REG_FILE.a3[4] ;
 wire \u_cpu.REG_FILE.rf[0][0] ;
 wire \u_cpu.REG_FILE.rf[0][10] ;
 wire \u_cpu.REG_FILE.rf[0][11] ;
 wire \u_cpu.REG_FILE.rf[0][12] ;
 wire \u_cpu.REG_FILE.rf[0][13] ;
 wire \u_cpu.REG_FILE.rf[0][14] ;
 wire \u_cpu.REG_FILE.rf[0][15] ;
 wire \u_cpu.REG_FILE.rf[0][16] ;
 wire \u_cpu.REG_FILE.rf[0][17] ;
 wire \u_cpu.REG_FILE.rf[0][18] ;
 wire \u_cpu.REG_FILE.rf[0][19] ;
 wire \u_cpu.REG_FILE.rf[0][1] ;
 wire \u_cpu.REG_FILE.rf[0][20] ;
 wire \u_cpu.REG_FILE.rf[0][21] ;
 wire \u_cpu.REG_FILE.rf[0][22] ;
 wire \u_cpu.REG_FILE.rf[0][23] ;
 wire \u_cpu.REG_FILE.rf[0][24] ;
 wire \u_cpu.REG_FILE.rf[0][25] ;
 wire \u_cpu.REG_FILE.rf[0][26] ;
 wire \u_cpu.REG_FILE.rf[0][27] ;
 wire \u_cpu.REG_FILE.rf[0][28] ;
 wire \u_cpu.REG_FILE.rf[0][29] ;
 wire \u_cpu.REG_FILE.rf[0][2] ;
 wire \u_cpu.REG_FILE.rf[0][30] ;
 wire \u_cpu.REG_FILE.rf[0][31] ;
 wire \u_cpu.REG_FILE.rf[0][3] ;
 wire \u_cpu.REG_FILE.rf[0][4] ;
 wire \u_cpu.REG_FILE.rf[0][5] ;
 wire \u_cpu.REG_FILE.rf[0][6] ;
 wire \u_cpu.REG_FILE.rf[0][7] ;
 wire \u_cpu.REG_FILE.rf[0][8] ;
 wire \u_cpu.REG_FILE.rf[0][9] ;
 wire \u_cpu.REG_FILE.rf[10][0] ;
 wire \u_cpu.REG_FILE.rf[10][10] ;
 wire \u_cpu.REG_FILE.rf[10][11] ;
 wire \u_cpu.REG_FILE.rf[10][12] ;
 wire \u_cpu.REG_FILE.rf[10][13] ;
 wire \u_cpu.REG_FILE.rf[10][14] ;
 wire \u_cpu.REG_FILE.rf[10][15] ;
 wire \u_cpu.REG_FILE.rf[10][16] ;
 wire \u_cpu.REG_FILE.rf[10][17] ;
 wire \u_cpu.REG_FILE.rf[10][18] ;
 wire \u_cpu.REG_FILE.rf[10][19] ;
 wire \u_cpu.REG_FILE.rf[10][1] ;
 wire \u_cpu.REG_FILE.rf[10][20] ;
 wire \u_cpu.REG_FILE.rf[10][21] ;
 wire \u_cpu.REG_FILE.rf[10][22] ;
 wire \u_cpu.REG_FILE.rf[10][23] ;
 wire \u_cpu.REG_FILE.rf[10][24] ;
 wire \u_cpu.REG_FILE.rf[10][25] ;
 wire \u_cpu.REG_FILE.rf[10][26] ;
 wire \u_cpu.REG_FILE.rf[10][27] ;
 wire \u_cpu.REG_FILE.rf[10][28] ;
 wire \u_cpu.REG_FILE.rf[10][29] ;
 wire \u_cpu.REG_FILE.rf[10][2] ;
 wire \u_cpu.REG_FILE.rf[10][30] ;
 wire \u_cpu.REG_FILE.rf[10][31] ;
 wire \u_cpu.REG_FILE.rf[10][3] ;
 wire \u_cpu.REG_FILE.rf[10][4] ;
 wire \u_cpu.REG_FILE.rf[10][5] ;
 wire \u_cpu.REG_FILE.rf[10][6] ;
 wire \u_cpu.REG_FILE.rf[10][7] ;
 wire \u_cpu.REG_FILE.rf[10][8] ;
 wire \u_cpu.REG_FILE.rf[10][9] ;
 wire \u_cpu.REG_FILE.rf[11][0] ;
 wire \u_cpu.REG_FILE.rf[11][10] ;
 wire \u_cpu.REG_FILE.rf[11][11] ;
 wire \u_cpu.REG_FILE.rf[11][12] ;
 wire \u_cpu.REG_FILE.rf[11][13] ;
 wire \u_cpu.REG_FILE.rf[11][14] ;
 wire \u_cpu.REG_FILE.rf[11][15] ;
 wire \u_cpu.REG_FILE.rf[11][16] ;
 wire \u_cpu.REG_FILE.rf[11][17] ;
 wire \u_cpu.REG_FILE.rf[11][18] ;
 wire \u_cpu.REG_FILE.rf[11][19] ;
 wire \u_cpu.REG_FILE.rf[11][1] ;
 wire \u_cpu.REG_FILE.rf[11][20] ;
 wire \u_cpu.REG_FILE.rf[11][21] ;
 wire \u_cpu.REG_FILE.rf[11][22] ;
 wire \u_cpu.REG_FILE.rf[11][23] ;
 wire \u_cpu.REG_FILE.rf[11][24] ;
 wire \u_cpu.REG_FILE.rf[11][25] ;
 wire \u_cpu.REG_FILE.rf[11][26] ;
 wire \u_cpu.REG_FILE.rf[11][27] ;
 wire \u_cpu.REG_FILE.rf[11][28] ;
 wire \u_cpu.REG_FILE.rf[11][29] ;
 wire \u_cpu.REG_FILE.rf[11][2] ;
 wire \u_cpu.REG_FILE.rf[11][30] ;
 wire \u_cpu.REG_FILE.rf[11][31] ;
 wire \u_cpu.REG_FILE.rf[11][3] ;
 wire \u_cpu.REG_FILE.rf[11][4] ;
 wire \u_cpu.REG_FILE.rf[11][5] ;
 wire \u_cpu.REG_FILE.rf[11][6] ;
 wire \u_cpu.REG_FILE.rf[11][7] ;
 wire \u_cpu.REG_FILE.rf[11][8] ;
 wire \u_cpu.REG_FILE.rf[11][9] ;
 wire \u_cpu.REG_FILE.rf[12][0] ;
 wire \u_cpu.REG_FILE.rf[12][10] ;
 wire \u_cpu.REG_FILE.rf[12][11] ;
 wire \u_cpu.REG_FILE.rf[12][12] ;
 wire \u_cpu.REG_FILE.rf[12][13] ;
 wire \u_cpu.REG_FILE.rf[12][14] ;
 wire \u_cpu.REG_FILE.rf[12][15] ;
 wire \u_cpu.REG_FILE.rf[12][16] ;
 wire \u_cpu.REG_FILE.rf[12][17] ;
 wire \u_cpu.REG_FILE.rf[12][18] ;
 wire \u_cpu.REG_FILE.rf[12][19] ;
 wire \u_cpu.REG_FILE.rf[12][1] ;
 wire \u_cpu.REG_FILE.rf[12][20] ;
 wire \u_cpu.REG_FILE.rf[12][21] ;
 wire \u_cpu.REG_FILE.rf[12][22] ;
 wire \u_cpu.REG_FILE.rf[12][23] ;
 wire \u_cpu.REG_FILE.rf[12][24] ;
 wire \u_cpu.REG_FILE.rf[12][25] ;
 wire \u_cpu.REG_FILE.rf[12][26] ;
 wire \u_cpu.REG_FILE.rf[12][27] ;
 wire \u_cpu.REG_FILE.rf[12][28] ;
 wire \u_cpu.REG_FILE.rf[12][29] ;
 wire \u_cpu.REG_FILE.rf[12][2] ;
 wire \u_cpu.REG_FILE.rf[12][30] ;
 wire \u_cpu.REG_FILE.rf[12][31] ;
 wire \u_cpu.REG_FILE.rf[12][3] ;
 wire \u_cpu.REG_FILE.rf[12][4] ;
 wire \u_cpu.REG_FILE.rf[12][5] ;
 wire \u_cpu.REG_FILE.rf[12][6] ;
 wire \u_cpu.REG_FILE.rf[12][7] ;
 wire \u_cpu.REG_FILE.rf[12][8] ;
 wire \u_cpu.REG_FILE.rf[12][9] ;
 wire \u_cpu.REG_FILE.rf[13][0] ;
 wire \u_cpu.REG_FILE.rf[13][10] ;
 wire \u_cpu.REG_FILE.rf[13][11] ;
 wire \u_cpu.REG_FILE.rf[13][12] ;
 wire \u_cpu.REG_FILE.rf[13][13] ;
 wire \u_cpu.REG_FILE.rf[13][14] ;
 wire \u_cpu.REG_FILE.rf[13][15] ;
 wire \u_cpu.REG_FILE.rf[13][16] ;
 wire \u_cpu.REG_FILE.rf[13][17] ;
 wire \u_cpu.REG_FILE.rf[13][18] ;
 wire \u_cpu.REG_FILE.rf[13][19] ;
 wire \u_cpu.REG_FILE.rf[13][1] ;
 wire \u_cpu.REG_FILE.rf[13][20] ;
 wire \u_cpu.REG_FILE.rf[13][21] ;
 wire \u_cpu.REG_FILE.rf[13][22] ;
 wire \u_cpu.REG_FILE.rf[13][23] ;
 wire \u_cpu.REG_FILE.rf[13][24] ;
 wire \u_cpu.REG_FILE.rf[13][25] ;
 wire \u_cpu.REG_FILE.rf[13][26] ;
 wire \u_cpu.REG_FILE.rf[13][27] ;
 wire \u_cpu.REG_FILE.rf[13][28] ;
 wire \u_cpu.REG_FILE.rf[13][29] ;
 wire \u_cpu.REG_FILE.rf[13][2] ;
 wire \u_cpu.REG_FILE.rf[13][30] ;
 wire \u_cpu.REG_FILE.rf[13][31] ;
 wire \u_cpu.REG_FILE.rf[13][3] ;
 wire \u_cpu.REG_FILE.rf[13][4] ;
 wire \u_cpu.REG_FILE.rf[13][5] ;
 wire \u_cpu.REG_FILE.rf[13][6] ;
 wire \u_cpu.REG_FILE.rf[13][7] ;
 wire \u_cpu.REG_FILE.rf[13][8] ;
 wire \u_cpu.REG_FILE.rf[13][9] ;
 wire \u_cpu.REG_FILE.rf[14][0] ;
 wire \u_cpu.REG_FILE.rf[14][10] ;
 wire \u_cpu.REG_FILE.rf[14][11] ;
 wire \u_cpu.REG_FILE.rf[14][12] ;
 wire \u_cpu.REG_FILE.rf[14][13] ;
 wire \u_cpu.REG_FILE.rf[14][14] ;
 wire \u_cpu.REG_FILE.rf[14][15] ;
 wire \u_cpu.REG_FILE.rf[14][16] ;
 wire \u_cpu.REG_FILE.rf[14][17] ;
 wire \u_cpu.REG_FILE.rf[14][18] ;
 wire \u_cpu.REG_FILE.rf[14][19] ;
 wire \u_cpu.REG_FILE.rf[14][1] ;
 wire \u_cpu.REG_FILE.rf[14][20] ;
 wire \u_cpu.REG_FILE.rf[14][21] ;
 wire \u_cpu.REG_FILE.rf[14][22] ;
 wire \u_cpu.REG_FILE.rf[14][23] ;
 wire \u_cpu.REG_FILE.rf[14][24] ;
 wire \u_cpu.REG_FILE.rf[14][25] ;
 wire \u_cpu.REG_FILE.rf[14][26] ;
 wire \u_cpu.REG_FILE.rf[14][27] ;
 wire \u_cpu.REG_FILE.rf[14][28] ;
 wire \u_cpu.REG_FILE.rf[14][29] ;
 wire \u_cpu.REG_FILE.rf[14][2] ;
 wire \u_cpu.REG_FILE.rf[14][30] ;
 wire \u_cpu.REG_FILE.rf[14][31] ;
 wire \u_cpu.REG_FILE.rf[14][3] ;
 wire \u_cpu.REG_FILE.rf[14][4] ;
 wire \u_cpu.REG_FILE.rf[14][5] ;
 wire \u_cpu.REG_FILE.rf[14][6] ;
 wire \u_cpu.REG_FILE.rf[14][7] ;
 wire \u_cpu.REG_FILE.rf[14][8] ;
 wire \u_cpu.REG_FILE.rf[14][9] ;
 wire \u_cpu.REG_FILE.rf[15][0] ;
 wire \u_cpu.REG_FILE.rf[15][10] ;
 wire \u_cpu.REG_FILE.rf[15][11] ;
 wire \u_cpu.REG_FILE.rf[15][12] ;
 wire \u_cpu.REG_FILE.rf[15][13] ;
 wire \u_cpu.REG_FILE.rf[15][14] ;
 wire \u_cpu.REG_FILE.rf[15][15] ;
 wire \u_cpu.REG_FILE.rf[15][16] ;
 wire \u_cpu.REG_FILE.rf[15][17] ;
 wire \u_cpu.REG_FILE.rf[15][18] ;
 wire \u_cpu.REG_FILE.rf[15][19] ;
 wire \u_cpu.REG_FILE.rf[15][1] ;
 wire \u_cpu.REG_FILE.rf[15][20] ;
 wire \u_cpu.REG_FILE.rf[15][21] ;
 wire \u_cpu.REG_FILE.rf[15][22] ;
 wire \u_cpu.REG_FILE.rf[15][23] ;
 wire \u_cpu.REG_FILE.rf[15][24] ;
 wire \u_cpu.REG_FILE.rf[15][25] ;
 wire \u_cpu.REG_FILE.rf[15][26] ;
 wire \u_cpu.REG_FILE.rf[15][27] ;
 wire \u_cpu.REG_FILE.rf[15][28] ;
 wire \u_cpu.REG_FILE.rf[15][29] ;
 wire \u_cpu.REG_FILE.rf[15][2] ;
 wire \u_cpu.REG_FILE.rf[15][30] ;
 wire \u_cpu.REG_FILE.rf[15][31] ;
 wire \u_cpu.REG_FILE.rf[15][3] ;
 wire \u_cpu.REG_FILE.rf[15][4] ;
 wire \u_cpu.REG_FILE.rf[15][5] ;
 wire \u_cpu.REG_FILE.rf[15][6] ;
 wire \u_cpu.REG_FILE.rf[15][7] ;
 wire \u_cpu.REG_FILE.rf[15][8] ;
 wire \u_cpu.REG_FILE.rf[15][9] ;
 wire \u_cpu.REG_FILE.rf[16][0] ;
 wire \u_cpu.REG_FILE.rf[16][10] ;
 wire \u_cpu.REG_FILE.rf[16][11] ;
 wire \u_cpu.REG_FILE.rf[16][12] ;
 wire \u_cpu.REG_FILE.rf[16][13] ;
 wire \u_cpu.REG_FILE.rf[16][14] ;
 wire \u_cpu.REG_FILE.rf[16][15] ;
 wire \u_cpu.REG_FILE.rf[16][16] ;
 wire \u_cpu.REG_FILE.rf[16][17] ;
 wire \u_cpu.REG_FILE.rf[16][18] ;
 wire \u_cpu.REG_FILE.rf[16][19] ;
 wire \u_cpu.REG_FILE.rf[16][1] ;
 wire \u_cpu.REG_FILE.rf[16][20] ;
 wire \u_cpu.REG_FILE.rf[16][21] ;
 wire \u_cpu.REG_FILE.rf[16][22] ;
 wire \u_cpu.REG_FILE.rf[16][23] ;
 wire \u_cpu.REG_FILE.rf[16][24] ;
 wire \u_cpu.REG_FILE.rf[16][25] ;
 wire \u_cpu.REG_FILE.rf[16][26] ;
 wire \u_cpu.REG_FILE.rf[16][27] ;
 wire \u_cpu.REG_FILE.rf[16][28] ;
 wire \u_cpu.REG_FILE.rf[16][29] ;
 wire \u_cpu.REG_FILE.rf[16][2] ;
 wire \u_cpu.REG_FILE.rf[16][30] ;
 wire \u_cpu.REG_FILE.rf[16][31] ;
 wire \u_cpu.REG_FILE.rf[16][3] ;
 wire \u_cpu.REG_FILE.rf[16][4] ;
 wire \u_cpu.REG_FILE.rf[16][5] ;
 wire \u_cpu.REG_FILE.rf[16][6] ;
 wire \u_cpu.REG_FILE.rf[16][7] ;
 wire \u_cpu.REG_FILE.rf[16][8] ;
 wire \u_cpu.REG_FILE.rf[16][9] ;
 wire \u_cpu.REG_FILE.rf[17][0] ;
 wire \u_cpu.REG_FILE.rf[17][10] ;
 wire \u_cpu.REG_FILE.rf[17][11] ;
 wire \u_cpu.REG_FILE.rf[17][12] ;
 wire \u_cpu.REG_FILE.rf[17][13] ;
 wire \u_cpu.REG_FILE.rf[17][14] ;
 wire \u_cpu.REG_FILE.rf[17][15] ;
 wire \u_cpu.REG_FILE.rf[17][16] ;
 wire \u_cpu.REG_FILE.rf[17][17] ;
 wire \u_cpu.REG_FILE.rf[17][18] ;
 wire \u_cpu.REG_FILE.rf[17][19] ;
 wire \u_cpu.REG_FILE.rf[17][1] ;
 wire \u_cpu.REG_FILE.rf[17][20] ;
 wire \u_cpu.REG_FILE.rf[17][21] ;
 wire \u_cpu.REG_FILE.rf[17][22] ;
 wire \u_cpu.REG_FILE.rf[17][23] ;
 wire \u_cpu.REG_FILE.rf[17][24] ;
 wire \u_cpu.REG_FILE.rf[17][25] ;
 wire \u_cpu.REG_FILE.rf[17][26] ;
 wire \u_cpu.REG_FILE.rf[17][27] ;
 wire \u_cpu.REG_FILE.rf[17][28] ;
 wire \u_cpu.REG_FILE.rf[17][29] ;
 wire \u_cpu.REG_FILE.rf[17][2] ;
 wire \u_cpu.REG_FILE.rf[17][30] ;
 wire \u_cpu.REG_FILE.rf[17][31] ;
 wire \u_cpu.REG_FILE.rf[17][3] ;
 wire \u_cpu.REG_FILE.rf[17][4] ;
 wire \u_cpu.REG_FILE.rf[17][5] ;
 wire \u_cpu.REG_FILE.rf[17][6] ;
 wire \u_cpu.REG_FILE.rf[17][7] ;
 wire \u_cpu.REG_FILE.rf[17][8] ;
 wire \u_cpu.REG_FILE.rf[17][9] ;
 wire \u_cpu.REG_FILE.rf[18][0] ;
 wire \u_cpu.REG_FILE.rf[18][10] ;
 wire \u_cpu.REG_FILE.rf[18][11] ;
 wire \u_cpu.REG_FILE.rf[18][12] ;
 wire \u_cpu.REG_FILE.rf[18][13] ;
 wire \u_cpu.REG_FILE.rf[18][14] ;
 wire \u_cpu.REG_FILE.rf[18][15] ;
 wire \u_cpu.REG_FILE.rf[18][16] ;
 wire \u_cpu.REG_FILE.rf[18][17] ;
 wire \u_cpu.REG_FILE.rf[18][18] ;
 wire \u_cpu.REG_FILE.rf[18][19] ;
 wire \u_cpu.REG_FILE.rf[18][1] ;
 wire \u_cpu.REG_FILE.rf[18][20] ;
 wire \u_cpu.REG_FILE.rf[18][21] ;
 wire \u_cpu.REG_FILE.rf[18][22] ;
 wire \u_cpu.REG_FILE.rf[18][23] ;
 wire \u_cpu.REG_FILE.rf[18][24] ;
 wire \u_cpu.REG_FILE.rf[18][25] ;
 wire \u_cpu.REG_FILE.rf[18][26] ;
 wire \u_cpu.REG_FILE.rf[18][27] ;
 wire \u_cpu.REG_FILE.rf[18][28] ;
 wire \u_cpu.REG_FILE.rf[18][29] ;
 wire \u_cpu.REG_FILE.rf[18][2] ;
 wire \u_cpu.REG_FILE.rf[18][30] ;
 wire \u_cpu.REG_FILE.rf[18][31] ;
 wire \u_cpu.REG_FILE.rf[18][3] ;
 wire \u_cpu.REG_FILE.rf[18][4] ;
 wire \u_cpu.REG_FILE.rf[18][5] ;
 wire \u_cpu.REG_FILE.rf[18][6] ;
 wire \u_cpu.REG_FILE.rf[18][7] ;
 wire \u_cpu.REG_FILE.rf[18][8] ;
 wire \u_cpu.REG_FILE.rf[18][9] ;
 wire \u_cpu.REG_FILE.rf[19][0] ;
 wire \u_cpu.REG_FILE.rf[19][10] ;
 wire \u_cpu.REG_FILE.rf[19][11] ;
 wire \u_cpu.REG_FILE.rf[19][12] ;
 wire \u_cpu.REG_FILE.rf[19][13] ;
 wire \u_cpu.REG_FILE.rf[19][14] ;
 wire \u_cpu.REG_FILE.rf[19][15] ;
 wire \u_cpu.REG_FILE.rf[19][16] ;
 wire \u_cpu.REG_FILE.rf[19][17] ;
 wire \u_cpu.REG_FILE.rf[19][18] ;
 wire \u_cpu.REG_FILE.rf[19][19] ;
 wire \u_cpu.REG_FILE.rf[19][1] ;
 wire \u_cpu.REG_FILE.rf[19][20] ;
 wire \u_cpu.REG_FILE.rf[19][21] ;
 wire \u_cpu.REG_FILE.rf[19][22] ;
 wire \u_cpu.REG_FILE.rf[19][23] ;
 wire \u_cpu.REG_FILE.rf[19][24] ;
 wire \u_cpu.REG_FILE.rf[19][25] ;
 wire \u_cpu.REG_FILE.rf[19][26] ;
 wire \u_cpu.REG_FILE.rf[19][27] ;
 wire \u_cpu.REG_FILE.rf[19][28] ;
 wire \u_cpu.REG_FILE.rf[19][29] ;
 wire \u_cpu.REG_FILE.rf[19][2] ;
 wire \u_cpu.REG_FILE.rf[19][30] ;
 wire \u_cpu.REG_FILE.rf[19][31] ;
 wire \u_cpu.REG_FILE.rf[19][3] ;
 wire \u_cpu.REG_FILE.rf[19][4] ;
 wire \u_cpu.REG_FILE.rf[19][5] ;
 wire \u_cpu.REG_FILE.rf[19][6] ;
 wire \u_cpu.REG_FILE.rf[19][7] ;
 wire \u_cpu.REG_FILE.rf[19][8] ;
 wire \u_cpu.REG_FILE.rf[19][9] ;
 wire \u_cpu.REG_FILE.rf[1][0] ;
 wire \u_cpu.REG_FILE.rf[1][10] ;
 wire \u_cpu.REG_FILE.rf[1][11] ;
 wire \u_cpu.REG_FILE.rf[1][12] ;
 wire \u_cpu.REG_FILE.rf[1][13] ;
 wire \u_cpu.REG_FILE.rf[1][14] ;
 wire \u_cpu.REG_FILE.rf[1][15] ;
 wire \u_cpu.REG_FILE.rf[1][16] ;
 wire \u_cpu.REG_FILE.rf[1][17] ;
 wire \u_cpu.REG_FILE.rf[1][18] ;
 wire \u_cpu.REG_FILE.rf[1][19] ;
 wire \u_cpu.REG_FILE.rf[1][1] ;
 wire \u_cpu.REG_FILE.rf[1][20] ;
 wire \u_cpu.REG_FILE.rf[1][21] ;
 wire \u_cpu.REG_FILE.rf[1][22] ;
 wire \u_cpu.REG_FILE.rf[1][23] ;
 wire \u_cpu.REG_FILE.rf[1][24] ;
 wire \u_cpu.REG_FILE.rf[1][25] ;
 wire \u_cpu.REG_FILE.rf[1][26] ;
 wire \u_cpu.REG_FILE.rf[1][27] ;
 wire \u_cpu.REG_FILE.rf[1][28] ;
 wire \u_cpu.REG_FILE.rf[1][29] ;
 wire \u_cpu.REG_FILE.rf[1][2] ;
 wire \u_cpu.REG_FILE.rf[1][30] ;
 wire \u_cpu.REG_FILE.rf[1][31] ;
 wire \u_cpu.REG_FILE.rf[1][3] ;
 wire \u_cpu.REG_FILE.rf[1][4] ;
 wire \u_cpu.REG_FILE.rf[1][5] ;
 wire \u_cpu.REG_FILE.rf[1][6] ;
 wire \u_cpu.REG_FILE.rf[1][7] ;
 wire \u_cpu.REG_FILE.rf[1][8] ;
 wire \u_cpu.REG_FILE.rf[1][9] ;
 wire \u_cpu.REG_FILE.rf[20][0] ;
 wire \u_cpu.REG_FILE.rf[20][10] ;
 wire \u_cpu.REG_FILE.rf[20][11] ;
 wire \u_cpu.REG_FILE.rf[20][12] ;
 wire \u_cpu.REG_FILE.rf[20][13] ;
 wire \u_cpu.REG_FILE.rf[20][14] ;
 wire \u_cpu.REG_FILE.rf[20][15] ;
 wire \u_cpu.REG_FILE.rf[20][16] ;
 wire \u_cpu.REG_FILE.rf[20][17] ;
 wire \u_cpu.REG_FILE.rf[20][18] ;
 wire \u_cpu.REG_FILE.rf[20][19] ;
 wire \u_cpu.REG_FILE.rf[20][1] ;
 wire \u_cpu.REG_FILE.rf[20][20] ;
 wire \u_cpu.REG_FILE.rf[20][21] ;
 wire \u_cpu.REG_FILE.rf[20][22] ;
 wire \u_cpu.REG_FILE.rf[20][23] ;
 wire \u_cpu.REG_FILE.rf[20][24] ;
 wire \u_cpu.REG_FILE.rf[20][25] ;
 wire \u_cpu.REG_FILE.rf[20][26] ;
 wire \u_cpu.REG_FILE.rf[20][27] ;
 wire \u_cpu.REG_FILE.rf[20][28] ;
 wire \u_cpu.REG_FILE.rf[20][29] ;
 wire \u_cpu.REG_FILE.rf[20][2] ;
 wire \u_cpu.REG_FILE.rf[20][30] ;
 wire \u_cpu.REG_FILE.rf[20][31] ;
 wire \u_cpu.REG_FILE.rf[20][3] ;
 wire \u_cpu.REG_FILE.rf[20][4] ;
 wire \u_cpu.REG_FILE.rf[20][5] ;
 wire \u_cpu.REG_FILE.rf[20][6] ;
 wire \u_cpu.REG_FILE.rf[20][7] ;
 wire \u_cpu.REG_FILE.rf[20][8] ;
 wire \u_cpu.REG_FILE.rf[20][9] ;
 wire \u_cpu.REG_FILE.rf[21][0] ;
 wire \u_cpu.REG_FILE.rf[21][10] ;
 wire \u_cpu.REG_FILE.rf[21][11] ;
 wire \u_cpu.REG_FILE.rf[21][12] ;
 wire \u_cpu.REG_FILE.rf[21][13] ;
 wire \u_cpu.REG_FILE.rf[21][14] ;
 wire \u_cpu.REG_FILE.rf[21][15] ;
 wire \u_cpu.REG_FILE.rf[21][16] ;
 wire \u_cpu.REG_FILE.rf[21][17] ;
 wire \u_cpu.REG_FILE.rf[21][18] ;
 wire \u_cpu.REG_FILE.rf[21][19] ;
 wire \u_cpu.REG_FILE.rf[21][1] ;
 wire \u_cpu.REG_FILE.rf[21][20] ;
 wire \u_cpu.REG_FILE.rf[21][21] ;
 wire \u_cpu.REG_FILE.rf[21][22] ;
 wire \u_cpu.REG_FILE.rf[21][23] ;
 wire \u_cpu.REG_FILE.rf[21][24] ;
 wire \u_cpu.REG_FILE.rf[21][25] ;
 wire \u_cpu.REG_FILE.rf[21][26] ;
 wire \u_cpu.REG_FILE.rf[21][27] ;
 wire \u_cpu.REG_FILE.rf[21][28] ;
 wire \u_cpu.REG_FILE.rf[21][29] ;
 wire \u_cpu.REG_FILE.rf[21][2] ;
 wire \u_cpu.REG_FILE.rf[21][30] ;
 wire \u_cpu.REG_FILE.rf[21][31] ;
 wire \u_cpu.REG_FILE.rf[21][3] ;
 wire \u_cpu.REG_FILE.rf[21][4] ;
 wire \u_cpu.REG_FILE.rf[21][5] ;
 wire \u_cpu.REG_FILE.rf[21][6] ;
 wire \u_cpu.REG_FILE.rf[21][7] ;
 wire \u_cpu.REG_FILE.rf[21][8] ;
 wire \u_cpu.REG_FILE.rf[21][9] ;
 wire \u_cpu.REG_FILE.rf[22][0] ;
 wire \u_cpu.REG_FILE.rf[22][10] ;
 wire \u_cpu.REG_FILE.rf[22][11] ;
 wire \u_cpu.REG_FILE.rf[22][12] ;
 wire \u_cpu.REG_FILE.rf[22][13] ;
 wire \u_cpu.REG_FILE.rf[22][14] ;
 wire \u_cpu.REG_FILE.rf[22][15] ;
 wire \u_cpu.REG_FILE.rf[22][16] ;
 wire \u_cpu.REG_FILE.rf[22][17] ;
 wire \u_cpu.REG_FILE.rf[22][18] ;
 wire \u_cpu.REG_FILE.rf[22][19] ;
 wire \u_cpu.REG_FILE.rf[22][1] ;
 wire \u_cpu.REG_FILE.rf[22][20] ;
 wire \u_cpu.REG_FILE.rf[22][21] ;
 wire \u_cpu.REG_FILE.rf[22][22] ;
 wire \u_cpu.REG_FILE.rf[22][23] ;
 wire \u_cpu.REG_FILE.rf[22][24] ;
 wire \u_cpu.REG_FILE.rf[22][25] ;
 wire \u_cpu.REG_FILE.rf[22][26] ;
 wire \u_cpu.REG_FILE.rf[22][27] ;
 wire \u_cpu.REG_FILE.rf[22][28] ;
 wire \u_cpu.REG_FILE.rf[22][29] ;
 wire \u_cpu.REG_FILE.rf[22][2] ;
 wire \u_cpu.REG_FILE.rf[22][30] ;
 wire \u_cpu.REG_FILE.rf[22][31] ;
 wire \u_cpu.REG_FILE.rf[22][3] ;
 wire \u_cpu.REG_FILE.rf[22][4] ;
 wire \u_cpu.REG_FILE.rf[22][5] ;
 wire \u_cpu.REG_FILE.rf[22][6] ;
 wire \u_cpu.REG_FILE.rf[22][7] ;
 wire \u_cpu.REG_FILE.rf[22][8] ;
 wire \u_cpu.REG_FILE.rf[22][9] ;
 wire \u_cpu.REG_FILE.rf[23][0] ;
 wire \u_cpu.REG_FILE.rf[23][10] ;
 wire \u_cpu.REG_FILE.rf[23][11] ;
 wire \u_cpu.REG_FILE.rf[23][12] ;
 wire \u_cpu.REG_FILE.rf[23][13] ;
 wire \u_cpu.REG_FILE.rf[23][14] ;
 wire \u_cpu.REG_FILE.rf[23][15] ;
 wire \u_cpu.REG_FILE.rf[23][16] ;
 wire \u_cpu.REG_FILE.rf[23][17] ;
 wire \u_cpu.REG_FILE.rf[23][18] ;
 wire \u_cpu.REG_FILE.rf[23][19] ;
 wire \u_cpu.REG_FILE.rf[23][1] ;
 wire \u_cpu.REG_FILE.rf[23][20] ;
 wire \u_cpu.REG_FILE.rf[23][21] ;
 wire \u_cpu.REG_FILE.rf[23][22] ;
 wire \u_cpu.REG_FILE.rf[23][23] ;
 wire \u_cpu.REG_FILE.rf[23][24] ;
 wire \u_cpu.REG_FILE.rf[23][25] ;
 wire \u_cpu.REG_FILE.rf[23][26] ;
 wire \u_cpu.REG_FILE.rf[23][27] ;
 wire \u_cpu.REG_FILE.rf[23][28] ;
 wire \u_cpu.REG_FILE.rf[23][29] ;
 wire \u_cpu.REG_FILE.rf[23][2] ;
 wire \u_cpu.REG_FILE.rf[23][30] ;
 wire \u_cpu.REG_FILE.rf[23][31] ;
 wire \u_cpu.REG_FILE.rf[23][3] ;
 wire \u_cpu.REG_FILE.rf[23][4] ;
 wire \u_cpu.REG_FILE.rf[23][5] ;
 wire \u_cpu.REG_FILE.rf[23][6] ;
 wire \u_cpu.REG_FILE.rf[23][7] ;
 wire \u_cpu.REG_FILE.rf[23][8] ;
 wire \u_cpu.REG_FILE.rf[23][9] ;
 wire \u_cpu.REG_FILE.rf[24][0] ;
 wire \u_cpu.REG_FILE.rf[24][10] ;
 wire \u_cpu.REG_FILE.rf[24][11] ;
 wire \u_cpu.REG_FILE.rf[24][12] ;
 wire \u_cpu.REG_FILE.rf[24][13] ;
 wire \u_cpu.REG_FILE.rf[24][14] ;
 wire \u_cpu.REG_FILE.rf[24][15] ;
 wire \u_cpu.REG_FILE.rf[24][16] ;
 wire \u_cpu.REG_FILE.rf[24][17] ;
 wire \u_cpu.REG_FILE.rf[24][18] ;
 wire \u_cpu.REG_FILE.rf[24][19] ;
 wire \u_cpu.REG_FILE.rf[24][1] ;
 wire \u_cpu.REG_FILE.rf[24][20] ;
 wire \u_cpu.REG_FILE.rf[24][21] ;
 wire \u_cpu.REG_FILE.rf[24][22] ;
 wire \u_cpu.REG_FILE.rf[24][23] ;
 wire \u_cpu.REG_FILE.rf[24][24] ;
 wire \u_cpu.REG_FILE.rf[24][25] ;
 wire \u_cpu.REG_FILE.rf[24][26] ;
 wire \u_cpu.REG_FILE.rf[24][27] ;
 wire \u_cpu.REG_FILE.rf[24][28] ;
 wire \u_cpu.REG_FILE.rf[24][29] ;
 wire \u_cpu.REG_FILE.rf[24][2] ;
 wire \u_cpu.REG_FILE.rf[24][30] ;
 wire \u_cpu.REG_FILE.rf[24][31] ;
 wire \u_cpu.REG_FILE.rf[24][3] ;
 wire \u_cpu.REG_FILE.rf[24][4] ;
 wire \u_cpu.REG_FILE.rf[24][5] ;
 wire \u_cpu.REG_FILE.rf[24][6] ;
 wire \u_cpu.REG_FILE.rf[24][7] ;
 wire \u_cpu.REG_FILE.rf[24][8] ;
 wire \u_cpu.REG_FILE.rf[24][9] ;
 wire \u_cpu.REG_FILE.rf[25][0] ;
 wire \u_cpu.REG_FILE.rf[25][10] ;
 wire \u_cpu.REG_FILE.rf[25][11] ;
 wire \u_cpu.REG_FILE.rf[25][12] ;
 wire \u_cpu.REG_FILE.rf[25][13] ;
 wire \u_cpu.REG_FILE.rf[25][14] ;
 wire \u_cpu.REG_FILE.rf[25][15] ;
 wire \u_cpu.REG_FILE.rf[25][16] ;
 wire \u_cpu.REG_FILE.rf[25][17] ;
 wire \u_cpu.REG_FILE.rf[25][18] ;
 wire \u_cpu.REG_FILE.rf[25][19] ;
 wire \u_cpu.REG_FILE.rf[25][1] ;
 wire \u_cpu.REG_FILE.rf[25][20] ;
 wire \u_cpu.REG_FILE.rf[25][21] ;
 wire \u_cpu.REG_FILE.rf[25][22] ;
 wire \u_cpu.REG_FILE.rf[25][23] ;
 wire \u_cpu.REG_FILE.rf[25][24] ;
 wire \u_cpu.REG_FILE.rf[25][25] ;
 wire \u_cpu.REG_FILE.rf[25][26] ;
 wire \u_cpu.REG_FILE.rf[25][27] ;
 wire \u_cpu.REG_FILE.rf[25][28] ;
 wire \u_cpu.REG_FILE.rf[25][29] ;
 wire \u_cpu.REG_FILE.rf[25][2] ;
 wire \u_cpu.REG_FILE.rf[25][30] ;
 wire \u_cpu.REG_FILE.rf[25][31] ;
 wire \u_cpu.REG_FILE.rf[25][3] ;
 wire \u_cpu.REG_FILE.rf[25][4] ;
 wire \u_cpu.REG_FILE.rf[25][5] ;
 wire \u_cpu.REG_FILE.rf[25][6] ;
 wire \u_cpu.REG_FILE.rf[25][7] ;
 wire \u_cpu.REG_FILE.rf[25][8] ;
 wire \u_cpu.REG_FILE.rf[25][9] ;
 wire \u_cpu.REG_FILE.rf[26][0] ;
 wire \u_cpu.REG_FILE.rf[26][10] ;
 wire \u_cpu.REG_FILE.rf[26][11] ;
 wire \u_cpu.REG_FILE.rf[26][12] ;
 wire \u_cpu.REG_FILE.rf[26][13] ;
 wire \u_cpu.REG_FILE.rf[26][14] ;
 wire \u_cpu.REG_FILE.rf[26][15] ;
 wire \u_cpu.REG_FILE.rf[26][16] ;
 wire \u_cpu.REG_FILE.rf[26][17] ;
 wire \u_cpu.REG_FILE.rf[26][18] ;
 wire \u_cpu.REG_FILE.rf[26][19] ;
 wire \u_cpu.REG_FILE.rf[26][1] ;
 wire \u_cpu.REG_FILE.rf[26][20] ;
 wire \u_cpu.REG_FILE.rf[26][21] ;
 wire \u_cpu.REG_FILE.rf[26][22] ;
 wire \u_cpu.REG_FILE.rf[26][23] ;
 wire \u_cpu.REG_FILE.rf[26][24] ;
 wire \u_cpu.REG_FILE.rf[26][25] ;
 wire \u_cpu.REG_FILE.rf[26][26] ;
 wire \u_cpu.REG_FILE.rf[26][27] ;
 wire \u_cpu.REG_FILE.rf[26][28] ;
 wire \u_cpu.REG_FILE.rf[26][29] ;
 wire \u_cpu.REG_FILE.rf[26][2] ;
 wire \u_cpu.REG_FILE.rf[26][30] ;
 wire \u_cpu.REG_FILE.rf[26][31] ;
 wire \u_cpu.REG_FILE.rf[26][3] ;
 wire \u_cpu.REG_FILE.rf[26][4] ;
 wire \u_cpu.REG_FILE.rf[26][5] ;
 wire \u_cpu.REG_FILE.rf[26][6] ;
 wire \u_cpu.REG_FILE.rf[26][7] ;
 wire \u_cpu.REG_FILE.rf[26][8] ;
 wire \u_cpu.REG_FILE.rf[26][9] ;
 wire \u_cpu.REG_FILE.rf[27][0] ;
 wire \u_cpu.REG_FILE.rf[27][10] ;
 wire \u_cpu.REG_FILE.rf[27][11] ;
 wire \u_cpu.REG_FILE.rf[27][12] ;
 wire \u_cpu.REG_FILE.rf[27][13] ;
 wire \u_cpu.REG_FILE.rf[27][14] ;
 wire \u_cpu.REG_FILE.rf[27][15] ;
 wire \u_cpu.REG_FILE.rf[27][16] ;
 wire \u_cpu.REG_FILE.rf[27][17] ;
 wire \u_cpu.REG_FILE.rf[27][18] ;
 wire \u_cpu.REG_FILE.rf[27][19] ;
 wire \u_cpu.REG_FILE.rf[27][1] ;
 wire \u_cpu.REG_FILE.rf[27][20] ;
 wire \u_cpu.REG_FILE.rf[27][21] ;
 wire \u_cpu.REG_FILE.rf[27][22] ;
 wire \u_cpu.REG_FILE.rf[27][23] ;
 wire \u_cpu.REG_FILE.rf[27][24] ;
 wire \u_cpu.REG_FILE.rf[27][25] ;
 wire \u_cpu.REG_FILE.rf[27][26] ;
 wire \u_cpu.REG_FILE.rf[27][27] ;
 wire \u_cpu.REG_FILE.rf[27][28] ;
 wire \u_cpu.REG_FILE.rf[27][29] ;
 wire \u_cpu.REG_FILE.rf[27][2] ;
 wire \u_cpu.REG_FILE.rf[27][30] ;
 wire \u_cpu.REG_FILE.rf[27][31] ;
 wire \u_cpu.REG_FILE.rf[27][3] ;
 wire \u_cpu.REG_FILE.rf[27][4] ;
 wire \u_cpu.REG_FILE.rf[27][5] ;
 wire \u_cpu.REG_FILE.rf[27][6] ;
 wire \u_cpu.REG_FILE.rf[27][7] ;
 wire \u_cpu.REG_FILE.rf[27][8] ;
 wire \u_cpu.REG_FILE.rf[27][9] ;
 wire \u_cpu.REG_FILE.rf[28][0] ;
 wire \u_cpu.REG_FILE.rf[28][10] ;
 wire \u_cpu.REG_FILE.rf[28][11] ;
 wire \u_cpu.REG_FILE.rf[28][12] ;
 wire \u_cpu.REG_FILE.rf[28][13] ;
 wire \u_cpu.REG_FILE.rf[28][14] ;
 wire \u_cpu.REG_FILE.rf[28][15] ;
 wire \u_cpu.REG_FILE.rf[28][16] ;
 wire \u_cpu.REG_FILE.rf[28][17] ;
 wire \u_cpu.REG_FILE.rf[28][18] ;
 wire \u_cpu.REG_FILE.rf[28][19] ;
 wire \u_cpu.REG_FILE.rf[28][1] ;
 wire \u_cpu.REG_FILE.rf[28][20] ;
 wire \u_cpu.REG_FILE.rf[28][21] ;
 wire \u_cpu.REG_FILE.rf[28][22] ;
 wire \u_cpu.REG_FILE.rf[28][23] ;
 wire \u_cpu.REG_FILE.rf[28][24] ;
 wire \u_cpu.REG_FILE.rf[28][25] ;
 wire \u_cpu.REG_FILE.rf[28][26] ;
 wire \u_cpu.REG_FILE.rf[28][27] ;
 wire \u_cpu.REG_FILE.rf[28][28] ;
 wire \u_cpu.REG_FILE.rf[28][29] ;
 wire \u_cpu.REG_FILE.rf[28][2] ;
 wire \u_cpu.REG_FILE.rf[28][30] ;
 wire \u_cpu.REG_FILE.rf[28][31] ;
 wire \u_cpu.REG_FILE.rf[28][3] ;
 wire \u_cpu.REG_FILE.rf[28][4] ;
 wire \u_cpu.REG_FILE.rf[28][5] ;
 wire \u_cpu.REG_FILE.rf[28][6] ;
 wire \u_cpu.REG_FILE.rf[28][7] ;
 wire \u_cpu.REG_FILE.rf[28][8] ;
 wire \u_cpu.REG_FILE.rf[28][9] ;
 wire \u_cpu.REG_FILE.rf[29][0] ;
 wire \u_cpu.REG_FILE.rf[29][10] ;
 wire \u_cpu.REG_FILE.rf[29][11] ;
 wire \u_cpu.REG_FILE.rf[29][12] ;
 wire \u_cpu.REG_FILE.rf[29][13] ;
 wire \u_cpu.REG_FILE.rf[29][14] ;
 wire \u_cpu.REG_FILE.rf[29][15] ;
 wire \u_cpu.REG_FILE.rf[29][16] ;
 wire \u_cpu.REG_FILE.rf[29][17] ;
 wire \u_cpu.REG_FILE.rf[29][18] ;
 wire \u_cpu.REG_FILE.rf[29][19] ;
 wire \u_cpu.REG_FILE.rf[29][1] ;
 wire \u_cpu.REG_FILE.rf[29][20] ;
 wire \u_cpu.REG_FILE.rf[29][21] ;
 wire \u_cpu.REG_FILE.rf[29][22] ;
 wire \u_cpu.REG_FILE.rf[29][23] ;
 wire \u_cpu.REG_FILE.rf[29][24] ;
 wire \u_cpu.REG_FILE.rf[29][25] ;
 wire \u_cpu.REG_FILE.rf[29][26] ;
 wire \u_cpu.REG_FILE.rf[29][27] ;
 wire \u_cpu.REG_FILE.rf[29][28] ;
 wire \u_cpu.REG_FILE.rf[29][29] ;
 wire \u_cpu.REG_FILE.rf[29][2] ;
 wire \u_cpu.REG_FILE.rf[29][30] ;
 wire \u_cpu.REG_FILE.rf[29][31] ;
 wire \u_cpu.REG_FILE.rf[29][3] ;
 wire \u_cpu.REG_FILE.rf[29][4] ;
 wire \u_cpu.REG_FILE.rf[29][5] ;
 wire \u_cpu.REG_FILE.rf[29][6] ;
 wire \u_cpu.REG_FILE.rf[29][7] ;
 wire \u_cpu.REG_FILE.rf[29][8] ;
 wire \u_cpu.REG_FILE.rf[29][9] ;
 wire \u_cpu.REG_FILE.rf[2][0] ;
 wire \u_cpu.REG_FILE.rf[2][10] ;
 wire \u_cpu.REG_FILE.rf[2][11] ;
 wire \u_cpu.REG_FILE.rf[2][12] ;
 wire \u_cpu.REG_FILE.rf[2][13] ;
 wire \u_cpu.REG_FILE.rf[2][14] ;
 wire \u_cpu.REG_FILE.rf[2][15] ;
 wire \u_cpu.REG_FILE.rf[2][16] ;
 wire \u_cpu.REG_FILE.rf[2][17] ;
 wire \u_cpu.REG_FILE.rf[2][18] ;
 wire \u_cpu.REG_FILE.rf[2][19] ;
 wire \u_cpu.REG_FILE.rf[2][1] ;
 wire \u_cpu.REG_FILE.rf[2][20] ;
 wire \u_cpu.REG_FILE.rf[2][21] ;
 wire \u_cpu.REG_FILE.rf[2][22] ;
 wire \u_cpu.REG_FILE.rf[2][23] ;
 wire \u_cpu.REG_FILE.rf[2][24] ;
 wire \u_cpu.REG_FILE.rf[2][25] ;
 wire \u_cpu.REG_FILE.rf[2][26] ;
 wire \u_cpu.REG_FILE.rf[2][27] ;
 wire \u_cpu.REG_FILE.rf[2][28] ;
 wire \u_cpu.REG_FILE.rf[2][29] ;
 wire \u_cpu.REG_FILE.rf[2][2] ;
 wire \u_cpu.REG_FILE.rf[2][30] ;
 wire \u_cpu.REG_FILE.rf[2][31] ;
 wire \u_cpu.REG_FILE.rf[2][3] ;
 wire \u_cpu.REG_FILE.rf[2][4] ;
 wire \u_cpu.REG_FILE.rf[2][5] ;
 wire \u_cpu.REG_FILE.rf[2][6] ;
 wire \u_cpu.REG_FILE.rf[2][7] ;
 wire \u_cpu.REG_FILE.rf[2][8] ;
 wire \u_cpu.REG_FILE.rf[2][9] ;
 wire \u_cpu.REG_FILE.rf[30][0] ;
 wire \u_cpu.REG_FILE.rf[30][10] ;
 wire \u_cpu.REG_FILE.rf[30][11] ;
 wire \u_cpu.REG_FILE.rf[30][12] ;
 wire \u_cpu.REG_FILE.rf[30][13] ;
 wire \u_cpu.REG_FILE.rf[30][14] ;
 wire \u_cpu.REG_FILE.rf[30][15] ;
 wire \u_cpu.REG_FILE.rf[30][16] ;
 wire \u_cpu.REG_FILE.rf[30][17] ;
 wire \u_cpu.REG_FILE.rf[30][18] ;
 wire \u_cpu.REG_FILE.rf[30][19] ;
 wire \u_cpu.REG_FILE.rf[30][1] ;
 wire \u_cpu.REG_FILE.rf[30][20] ;
 wire \u_cpu.REG_FILE.rf[30][21] ;
 wire \u_cpu.REG_FILE.rf[30][22] ;
 wire \u_cpu.REG_FILE.rf[30][23] ;
 wire \u_cpu.REG_FILE.rf[30][24] ;
 wire \u_cpu.REG_FILE.rf[30][25] ;
 wire \u_cpu.REG_FILE.rf[30][26] ;
 wire \u_cpu.REG_FILE.rf[30][27] ;
 wire \u_cpu.REG_FILE.rf[30][28] ;
 wire \u_cpu.REG_FILE.rf[30][29] ;
 wire \u_cpu.REG_FILE.rf[30][2] ;
 wire \u_cpu.REG_FILE.rf[30][30] ;
 wire \u_cpu.REG_FILE.rf[30][31] ;
 wire \u_cpu.REG_FILE.rf[30][3] ;
 wire \u_cpu.REG_FILE.rf[30][4] ;
 wire \u_cpu.REG_FILE.rf[30][5] ;
 wire \u_cpu.REG_FILE.rf[30][6] ;
 wire \u_cpu.REG_FILE.rf[30][7] ;
 wire \u_cpu.REG_FILE.rf[30][8] ;
 wire \u_cpu.REG_FILE.rf[30][9] ;
 wire \u_cpu.REG_FILE.rf[31][0] ;
 wire \u_cpu.REG_FILE.rf[31][10] ;
 wire \u_cpu.REG_FILE.rf[31][11] ;
 wire \u_cpu.REG_FILE.rf[31][12] ;
 wire \u_cpu.REG_FILE.rf[31][13] ;
 wire \u_cpu.REG_FILE.rf[31][14] ;
 wire \u_cpu.REG_FILE.rf[31][15] ;
 wire \u_cpu.REG_FILE.rf[31][16] ;
 wire \u_cpu.REG_FILE.rf[31][17] ;
 wire \u_cpu.REG_FILE.rf[31][18] ;
 wire \u_cpu.REG_FILE.rf[31][19] ;
 wire \u_cpu.REG_FILE.rf[31][1] ;
 wire \u_cpu.REG_FILE.rf[31][20] ;
 wire \u_cpu.REG_FILE.rf[31][21] ;
 wire \u_cpu.REG_FILE.rf[31][22] ;
 wire \u_cpu.REG_FILE.rf[31][23] ;
 wire \u_cpu.REG_FILE.rf[31][24] ;
 wire \u_cpu.REG_FILE.rf[31][25] ;
 wire \u_cpu.REG_FILE.rf[31][26] ;
 wire \u_cpu.REG_FILE.rf[31][27] ;
 wire \u_cpu.REG_FILE.rf[31][28] ;
 wire \u_cpu.REG_FILE.rf[31][29] ;
 wire \u_cpu.REG_FILE.rf[31][2] ;
 wire \u_cpu.REG_FILE.rf[31][30] ;
 wire \u_cpu.REG_FILE.rf[31][31] ;
 wire \u_cpu.REG_FILE.rf[31][3] ;
 wire \u_cpu.REG_FILE.rf[31][4] ;
 wire \u_cpu.REG_FILE.rf[31][5] ;
 wire \u_cpu.REG_FILE.rf[31][6] ;
 wire \u_cpu.REG_FILE.rf[31][7] ;
 wire \u_cpu.REG_FILE.rf[31][8] ;
 wire \u_cpu.REG_FILE.rf[31][9] ;
 wire \u_cpu.REG_FILE.rf[3][0] ;
 wire \u_cpu.REG_FILE.rf[3][10] ;
 wire \u_cpu.REG_FILE.rf[3][11] ;
 wire \u_cpu.REG_FILE.rf[3][12] ;
 wire \u_cpu.REG_FILE.rf[3][13] ;
 wire \u_cpu.REG_FILE.rf[3][14] ;
 wire \u_cpu.REG_FILE.rf[3][15] ;
 wire \u_cpu.REG_FILE.rf[3][16] ;
 wire \u_cpu.REG_FILE.rf[3][17] ;
 wire \u_cpu.REG_FILE.rf[3][18] ;
 wire \u_cpu.REG_FILE.rf[3][19] ;
 wire \u_cpu.REG_FILE.rf[3][1] ;
 wire \u_cpu.REG_FILE.rf[3][20] ;
 wire \u_cpu.REG_FILE.rf[3][21] ;
 wire \u_cpu.REG_FILE.rf[3][22] ;
 wire \u_cpu.REG_FILE.rf[3][23] ;
 wire \u_cpu.REG_FILE.rf[3][24] ;
 wire \u_cpu.REG_FILE.rf[3][25] ;
 wire \u_cpu.REG_FILE.rf[3][26] ;
 wire \u_cpu.REG_FILE.rf[3][27] ;
 wire \u_cpu.REG_FILE.rf[3][28] ;
 wire \u_cpu.REG_FILE.rf[3][29] ;
 wire \u_cpu.REG_FILE.rf[3][2] ;
 wire \u_cpu.REG_FILE.rf[3][30] ;
 wire \u_cpu.REG_FILE.rf[3][31] ;
 wire \u_cpu.REG_FILE.rf[3][3] ;
 wire \u_cpu.REG_FILE.rf[3][4] ;
 wire \u_cpu.REG_FILE.rf[3][5] ;
 wire \u_cpu.REG_FILE.rf[3][6] ;
 wire \u_cpu.REG_FILE.rf[3][7] ;
 wire \u_cpu.REG_FILE.rf[3][8] ;
 wire \u_cpu.REG_FILE.rf[3][9] ;
 wire \u_cpu.REG_FILE.rf[4][0] ;
 wire \u_cpu.REG_FILE.rf[4][10] ;
 wire \u_cpu.REG_FILE.rf[4][11] ;
 wire \u_cpu.REG_FILE.rf[4][12] ;
 wire \u_cpu.REG_FILE.rf[4][13] ;
 wire \u_cpu.REG_FILE.rf[4][14] ;
 wire \u_cpu.REG_FILE.rf[4][15] ;
 wire \u_cpu.REG_FILE.rf[4][16] ;
 wire \u_cpu.REG_FILE.rf[4][17] ;
 wire \u_cpu.REG_FILE.rf[4][18] ;
 wire \u_cpu.REG_FILE.rf[4][19] ;
 wire \u_cpu.REG_FILE.rf[4][1] ;
 wire \u_cpu.REG_FILE.rf[4][20] ;
 wire \u_cpu.REG_FILE.rf[4][21] ;
 wire \u_cpu.REG_FILE.rf[4][22] ;
 wire \u_cpu.REG_FILE.rf[4][23] ;
 wire \u_cpu.REG_FILE.rf[4][24] ;
 wire \u_cpu.REG_FILE.rf[4][25] ;
 wire \u_cpu.REG_FILE.rf[4][26] ;
 wire \u_cpu.REG_FILE.rf[4][27] ;
 wire \u_cpu.REG_FILE.rf[4][28] ;
 wire \u_cpu.REG_FILE.rf[4][29] ;
 wire \u_cpu.REG_FILE.rf[4][2] ;
 wire \u_cpu.REG_FILE.rf[4][30] ;
 wire \u_cpu.REG_FILE.rf[4][31] ;
 wire \u_cpu.REG_FILE.rf[4][3] ;
 wire \u_cpu.REG_FILE.rf[4][4] ;
 wire \u_cpu.REG_FILE.rf[4][5] ;
 wire \u_cpu.REG_FILE.rf[4][6] ;
 wire \u_cpu.REG_FILE.rf[4][7] ;
 wire \u_cpu.REG_FILE.rf[4][8] ;
 wire \u_cpu.REG_FILE.rf[4][9] ;
 wire \u_cpu.REG_FILE.rf[5][0] ;
 wire \u_cpu.REG_FILE.rf[5][10] ;
 wire \u_cpu.REG_FILE.rf[5][11] ;
 wire \u_cpu.REG_FILE.rf[5][12] ;
 wire \u_cpu.REG_FILE.rf[5][13] ;
 wire \u_cpu.REG_FILE.rf[5][14] ;
 wire \u_cpu.REG_FILE.rf[5][15] ;
 wire \u_cpu.REG_FILE.rf[5][16] ;
 wire \u_cpu.REG_FILE.rf[5][17] ;
 wire \u_cpu.REG_FILE.rf[5][18] ;
 wire \u_cpu.REG_FILE.rf[5][19] ;
 wire \u_cpu.REG_FILE.rf[5][1] ;
 wire \u_cpu.REG_FILE.rf[5][20] ;
 wire \u_cpu.REG_FILE.rf[5][21] ;
 wire \u_cpu.REG_FILE.rf[5][22] ;
 wire \u_cpu.REG_FILE.rf[5][23] ;
 wire \u_cpu.REG_FILE.rf[5][24] ;
 wire \u_cpu.REG_FILE.rf[5][25] ;
 wire \u_cpu.REG_FILE.rf[5][26] ;
 wire \u_cpu.REG_FILE.rf[5][27] ;
 wire \u_cpu.REG_FILE.rf[5][28] ;
 wire \u_cpu.REG_FILE.rf[5][29] ;
 wire \u_cpu.REG_FILE.rf[5][2] ;
 wire \u_cpu.REG_FILE.rf[5][30] ;
 wire \u_cpu.REG_FILE.rf[5][31] ;
 wire \u_cpu.REG_FILE.rf[5][3] ;
 wire \u_cpu.REG_FILE.rf[5][4] ;
 wire \u_cpu.REG_FILE.rf[5][5] ;
 wire \u_cpu.REG_FILE.rf[5][6] ;
 wire \u_cpu.REG_FILE.rf[5][7] ;
 wire \u_cpu.REG_FILE.rf[5][8] ;
 wire \u_cpu.REG_FILE.rf[5][9] ;
 wire \u_cpu.REG_FILE.rf[6][0] ;
 wire \u_cpu.REG_FILE.rf[6][10] ;
 wire \u_cpu.REG_FILE.rf[6][11] ;
 wire \u_cpu.REG_FILE.rf[6][12] ;
 wire \u_cpu.REG_FILE.rf[6][13] ;
 wire \u_cpu.REG_FILE.rf[6][14] ;
 wire \u_cpu.REG_FILE.rf[6][15] ;
 wire \u_cpu.REG_FILE.rf[6][16] ;
 wire \u_cpu.REG_FILE.rf[6][17] ;
 wire \u_cpu.REG_FILE.rf[6][18] ;
 wire \u_cpu.REG_FILE.rf[6][19] ;
 wire \u_cpu.REG_FILE.rf[6][1] ;
 wire \u_cpu.REG_FILE.rf[6][20] ;
 wire \u_cpu.REG_FILE.rf[6][21] ;
 wire \u_cpu.REG_FILE.rf[6][22] ;
 wire \u_cpu.REG_FILE.rf[6][23] ;
 wire \u_cpu.REG_FILE.rf[6][24] ;
 wire \u_cpu.REG_FILE.rf[6][25] ;
 wire \u_cpu.REG_FILE.rf[6][26] ;
 wire \u_cpu.REG_FILE.rf[6][27] ;
 wire \u_cpu.REG_FILE.rf[6][28] ;
 wire \u_cpu.REG_FILE.rf[6][29] ;
 wire \u_cpu.REG_FILE.rf[6][2] ;
 wire \u_cpu.REG_FILE.rf[6][30] ;
 wire \u_cpu.REG_FILE.rf[6][31] ;
 wire \u_cpu.REG_FILE.rf[6][3] ;
 wire \u_cpu.REG_FILE.rf[6][4] ;
 wire \u_cpu.REG_FILE.rf[6][5] ;
 wire \u_cpu.REG_FILE.rf[6][6] ;
 wire \u_cpu.REG_FILE.rf[6][7] ;
 wire \u_cpu.REG_FILE.rf[6][8] ;
 wire \u_cpu.REG_FILE.rf[6][9] ;
 wire \u_cpu.REG_FILE.rf[7][0] ;
 wire \u_cpu.REG_FILE.rf[7][10] ;
 wire \u_cpu.REG_FILE.rf[7][11] ;
 wire \u_cpu.REG_FILE.rf[7][12] ;
 wire \u_cpu.REG_FILE.rf[7][13] ;
 wire \u_cpu.REG_FILE.rf[7][14] ;
 wire \u_cpu.REG_FILE.rf[7][15] ;
 wire \u_cpu.REG_FILE.rf[7][16] ;
 wire \u_cpu.REG_FILE.rf[7][17] ;
 wire \u_cpu.REG_FILE.rf[7][18] ;
 wire \u_cpu.REG_FILE.rf[7][19] ;
 wire \u_cpu.REG_FILE.rf[7][1] ;
 wire \u_cpu.REG_FILE.rf[7][20] ;
 wire \u_cpu.REG_FILE.rf[7][21] ;
 wire \u_cpu.REG_FILE.rf[7][22] ;
 wire \u_cpu.REG_FILE.rf[7][23] ;
 wire \u_cpu.REG_FILE.rf[7][24] ;
 wire \u_cpu.REG_FILE.rf[7][25] ;
 wire \u_cpu.REG_FILE.rf[7][26] ;
 wire \u_cpu.REG_FILE.rf[7][27] ;
 wire \u_cpu.REG_FILE.rf[7][28] ;
 wire \u_cpu.REG_FILE.rf[7][29] ;
 wire \u_cpu.REG_FILE.rf[7][2] ;
 wire \u_cpu.REG_FILE.rf[7][30] ;
 wire \u_cpu.REG_FILE.rf[7][31] ;
 wire \u_cpu.REG_FILE.rf[7][3] ;
 wire \u_cpu.REG_FILE.rf[7][4] ;
 wire \u_cpu.REG_FILE.rf[7][5] ;
 wire \u_cpu.REG_FILE.rf[7][6] ;
 wire \u_cpu.REG_FILE.rf[7][7] ;
 wire \u_cpu.REG_FILE.rf[7][8] ;
 wire \u_cpu.REG_FILE.rf[7][9] ;
 wire \u_cpu.REG_FILE.rf[8][0] ;
 wire \u_cpu.REG_FILE.rf[8][10] ;
 wire \u_cpu.REG_FILE.rf[8][11] ;
 wire \u_cpu.REG_FILE.rf[8][12] ;
 wire \u_cpu.REG_FILE.rf[8][13] ;
 wire \u_cpu.REG_FILE.rf[8][14] ;
 wire \u_cpu.REG_FILE.rf[8][15] ;
 wire \u_cpu.REG_FILE.rf[8][16] ;
 wire \u_cpu.REG_FILE.rf[8][17] ;
 wire \u_cpu.REG_FILE.rf[8][18] ;
 wire \u_cpu.REG_FILE.rf[8][19] ;
 wire \u_cpu.REG_FILE.rf[8][1] ;
 wire \u_cpu.REG_FILE.rf[8][20] ;
 wire \u_cpu.REG_FILE.rf[8][21] ;
 wire \u_cpu.REG_FILE.rf[8][22] ;
 wire \u_cpu.REG_FILE.rf[8][23] ;
 wire \u_cpu.REG_FILE.rf[8][24] ;
 wire \u_cpu.REG_FILE.rf[8][25] ;
 wire \u_cpu.REG_FILE.rf[8][26] ;
 wire \u_cpu.REG_FILE.rf[8][27] ;
 wire \u_cpu.REG_FILE.rf[8][28] ;
 wire \u_cpu.REG_FILE.rf[8][29] ;
 wire \u_cpu.REG_FILE.rf[8][2] ;
 wire \u_cpu.REG_FILE.rf[8][30] ;
 wire \u_cpu.REG_FILE.rf[8][31] ;
 wire \u_cpu.REG_FILE.rf[8][3] ;
 wire \u_cpu.REG_FILE.rf[8][4] ;
 wire \u_cpu.REG_FILE.rf[8][5] ;
 wire \u_cpu.REG_FILE.rf[8][6] ;
 wire \u_cpu.REG_FILE.rf[8][7] ;
 wire \u_cpu.REG_FILE.rf[8][8] ;
 wire \u_cpu.REG_FILE.rf[8][9] ;
 wire \u_cpu.REG_FILE.rf[9][0] ;
 wire \u_cpu.REG_FILE.rf[9][10] ;
 wire \u_cpu.REG_FILE.rf[9][11] ;
 wire \u_cpu.REG_FILE.rf[9][12] ;
 wire \u_cpu.REG_FILE.rf[9][13] ;
 wire \u_cpu.REG_FILE.rf[9][14] ;
 wire \u_cpu.REG_FILE.rf[9][15] ;
 wire \u_cpu.REG_FILE.rf[9][16] ;
 wire \u_cpu.REG_FILE.rf[9][17] ;
 wire \u_cpu.REG_FILE.rf[9][18] ;
 wire \u_cpu.REG_FILE.rf[9][19] ;
 wire \u_cpu.REG_FILE.rf[9][1] ;
 wire \u_cpu.REG_FILE.rf[9][20] ;
 wire \u_cpu.REG_FILE.rf[9][21] ;
 wire \u_cpu.REG_FILE.rf[9][22] ;
 wire \u_cpu.REG_FILE.rf[9][23] ;
 wire \u_cpu.REG_FILE.rf[9][24] ;
 wire \u_cpu.REG_FILE.rf[9][25] ;
 wire \u_cpu.REG_FILE.rf[9][26] ;
 wire \u_cpu.REG_FILE.rf[9][27] ;
 wire \u_cpu.REG_FILE.rf[9][28] ;
 wire \u_cpu.REG_FILE.rf[9][29] ;
 wire \u_cpu.REG_FILE.rf[9][2] ;
 wire \u_cpu.REG_FILE.rf[9][30] ;
 wire \u_cpu.REG_FILE.rf[9][31] ;
 wire \u_cpu.REG_FILE.rf[9][3] ;
 wire \u_cpu.REG_FILE.rf[9][4] ;
 wire \u_cpu.REG_FILE.rf[9][5] ;
 wire \u_cpu.REG_FILE.rf[9][6] ;
 wire \u_cpu.REG_FILE.rf[9][7] ;
 wire \u_cpu.REG_FILE.rf[9][8] ;
 wire \u_cpu.REG_FILE.rf[9][9] ;
 wire \u_cpu.REG_FILE.wd3[0] ;
 wire \u_cpu.REG_FILE.wd3[10] ;
 wire \u_cpu.REG_FILE.wd3[11] ;
 wire \u_cpu.REG_FILE.wd3[12] ;
 wire \u_cpu.REG_FILE.wd3[13] ;
 wire \u_cpu.REG_FILE.wd3[14] ;
 wire \u_cpu.REG_FILE.wd3[15] ;
 wire \u_cpu.REG_FILE.wd3[16] ;
 wire \u_cpu.REG_FILE.wd3[17] ;
 wire \u_cpu.REG_FILE.wd3[18] ;
 wire \u_cpu.REG_FILE.wd3[19] ;
 wire \u_cpu.REG_FILE.wd3[1] ;
 wire \u_cpu.REG_FILE.wd3[20] ;
 wire \u_cpu.REG_FILE.wd3[21] ;
 wire \u_cpu.REG_FILE.wd3[22] ;
 wire \u_cpu.REG_FILE.wd3[23] ;
 wire \u_cpu.REG_FILE.wd3[24] ;
 wire \u_cpu.REG_FILE.wd3[25] ;
 wire \u_cpu.REG_FILE.wd3[26] ;
 wire \u_cpu.REG_FILE.wd3[27] ;
 wire \u_cpu.REG_FILE.wd3[28] ;
 wire \u_cpu.REG_FILE.wd3[29] ;
 wire \u_cpu.REG_FILE.wd3[2] ;
 wire \u_cpu.REG_FILE.wd3[30] ;
 wire \u_cpu.REG_FILE.wd3[31] ;
 wire \u_cpu.REG_FILE.wd3[3] ;
 wire \u_cpu.REG_FILE.wd3[4] ;
 wire \u_cpu.REG_FILE.wd3[5] ;
 wire \u_cpu.REG_FILE.wd3[6] ;
 wire \u_cpu.REG_FILE.wd3[7] ;
 wire \u_cpu.REG_FILE.wd3[8] ;
 wire \u_cpu.REG_FILE.wd3[9] ;
 wire \u_cpu.REG_FILE.we3 ;
 wire \u_cpu._0000_ ;
 wire \u_cpu._0001_ ;
 wire \u_cpu._0002_ ;
 wire \u_cpu._0003_ ;
 wire \u_cpu._0004_ ;
 wire \u_cpu._0005_ ;
 wire \u_cpu._0006_ ;
 wire \u_cpu._0007_ ;
 wire \u_cpu._0008_ ;
 wire \u_cpu._0009_ ;
 wire \u_cpu._0010_ ;
 wire \u_cpu._0011_ ;
 wire \u_cpu._0012_ ;
 wire \u_cpu._0013_ ;
 wire \u_cpu._0014_ ;
 wire \u_cpu._0015_ ;
 wire \u_cpu._0016_ ;
 wire \u_cpu._0017_ ;
 wire \u_cpu._0018_ ;
 wire \u_cpu._0019_ ;
 wire \u_cpu._0020_ ;
 wire \u_cpu._0021_ ;
 wire \u_cpu._0022_ ;
 wire \u_cpu._0023_ ;
 wire \u_cpu._0024_ ;
 wire \u_cpu._0025_ ;
 wire \u_cpu._0026_ ;
 wire \u_cpu._0027_ ;
 wire \u_cpu._0028_ ;
 wire \u_cpu._0029_ ;
 wire \u_cpu._0030_ ;
 wire \u_cpu._0031_ ;
 wire \u_cpu._0032_ ;
 wire \u_cpu._0033_ ;
 wire \u_cpu._0034_ ;
 wire \u_cpu._0035_ ;
 wire \u_cpu._0036_ ;
 wire \u_cpu._0037_ ;
 wire \u_cpu._0038_ ;
 wire \u_cpu._0039_ ;
 wire \u_cpu._0040_ ;
 wire \u_cpu._0041_ ;
 wire \u_cpu._0042_ ;
 wire \u_cpu._0043_ ;
 wire \u_cpu._0044_ ;
 wire \u_cpu._0045_ ;
 wire \u_cpu._0046_ ;
 wire \u_cpu._0047_ ;
 wire \u_cpu._0048_ ;
 wire \u_cpu._0049_ ;
 wire \u_cpu._0050_ ;
 wire \u_cpu._0051_ ;
 wire \u_cpu._0052_ ;
 wire \u_cpu._0053_ ;
 wire \u_cpu._0054_ ;
 wire \u_cpu._0055_ ;
 wire \u_cpu._0056_ ;
 wire \u_cpu._0057_ ;
 wire \u_cpu._0058_ ;
 wire \u_cpu._0059_ ;
 wire \u_cpu._0060_ ;
 wire \u_cpu._0061_ ;
 wire \u_cpu._0062_ ;
 wire \u_cpu._0063_ ;
 wire \u_cpu._0064_ ;
 wire \u_cpu._0065_ ;
 wire \u_cpu._0066_ ;
 wire \u_cpu._0067_ ;
 wire \u_cpu._0068_ ;
 wire \u_cpu._0069_ ;
 wire \u_cpu._0070_ ;
 wire \u_cpu._0071_ ;
 wire \u_cpu._0072_ ;
 wire \u_cpu._0073_ ;
 wire \u_cpu._0074_ ;
 wire \u_cpu._0075_ ;
 wire \u_cpu._0076_ ;
 wire \u_cpu._0077_ ;
 wire \u_cpu._0078_ ;
 wire \u_cpu._0079_ ;
 wire \u_cpu._0080_ ;
 wire \u_cpu._0081_ ;
 wire \u_cpu._0082_ ;
 wire \u_cpu._0083_ ;
 wire \u_cpu._0084_ ;
 wire \u_cpu._0085_ ;
 wire \u_cpu._0086_ ;
 wire \u_cpu._0087_ ;
 wire \u_cpu._0088_ ;
 wire \u_cpu._0089_ ;
 wire \u_cpu._0090_ ;
 wire \u_cpu._0091_ ;
 wire \u_cpu._0092_ ;
 wire \u_cpu._0093_ ;
 wire \u_cpu._0094_ ;
 wire \u_cpu._0095_ ;
 wire \u_cpu._0096_ ;
 wire \u_cpu._0097_ ;
 wire \u_cpu._0098_ ;
 wire \u_cpu._0099_ ;
 wire \u_cpu._0100_ ;
 wire \u_cpu._0101_ ;
 wire \u_cpu._0102_ ;
 wire \u_cpu._0103_ ;
 wire \u_cpu._0104_ ;
 wire \u_cpu._0105_ ;
 wire \u_cpu._0106_ ;
 wire \u_cpu._0107_ ;
 wire \u_cpu._0108_ ;
 wire \u_cpu._0109_ ;
 wire \u_cpu._0110_ ;
 wire \u_cpu._0111_ ;
 wire \u_cpu._0112_ ;
 wire \u_cpu._0113_ ;
 wire \u_cpu._0114_ ;
 wire \u_cpu._0115_ ;
 wire \u_cpu._0116_ ;
 wire \u_cpu._0117_ ;
 wire \u_cpu._0118_ ;
 wire \u_cpu._0119_ ;
 wire \u_cpu._0120_ ;
 wire \u_cpu._0121_ ;
 wire \u_cpu._0122_ ;
 wire \u_cpu._0123_ ;
 wire \u_cpu._0124_ ;
 wire \u_cpu._0125_ ;
 wire \u_cpu._0126_ ;
 wire \u_cpu._0127_ ;
 wire \u_cpu._0128_ ;
 wire \u_cpu._0129_ ;
 wire \u_cpu._0130_ ;
 wire \u_cpu._0131_ ;
 wire \u_cpu._0132_ ;
 wire \u_cpu._0133_ ;
 wire \u_cpu._0134_ ;
 wire \u_cpu._0135_ ;
 wire \u_cpu._0136_ ;
 wire \u_cpu._0137_ ;
 wire \u_cpu._0138_ ;
 wire \u_cpu._0139_ ;
 wire \u_cpu._0140_ ;
 wire \u_cpu._0141_ ;
 wire \u_cpu._0142_ ;
 wire \u_cpu._0143_ ;
 wire \u_cpu._0144_ ;
 wire \u_cpu._0145_ ;
 wire \u_cpu._0146_ ;
 wire \u_cpu._0147_ ;
 wire \u_cpu._0148_ ;
 wire \u_cpu._0149_ ;
 wire \u_cpu._0150_ ;
 wire \u_cpu._0151_ ;
 wire \u_cpu._0152_ ;
 wire \u_cpu._0153_ ;
 wire \u_cpu._0154_ ;
 wire \u_cpu._0155_ ;
 wire \u_cpu._0156_ ;
 wire \u_cpu._0157_ ;
 wire \u_cpu._0158_ ;
 wire \u_cpu._0159_ ;
 wire \u_cpu._0160_ ;
 wire \u_cpu._0161_ ;
 wire \u_cpu._0162_ ;
 wire \u_cpu._0163_ ;
 wire \u_cpu._0164_ ;
 wire \u_cpu._0165_ ;
 wire \u_cpu._0166_ ;
 wire \u_cpu._0167_ ;
 wire \u_cpu._0168_ ;
 wire \u_cpu._0169_ ;
 wire \u_cpu._0170_ ;
 wire \u_cpu._0171_ ;
 wire \u_cpu._0172_ ;
 wire \u_cpu._0173_ ;
 wire \u_cpu._0174_ ;
 wire \u_cpu._0175_ ;
 wire \u_cpu._0176_ ;
 wire \u_cpu._0177_ ;
 wire \u_cpu._0178_ ;
 wire \u_cpu._0179_ ;
 wire \u_cpu._0180_ ;
 wire \u_cpu._0181_ ;
 wire \u_cpu._0182_ ;
 wire \u_cpu._0183_ ;
 wire \u_cpu._0184_ ;
 wire \u_cpu._0185_ ;
 wire \u_cpu._0186_ ;
 wire \u_cpu._0187_ ;
 wire \u_cpu._0188_ ;
 wire \u_cpu._0189_ ;
 wire \u_cpu._0190_ ;
 wire \u_cpu._0191_ ;
 wire \u_cpu._0192_ ;
 wire \u_cpu._0193_ ;
 wire \u_cpu._0194_ ;
 wire \u_cpu._0195_ ;
 wire \u_cpu._0196_ ;
 wire \u_cpu._0197_ ;
 wire \u_cpu._0198_ ;
 wire \u_cpu._0199_ ;
 wire \u_cpu._0200_ ;
 wire \u_cpu._0201_ ;
 wire \u_cpu._0202_ ;
 wire \u_cpu._0203_ ;
 wire \u_cpu._0204_ ;
 wire \u_cpu._0205_ ;
 wire \u_cpu._0206_ ;
 wire \u_cpu._0207_ ;
 wire \u_cpu._0208_ ;
 wire \u_cpu._0209_ ;
 wire \u_cpu._0210_ ;
 wire \u_cpu._0211_ ;
 wire \u_cpu._0212_ ;
 wire \u_cpu._0213_ ;
 wire \u_cpu._0214_ ;
 wire \u_cpu._0215_ ;
 wire \u_cpu._0216_ ;
 wire \u_cpu._0217_ ;
 wire \u_cpu._0218_ ;
 wire \u_cpu._0219_ ;
 wire \u_cpu._0220_ ;
 wire \u_cpu._0221_ ;
 wire \u_cpu._0222_ ;
 wire \u_cpu._0223_ ;
 wire \u_cpu._0224_ ;
 wire \u_cpu._0225_ ;
 wire \u_cpu._0226_ ;
 wire \u_cpu._0227_ ;
 wire \u_cpu._0228_ ;
 wire \u_cpu._0229_ ;
 wire \u_cpu._0230_ ;
 wire \u_cpu._0231_ ;
 wire \u_cpu._0232_ ;
 wire \u_cpu._0233_ ;
 wire \u_cpu._0234_ ;
 wire \u_cpu._0235_ ;
 wire \u_cpu._0236_ ;
 wire \u_cpu._0237_ ;
 wire \u_cpu._0238_ ;
 wire \u_cpu._0239_ ;
 wire \u_cpu._0240_ ;
 wire \u_cpu._0241_ ;
 wire \u_cpu._0242_ ;
 wire \u_cpu._0243_ ;
 wire \u_cpu._0244_ ;
 wire \u_cpu._0245_ ;
 wire \u_cpu._0246_ ;
 wire \u_cpu._0247_ ;
 wire \u_cpu._0248_ ;
 wire \u_cpu._0249_ ;
 wire \u_cpu._0250_ ;
 wire \u_cpu._0251_ ;
 wire \u_cpu._0252_ ;
 wire \u_cpu._0253_ ;
 wire \u_cpu._0254_ ;
 wire \u_cpu._0255_ ;
 wire \u_cpu._0256_ ;
 wire \u_cpu._0257_ ;
 wire \u_cpu._0258_ ;
 wire \u_cpu._0259_ ;
 wire \u_cpu._0260_ ;
 wire \u_cpu._0261_ ;
 wire \u_cpu._0262_ ;
 wire \u_cpu._0263_ ;
 wire \u_cpu._0264_ ;
 wire \u_cpu._0265_ ;
 wire \u_cpu._0266_ ;
 wire \u_cpu._0267_ ;
 wire \u_cpu._0268_ ;
 wire \u_cpu._0269_ ;
 wire \u_cpu._0270_ ;
 wire \u_cpu._0271_ ;
 wire \u_cpu._0272_ ;
 wire \u_cpu._0273_ ;
 wire \u_cpu._0274_ ;
 wire \u_cpu._0275_ ;
 wire \u_cpu._0276_ ;
 wire \u_cpu._0277_ ;
 wire \u_cpu._0278_ ;
 wire \u_cpu._0279_ ;
 wire \u_cpu._0280_ ;
 wire \u_cpu._0281_ ;
 wire \u_cpu._0282_ ;
 wire \u_cpu._0283_ ;
 wire \u_cpu._0284_ ;
 wire \u_cpu._0285_ ;
 wire \u_cpu._0286_ ;
 wire \u_cpu._0287_ ;
 wire \u_cpu._0288_ ;
 wire \u_cpu._0289_ ;
 wire \u_cpu._0290_ ;
 wire \u_cpu._0291_ ;
 wire \u_cpu._0292_ ;
 wire \u_cpu._0293_ ;
 wire \u_cpu._0294_ ;
 wire \u_cpu._0295_ ;
 wire \u_cpu._0296_ ;
 wire \u_cpu._0297_ ;
 wire \u_cpu._0298_ ;
 wire \u_cpu._0299_ ;
 wire \u_cpu._0300_ ;
 wire \u_cpu._0301_ ;
 wire \u_cpu._0302_ ;
 wire \u_cpu._0303_ ;
 wire \u_cpu._0304_ ;
 wire \u_cpu._0305_ ;
 wire \u_cpu._0306_ ;
 wire \u_cpu._0307_ ;
 wire \u_cpu._0308_ ;
 wire \u_cpu._0309_ ;
 wire \u_cpu._0310_ ;
 wire \u_cpu._0311_ ;
 wire \u_cpu._0312_ ;
 wire \u_cpu._0313_ ;
 wire \u_cpu._0314_ ;
 wire \u_cpu._0315_ ;
 wire \u_cpu._0316_ ;
 wire \u_cpu._0317_ ;
 wire \u_cpu._0318_ ;
 wire \u_cpu._0319_ ;
 wire \u_cpu._0320_ ;
 wire \u_cpu._0321_ ;
 wire \u_cpu._0322_ ;
 wire \u_cpu._0323_ ;
 wire \u_cpu._0324_ ;
 wire \u_cpu._0325_ ;
 wire \u_cpu._0326_ ;
 wire \u_cpu._0327_ ;
 wire \u_cpu._0328_ ;
 wire \u_cpu._0329_ ;
 wire \u_cpu._0330_ ;
 wire \u_cpu._0331_ ;
 wire \u_cpu._0332_ ;
 wire \u_cpu._0333_ ;
 wire \u_cpu._0334_ ;
 wire \u_cpu._0335_ ;
 wire \u_cpu._0336_ ;
 wire \u_cpu._0337_ ;
 wire \u_cpu._0338_ ;
 wire \u_cpu._0339_ ;
 wire \u_cpu._0340_ ;
 wire \u_cpu._0341_ ;
 wire \u_cpu._0342_ ;
 wire \u_cpu._0343_ ;
 wire \u_cpu._0344_ ;
 wire \u_cpu._0345_ ;
 wire \u_cpu._0346_ ;
 wire \u_cpu._0347_ ;
 wire \u_cpu._0348_ ;
 wire \u_cpu._0349_ ;
 wire \u_cpu._0350_ ;
 wire \u_cpu._0351_ ;
 wire \u_cpu._0352_ ;
 wire \u_cpu._0353_ ;
 wire \u_cpu._0354_ ;
 wire \u_cpu._0355_ ;
 wire \u_cpu._0356_ ;
 wire \u_cpu._0357_ ;
 wire \u_cpu._0358_ ;
 wire \u_cpu._0359_ ;
 wire \u_cpu._0360_ ;
 wire \u_cpu._0361_ ;
 wire \u_cpu._0362_ ;
 wire \u_cpu._0363_ ;
 wire \u_cpu._0364_ ;
 wire \u_cpu._0365_ ;
 wire \u_cpu._0366_ ;
 wire \u_cpu._0367_ ;
 wire \u_cpu._0368_ ;
 wire \u_cpu._0369_ ;
 wire \u_cpu._0370_ ;
 wire \u_cpu._0371_ ;
 wire \u_cpu._0372_ ;
 wire \u_cpu._0373_ ;
 wire \u_cpu._0374_ ;
 wire \u_cpu._0375_ ;
 wire \u_cpu._0376_ ;
 wire \u_cpu._0377_ ;
 wire \u_cpu._0378_ ;
 wire \u_cpu._0379_ ;
 wire \u_cpu._0380_ ;
 wire \u_cpu._0381_ ;
 wire \u_cpu._0382_ ;
 wire \u_cpu._0383_ ;
 wire \u_cpu._0384_ ;
 wire \u_cpu._0385_ ;
 wire \u_cpu._0386_ ;
 wire \u_cpu._0387_ ;
 wire \u_cpu._0388_ ;
 wire \u_cpu._0389_ ;
 wire \u_cpu._0390_ ;
 wire \u_cpu._0391_ ;
 wire \u_cpu._0392_ ;
 wire \u_cpu._0393_ ;
 wire \u_cpu._0394_ ;
 wire \u_cpu._0395_ ;
 wire \u_cpu._0396_ ;
 wire \u_cpu._0397_ ;
 wire \u_cpu._0398_ ;
 wire \u_cpu._0399_ ;
 wire \u_cpu._0400_ ;
 wire \u_cpu._0401_ ;
 wire \u_cpu._0402_ ;
 wire \u_cpu._0403_ ;
 wire \u_cpu._0404_ ;
 wire \u_cpu._0405_ ;
 wire \u_cpu._0406_ ;
 wire \u_cpu._0407_ ;
 wire \u_cpu._0408_ ;
 wire \u_cpu._0409_ ;
 wire \u_cpu._0410_ ;
 wire \u_cpu._0411_ ;
 wire \u_cpu._0412_ ;
 wire \u_cpu._0413_ ;
 wire \u_cpu._0414_ ;
 wire \u_cpu._0415_ ;
 wire \u_cpu._0416_ ;
 wire \u_cpu._0417_ ;
 wire \u_cpu._0418_ ;
 wire \u_cpu._0419_ ;
 wire \u_cpu._0420_ ;
 wire \u_cpu._0421_ ;
 wire \u_cpu._0422_ ;
 wire \u_cpu._0423_ ;
 wire \u_cpu._0424_ ;
 wire \u_cpu._0425_ ;
 wire \u_cpu._0426_ ;
 wire \u_cpu._0427_ ;
 wire \u_cpu._0428_ ;
 wire \u_cpu._0429_ ;
 wire \u_cpu._0430_ ;
 wire \u_cpu._0431_ ;
 wire \u_cpu._0432_ ;
 wire \u_cpu._0433_ ;
 wire \u_cpu._0434_ ;
 wire \u_cpu._0435_ ;
 wire \u_cpu._0436_ ;
 wire \u_cpu._0437_ ;
 wire \u_cpu._0438_ ;
 wire \u_cpu._0439_ ;
 wire \u_cpu._0440_ ;
 wire \u_cpu._0441_ ;
 wire \u_cpu._0442_ ;
 wire \u_cpu._0443_ ;
 wire \u_cpu._0444_ ;
 wire \u_cpu._0445_ ;
 wire \u_cpu._0446_ ;
 wire \u_cpu._0447_ ;
 wire \u_cpu._0448_ ;
 wire \u_cpu._0449_ ;
 wire \u_cpu._0450_ ;
 wire \u_cpu._0451_ ;
 wire \u_cpu._0452_ ;
 wire \u_cpu._0453_ ;
 wire \u_cpu._0454_ ;
 wire \u_cpu._0455_ ;
 wire \u_cpu._0456_ ;
 wire \u_cpu._0457_ ;
 wire \u_cpu._0458_ ;
 wire \u_cpu._0459_ ;
 wire \u_cpu._0460_ ;
 wire \u_cpu._0461_ ;
 wire \u_cpu._0462_ ;
 wire \u_cpu._0463_ ;
 wire \u_cpu._0464_ ;
 wire \u_cpu._0465_ ;
 wire \u_cpu._0466_ ;
 wire \u_cpu._0467_ ;
 wire \u_cpu._0468_ ;
 wire \u_cpu._0469_ ;
 wire \u_cpu._0470_ ;
 wire \u_cpu._0471_ ;
 wire \u_cpu._0472_ ;
 wire \u_cpu._0473_ ;
 wire \u_cpu._0474_ ;
 wire \u_cpu._0475_ ;
 wire \u_cpu._0476_ ;
 wire \u_cpu._0477_ ;
 wire \u_cpu._0478_ ;
 wire \u_cpu._0479_ ;
 wire \u_cpu._0480_ ;
 wire \u_cpu._0481_ ;
 wire \u_cpu._0482_ ;
 wire \u_cpu._0483_ ;
 wire \u_cpu._0484_ ;
 wire \u_cpu._0485_ ;
 wire \u_cpu._0486_ ;
 wire \u_cpu._0487_ ;
 wire \u_cpu._0488_ ;
 wire \u_cpu._0489_ ;
 wire \u_cpu._0490_ ;
 wire \u_cpu._0491_ ;
 wire \u_cpu._0492_ ;
 wire \u_cpu._0493_ ;
 wire \u_cpu._0494_ ;
 wire \u_cpu._0495_ ;
 wire \u_cpu._0496_ ;
 wire \u_cpu._0497_ ;
 wire \u_cpu._0498_ ;
 wire \u_cpu._0499_ ;
 wire \u_cpu._0500_ ;
 wire \u_cpu._0501_ ;
 wire \u_cpu._0502_ ;
 wire \u_cpu._0503_ ;
 wire \u_cpu._0504_ ;
 wire \u_cpu._0505_ ;
 wire \u_cpu._0506_ ;
 wire \u_cpu._0507_ ;
 wire \u_cpu._0508_ ;
 wire \u_cpu._0509_ ;
 wire \u_cpu._0510_ ;
 wire \u_cpu._0511_ ;
 wire \u_cpu._0512_ ;
 wire \u_cpu._0513_ ;
 wire \u_cpu._0514_ ;
 wire \u_cpu._0515_ ;
 wire \u_cpu._0516_ ;
 wire \u_cpu._0517_ ;
 wire \u_cpu._0518_ ;
 wire \u_cpu._0519_ ;
 wire \u_cpu._0520_ ;
 wire \u_cpu._0521_ ;
 wire \u_cpu._0522_ ;
 wire \u_cpu._0523_ ;
 wire \u_cpu._0524_ ;
 wire \u_cpu._0525_ ;
 wire \u_cpu._0526_ ;
 wire \u_cpu._0527_ ;
 wire \u_cpu._0528_ ;
 wire \u_cpu._0529_ ;
 wire \u_cpu._0530_ ;
 wire \u_cpu._0531_ ;
 wire \u_cpu._0532_ ;
 wire \u_cpu._0533_ ;
 wire \u_cpu._0534_ ;
 wire \u_cpu._0535_ ;
 wire \u_cpu._0536_ ;
 wire \u_cpu._0537_ ;
 wire \u_cpu._0538_ ;
 wire \u_cpu._0539_ ;
 wire \u_cpu._0540_ ;
 wire \u_cpu._0541_ ;
 wire \u_cpu._0542_ ;
 wire \u_cpu._0543_ ;
 wire \u_cpu._0544_ ;
 wire \u_cpu._0545_ ;
 wire \u_cpu._0546_ ;
 wire \u_cpu._0547_ ;
 wire \u_cpu._0548_ ;
 wire \u_cpu._0549_ ;
 wire \u_cpu._0550_ ;
 wire \u_cpu._0551_ ;
 wire \u_cpu._0552_ ;
 wire \u_cpu._0553_ ;
 wire \u_cpu._0554_ ;
 wire \u_cpu._0555_ ;
 wire \u_cpu._0556_ ;
 wire \u_cpu._0557_ ;
 wire \u_cpu._0558_ ;
 wire \u_cpu._0559_ ;
 wire \u_cpu._0560_ ;
 wire \u_cpu._0561_ ;
 wire \u_cpu._0562_ ;
 wire \u_cpu._0563_ ;
 wire \u_cpu._0564_ ;
 wire \u_cpu._0565_ ;
 wire \u_cpu._0566_ ;
 wire \u_cpu._0567_ ;
 wire \u_cpu._0568_ ;
 wire \u_cpu._0569_ ;
 wire \u_cpu._0570_ ;
 wire \u_cpu._0571_ ;
 wire \u_cpu._0572_ ;
 wire \u_cpu._0573_ ;
 wire \u_cpu._0574_ ;
 wire \u_cpu._0575_ ;
 wire \u_cpu._0576_ ;
 wire \u_cpu._0577_ ;
 wire \u_cpu._0578_ ;
 wire \u_cpu._0579_ ;
 wire \u_cpu._0580_ ;
 wire \u_cpu._0581_ ;
 wire \u_cpu._0582_ ;
 wire \u_cpu._0583_ ;
 wire \u_cpu._0584_ ;
 wire \u_cpu._0585_ ;
 wire \u_cpu._0586_ ;
 wire \u_cpu._0587_ ;
 wire \u_cpu._0588_ ;
 wire \u_cpu._0589_ ;
 wire \u_cpu._0590_ ;
 wire \u_cpu._0591_ ;
 wire \u_cpu._0592_ ;
 wire \u_cpu._0593_ ;
 wire \u_cpu._0594_ ;
 wire \u_cpu._0595_ ;
 wire \u_cpu._0596_ ;
 wire \u_cpu._0597_ ;
 wire \u_cpu._0598_ ;
 wire \u_cpu._0599_ ;
 wire \u_cpu._0600_ ;
 wire \u_cpu._0601_ ;
 wire \u_cpu._0602_ ;
 wire \u_cpu._0603_ ;
 wire \u_cpu._0604_ ;
 wire \u_cpu._0605_ ;
 wire \u_cpu._0606_ ;
 wire \u_cpu._0607_ ;
 wire \u_cpu._0608_ ;
 wire \u_cpu._0609_ ;
 wire \u_cpu._0610_ ;
 wire \u_cpu._0611_ ;
 wire \u_cpu._0612_ ;
 wire \u_cpu._0613_ ;
 wire \u_cpu._0614_ ;
 wire \u_cpu._0615_ ;
 wire \u_cpu._0616_ ;
 wire \u_cpu._0617_ ;
 wire \u_cpu._0618_ ;
 wire \u_cpu._0619_ ;
 wire \u_cpu._0620_ ;
 wire \u_cpu._0621_ ;
 wire \u_cpu._0622_ ;
 wire \u_cpu._0623_ ;
 wire \u_cpu._0624_ ;
 wire \u_cpu._0625_ ;
 wire \u_cpu._0626_ ;
 wire \u_cpu._0627_ ;
 wire \u_cpu._0628_ ;
 wire \u_cpu._0629_ ;
 wire \u_cpu._0630_ ;
 wire \u_cpu._0631_ ;
 wire \u_cpu._0632_ ;
 wire \u_cpu._0633_ ;
 wire \u_cpu._0634_ ;
 wire \u_cpu._0635_ ;
 wire \u_cpu._0636_ ;
 wire \u_cpu._0637_ ;
 wire \u_cpu._0638_ ;
 wire \u_cpu._0639_ ;
 wire \u_cpu._0640_ ;
 wire \u_cpu._0641_ ;
 wire \u_cpu._0642_ ;
 wire \u_cpu._0643_ ;
 wire \u_cpu._0644_ ;
 wire \u_cpu._0645_ ;
 wire \u_cpu._0646_ ;
 wire \u_cpu._0647_ ;
 wire \u_cpu._0648_ ;
 wire \u_cpu._0649_ ;
 wire \u_cpu._0650_ ;
 wire \u_cpu._0651_ ;
 wire \u_cpu._0652_ ;
 wire \u_cpu._0653_ ;
 wire \u_cpu._0654_ ;
 wire \u_cpu.counter[0] ;
 wire \u_cpu.counter[10] ;
 wire \u_cpu.counter[11] ;
 wire \u_cpu.counter[12] ;
 wire \u_cpu.counter[13] ;
 wire \u_cpu.counter[14] ;
 wire \u_cpu.counter[15] ;
 wire \u_cpu.counter[16] ;
 wire \u_cpu.counter[17] ;
 wire \u_cpu.counter[18] ;
 wire \u_cpu.counter[19] ;
 wire \u_cpu.counter[1] ;
 wire \u_cpu.counter[20] ;
 wire \u_cpu.counter[21] ;
 wire \u_cpu.counter[22] ;
 wire \u_cpu.counter[23] ;
 wire \u_cpu.counter[24] ;
 wire \u_cpu.counter[25] ;
 wire \u_cpu.counter[2] ;
 wire \u_cpu.counter[3] ;
 wire \u_cpu.counter[4] ;
 wire \u_cpu.counter[5] ;
 wire \u_cpu.counter[6] ;
 wire \u_cpu.counter[7] ;
 wire \u_cpu.counter[8] ;
 wire \u_cpu.counter[9] ;
 wire \u_cpu.led[0] ;
 wire \u_cpu.led[1] ;
 wire \u_cpu.led[2] ;
 wire \u_cpu.led[3] ;
 wire \u_cpu.led[4] ;
 wire \u_cpu.led[5] ;
 wire \u_cpu.led[6] ;
 wire \u_cpu.led[7] ;
 wire \u_cpu.led[8] ;
 wire \u_cpu.led[9] ;
 wire \u_cpu.rst_n ;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_64_wb_clk_i;
 wire clknet_leaf_65_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_70_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_72_wb_clk_i;
 wire clknet_leaf_73_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_75_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_78_wb_clk_i;
 wire clknet_leaf_79_wb_clk_i;
 wire clknet_leaf_80_wb_clk_i;
 wire clknet_leaf_81_wb_clk_i;
 wire clknet_leaf_82_wb_clk_i;
 wire clknet_leaf_83_wb_clk_i;
 wire clknet_leaf_84_wb_clk_i;
 wire clknet_leaf_85_wb_clk_i;
 wire clknet_leaf_86_wb_clk_i;
 wire clknet_leaf_87_wb_clk_i;
 wire clknet_leaf_88_wb_clk_i;
 wire clknet_leaf_89_wb_clk_i;
 wire clknet_leaf_90_wb_clk_i;
 wire clknet_leaf_91_wb_clk_i;
 wire clknet_leaf_92_wb_clk_i;
 wire clknet_leaf_93_wb_clk_i;
 wire clknet_leaf_94_wb_clk_i;
 wire clknet_leaf_95_wb_clk_i;
 wire clknet_leaf_96_wb_clk_i;
 wire clknet_leaf_97_wb_clk_i;
 wire clknet_leaf_98_wb_clk_i;
 wire clknet_leaf_99_wb_clk_i;
 wire clknet_leaf_100_wb_clk_i;
 wire clknet_leaf_101_wb_clk_i;
 wire clknet_leaf_102_wb_clk_i;
 wire clknet_leaf_103_wb_clk_i;
 wire clknet_leaf_104_wb_clk_i;
 wire clknet_leaf_105_wb_clk_i;
 wire clknet_leaf_106_wb_clk_i;
 wire clknet_leaf_107_wb_clk_i;
 wire clknet_leaf_108_wb_clk_i;
 wire clknet_leaf_109_wb_clk_i;
 wire clknet_leaf_110_wb_clk_i;
 wire clknet_leaf_111_wb_clk_i;
 wire clknet_leaf_112_wb_clk_i;
 wire clknet_leaf_113_wb_clk_i;
 wire clknet_leaf_114_wb_clk_i;
 wire clknet_leaf_115_wb_clk_i;
 wire clknet_leaf_116_wb_clk_i;
 wire clknet_leaf_117_wb_clk_i;
 wire clknet_leaf_118_wb_clk_i;
 wire clknet_leaf_119_wb_clk_i;
 wire clknet_leaf_120_wb_clk_i;
 wire clknet_leaf_121_wb_clk_i;
 wire clknet_leaf_122_wb_clk_i;
 wire clknet_leaf_123_wb_clk_i;
 wire clknet_leaf_124_wb_clk_i;
 wire clknet_leaf_125_wb_clk_i;
 wire clknet_leaf_126_wb_clk_i;
 wire clknet_leaf_127_wb_clk_i;
 wire clknet_leaf_128_wb_clk_i;
 wire clknet_leaf_129_wb_clk_i;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_4_0__leaf_wb_clk_i;
 wire clknet_4_1__leaf_wb_clk_i;
 wire clknet_4_2__leaf_wb_clk_i;
 wire clknet_4_3__leaf_wb_clk_i;
 wire clknet_4_4__leaf_wb_clk_i;
 wire clknet_4_5__leaf_wb_clk_i;
 wire clknet_4_6__leaf_wb_clk_i;
 wire clknet_4_7__leaf_wb_clk_i;
 wire clknet_4_8__leaf_wb_clk_i;
 wire clknet_4_9__leaf_wb_clk_i;
 wire clknet_4_10__leaf_wb_clk_i;
 wire clknet_4_11__leaf_wb_clk_i;
 wire clknet_4_12__leaf_wb_clk_i;
 wire clknet_4_13__leaf_wb_clk_i;
 wire clknet_4_14__leaf_wb_clk_i;
 wire clknet_4_15__leaf_wb_clk_i;

 sky130_fd_sc_hd__inv_2 _48696_ (.A(wb_rst_i),
    .Y(_08226_));
 sky130_fd_sc_hd__buf_1 _48697_ (.A(_08226_),
    .X(\u_cpu.rst_n ));
 sky130_fd_sc_hd__conb_1 _71895_ (.LO(io_oeb[0]));
 sky130_fd_sc_hd__conb_1 _71896_ (.LO(io_oeb[1]));
 sky130_fd_sc_hd__conb_1 _71897_ (.LO(io_oeb[2]));
 sky130_fd_sc_hd__conb_1 _71898_ (.LO(io_oeb[3]));
 sky130_fd_sc_hd__conb_1 _71899_ (.LO(io_oeb[4]));
 sky130_fd_sc_hd__conb_1 _71900_ (.LO(io_oeb[5]));
 sky130_fd_sc_hd__conb_1 _71901_ (.LO(io_oeb[6]));
 sky130_fd_sc_hd__conb_1 _71902_ (.LO(io_oeb[7]));
 sky130_fd_sc_hd__conb_1 _71903_ (.LO(io_oeb[8]));
 sky130_fd_sc_hd__conb_1 _71904_ (.LO(io_oeb[9]));
 sky130_fd_sc_hd__conb_1 _71905_ (.LO(io_oeb[10]));
 sky130_fd_sc_hd__conb_1 _71906_ (.LO(io_oeb[11]));
 sky130_fd_sc_hd__conb_1 _71907_ (.LO(io_oeb[12]));
 sky130_fd_sc_hd__conb_1 _71908_ (.LO(io_oeb[13]));
 sky130_fd_sc_hd__conb_1 _71909_ (.LO(io_oeb[14]));
 sky130_fd_sc_hd__conb_1 _71910_ (.LO(io_oeb[15]));
 sky130_fd_sc_hd__conb_1 _71911_ (.LO(io_oeb[16]));
 sky130_fd_sc_hd__conb_1 _71912_ (.LO(io_oeb[17]));
 sky130_fd_sc_hd__conb_1 _71913_ (.LO(io_oeb[18]));
 sky130_fd_sc_hd__conb_1 _71914_ (.LO(io_oeb[19]));
 sky130_fd_sc_hd__conb_1 _71915_ (.LO(io_oeb[20]));
 sky130_fd_sc_hd__conb_1 _71916_ (.LO(io_oeb[21]));
 sky130_fd_sc_hd__conb_1 _71917_ (.LO(io_oeb[22]));
 sky130_fd_sc_hd__conb_1 _71918_ (.LO(io_oeb[23]));
 sky130_fd_sc_hd__conb_1 _71919_ (.LO(io_oeb[24]));
 sky130_fd_sc_hd__conb_1 _71920_ (.LO(io_oeb[25]));
 sky130_fd_sc_hd__conb_1 _71921_ (.LO(io_oeb[26]));
 sky130_fd_sc_hd__conb_1 _71922_ (.LO(io_oeb[27]));
 sky130_fd_sc_hd__conb_1 _71923_ (.LO(io_oeb[28]));
 sky130_fd_sc_hd__conb_1 _71924_ (.LO(io_oeb[29]));
 sky130_fd_sc_hd__conb_1 _71925_ (.LO(io_oeb[30]));
 sky130_fd_sc_hd__conb_1 _71926_ (.LO(io_oeb[31]));
 sky130_fd_sc_hd__conb_1 _71927_ (.LO(io_oeb[32]));
 sky130_fd_sc_hd__conb_1 _71928_ (.LO(io_oeb[33]));
 sky130_fd_sc_hd__conb_1 _71929_ (.LO(io_oeb[34]));
 sky130_fd_sc_hd__conb_1 _71930_ (.LO(io_oeb[35]));
 sky130_fd_sc_hd__conb_1 _71931_ (.LO(io_oeb[36]));
 sky130_fd_sc_hd__conb_1 _71932_ (.LO(io_oeb[37]));
 sky130_fd_sc_hd__conb_1 _71956_ (.LO(_71933_));
 sky130_fd_sc_hd__conb_1 _71957_ (.LO(_71934_));
 sky130_fd_sc_hd__conb_1 _71958_ (.LO(_71935_));
 sky130_fd_sc_hd__conb_1 _71959_ (.LO(_71936_));
 sky130_fd_sc_hd__conb_1 _71960_ (.LO(_71937_));
 sky130_fd_sc_hd__conb_1 _71961_ (.LO(_71938_));
 sky130_fd_sc_hd__conb_1 _71962_ (.LO(_71939_));
 sky130_fd_sc_hd__conb_1 _71963_ (.LO(_71940_));
 sky130_fd_sc_hd__conb_1 _71964_ (.LO(_71941_));
 sky130_fd_sc_hd__conb_1 _71965_ (.LO(_71942_));
 sky130_fd_sc_hd__conb_1 _71966_ (.LO(_71943_));
 sky130_fd_sc_hd__conb_1 _71967_ (.LO(_71944_));
 sky130_fd_sc_hd__conb_1 _71968_ (.LO(_71945_));
 sky130_fd_sc_hd__conb_1 _71969_ (.LO(_71946_));
 sky130_fd_sc_hd__conb_1 _71970_ (.LO(_71947_));
 sky130_fd_sc_hd__conb_1 _71971_ (.LO(_71948_));
 sky130_fd_sc_hd__conb_1 _71972_ (.LO(_71949_));
 sky130_fd_sc_hd__conb_1 _71973_ (.LO(_71950_));
 sky130_fd_sc_hd__conb_1 _71974_ (.LO(_71951_));
 sky130_fd_sc_hd__conb_1 _71975_ (.LO(_71952_));
 sky130_fd_sc_hd__conb_1 _71976_ (.LO(_71953_));
 sky130_fd_sc_hd__conb_1 _71977_ (.LO(_71954_));
 sky130_fd_sc_hd__conb_1 _71978_ (.LO(_71955_));
 sky130_fd_sc_hd__buf_2 _71979_ (.A(\u_cpu.led[0] ),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_2 _71980_ (.A(\u_cpu.led[1] ),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_2 _71981_ (.A(\u_cpu.led[2] ),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_2 _71982_ (.A(\u_cpu.led[3] ),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_2 _71983_ (.A(\u_cpu.led[4] ),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_2 _71984_ (.A(\u_cpu.led[5] ),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_2 _71985_ (.A(\u_cpu.led[6] ),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_2 _71986_ (.A(\u_cpu.led[7] ),
    .X(io_out[7]));
 sky130_fd_sc_hd__buf_2 _71987_ (.A(\u_cpu.led[8] ),
    .X(io_out[8]));
 sky130_fd_sc_hd__buf_2 _71988_ (.A(\u_cpu.led[9] ),
    .X(io_out[9]));
 sky130_fd_sc_hd__buf_2 _71989_ (.A(\u_cpu.M_AXI_WDATA[0] ),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_2 _71990_ (.A(\u_cpu.M_AXI_WDATA[1] ),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_2 _71991_ (.A(\u_cpu.M_AXI_WDATA[2] ),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_2 _71992_ (.A(\u_cpu.M_AXI_WDATA[3] ),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_2 _71993_ (.A(\u_cpu.M_AXI_WDATA[4] ),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_2 _71994_ (.A(\u_cpu.M_AXI_WDATA[5] ),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_2 _71995_ (.A(\u_cpu.M_AXI_WDATA[6] ),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_2 _71996_ (.A(\u_cpu.M_AXI_WDATA[7] ),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_2 _71997_ (.A(\u_cpu.M_AXI_WDATA[8] ),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_2 _71998_ (.A(\u_cpu.M_AXI_WDATA[9] ),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_2 _71999_ (.A(\u_cpu.M_AXI_WDATA[10] ),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_2 _72000_ (.A(\u_cpu.M_AXI_WDATA[11] ),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_2 _72001_ (.A(\u_cpu.M_AXI_AWADDR[0] ),
    .X(io_out[22]));
 sky130_fd_sc_hd__buf_2 _72002_ (.A(\u_cpu.M_AXI_AWADDR[1] ),
    .X(io_out[23]));
 sky130_fd_sc_hd__buf_2 _72003_ (.A(\u_cpu.M_AXI_AWADDR[2] ),
    .X(io_out[24]));
 sky130_fd_sc_hd__buf_2 _72004_ (.A(\u_cpu.M_AXI_AWADDR[3] ),
    .X(io_out[25]));
 sky130_fd_sc_hd__buf_2 _72005_ (.A(\u_cpu.M_AXI_AWADDR[4] ),
    .X(io_out[26]));
 sky130_fd_sc_hd__buf_2 _72006_ (.A(\u_cpu.M_AXI_AWADDR[5] ),
    .X(io_out[27]));
 sky130_fd_sc_hd__buf_2 _72007_ (.A(\u_cpu.M_AXI_AWADDR[6] ),
    .X(io_out[28]));
 sky130_fd_sc_hd__buf_2 _72008_ (.A(\u_cpu.M_AXI_AWADDR[7] ),
    .X(io_out[29]));
 sky130_fd_sc_hd__buf_2 _72009_ (.A(\u_cpu.M_AXI_AWADDR[8] ),
    .X(io_out[30]));
 sky130_fd_sc_hd__buf_2 _72010_ (.A(\u_cpu.M_AXI_AWADDR[9] ),
    .X(io_out[31]));
 sky130_fd_sc_hd__buf_2 _72011_ (.A(\u_cpu.M_AXI_AWADDR[10] ),
    .X(io_out[32]));
 sky130_fd_sc_hd__buf_2 _72012_ (.A(\u_cpu.M_AXI_AWADDR[11] ),
    .X(io_out[33]));
 sky130_fd_sc_hd__buf_2 _72013_ (.A(\u_cpu.M_AXI_AWADDR[12] ),
    .X(io_out[34]));
 sky130_fd_sc_hd__buf_2 _72014_ (.A(\u_cpu.M_AXI_AWADDR[13] ),
    .X(io_out[35]));
 sky130_fd_sc_hd__buf_2 _72015_ (.A(\u_cpu.M_AXI_AWADDR[14] ),
    .X(io_out[36]));
 sky130_fd_sc_hd__buf_2 _72016_ (.A(\u_cpu.M_AXI_AWADDR[15] ),
    .X(io_out[37]));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1351_  (.A(\u_cpu.ALU.SrcA[27] ),
    .X(\u_cpu.ALU._0338_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1352_  (.A(\u_cpu.ALU._0338_ ),
    .B(\u_cpu.ALU.SrcB[27] ),
    .Y(\u_cpu.ALU._0348_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1353_  (.A(\u_cpu.ALU.SrcA[27] ),
    .Y(\u_cpu.ALU._0359_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1354_  (.A(\u_cpu.ALU.SrcB[27] ),
    .Y(\u_cpu.ALU._0370_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1355_  (.A(\u_cpu.ALU._0359_ ),
    .B(\u_cpu.ALU._0370_ ),
    .Y(\u_cpu.ALU._0380_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1356_  (.A(\u_cpu.ALU._0348_ ),
    .B(\u_cpu.ALU._0380_ ),
    .Y(\u_cpu.ALU._0391_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1357_  (.A(\u_cpu.ALU.SrcA[26] ),
    .B(\u_cpu.ALU.SrcB[26] ),
    .Y(\u_cpu.ALU._0401_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1358_  (.A(\u_cpu.ALU.SrcA[26] ),
    .B(\u_cpu.ALU.SrcB[26] ),
    .X(\u_cpu.ALU._0412_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1359_  (.A(\u_cpu.ALU._0401_ ),
    .B(\u_cpu.ALU._0412_ ),
    .Y(\u_cpu.ALU._0423_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1360_  (.A(\u_cpu.ALU.SrcA[24] ),
    .X(\u_cpu.ALU._0433_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1361_  (.A(\u_cpu.ALU.SrcB[24] ),
    .X(\u_cpu.ALU._0444_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU._1362_  (.A(\u_cpu.ALU._0433_ ),
    .B(\u_cpu.ALU._0444_ ),
    .X(\u_cpu.ALU._0454_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1363_  (.A(\u_cpu.ALU._0433_ ),
    .B(\u_cpu.ALU._0444_ ),
    .Y(\u_cpu.ALU._0465_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1364_  (.A(\u_cpu.ALU.SrcA[25] ),
    .X(\u_cpu.ALU._0475_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1365_  (.A(\u_cpu.ALU._0475_ ),
    .B(\u_cpu.ALU.SrcB[25] ),
    .Y(\u_cpu.ALU._0486_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1366_  (.A(\u_cpu.ALU.SrcA[25] ),
    .B(\u_cpu.ALU.SrcB[25] ),
    .X(\u_cpu.ALU._0496_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1367_  (.A(\u_cpu.ALU._0486_ ),
    .B(\u_cpu.ALU._0496_ ),
    .Y(\u_cpu.ALU._0507_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1368_  (.A1(\u_cpu.ALU._0454_ ),
    .A2(\u_cpu.ALU._0465_ ),
    .B1(\u_cpu.ALU._0507_ ),
    .Y(\u_cpu.ALU._0515_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1369_  (.A(\u_cpu.ALU.SrcA[30] ),
    .X(\u_cpu.ALU._0516_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1370_  (.A(\u_cpu.ALU._0516_ ),
    .B(\u_cpu.ALU.SrcB[30] ),
    .Y(\u_cpu.ALU._0517_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1371_  (.A(\u_cpu.ALU.SrcA[30] ),
    .B(\u_cpu.ALU.SrcB[30] ),
    .X(\u_cpu.ALU._0518_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU._1372_  (.A(\u_cpu.ALU.SrcA[28] ),
    .B(\u_cpu.ALU.SrcB[28] ),
    .X(\u_cpu.ALU._0519_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1373_  (.A(\u_cpu.ALU.SrcA[28] ),
    .B(\u_cpu.ALU.SrcB[28] ),
    .Y(\u_cpu.ALU._0520_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1374_  (.A(\u_cpu.ALU.SrcA[29] ),
    .B(\u_cpu.ALU.SrcB[29] ),
    .Y(\u_cpu.ALU._0521_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1375_  (.A(\u_cpu.ALU.SrcA[29] ),
    .B(\u_cpu.ALU.SrcB[29] ),
    .X(\u_cpu.ALU._0522_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU._1376_  (.A1_N(\u_cpu.ALU._0519_ ),
    .A2_N(\u_cpu.ALU._0520_ ),
    .B1(\u_cpu.ALU._0521_ ),
    .B2(\u_cpu.ALU._0522_ ),
    .X(\u_cpu.ALU._0523_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1377_  (.A(\u_cpu.ALU.SrcA[31] ),
    .B(\u_cpu.ALU.SrcB[31] ),
    .X(\u_cpu.ALU._0524_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1378_  (.A(\u_cpu.ALU.SrcA[31] ),
    .B(\u_cpu.ALU.SrcB[31] ),
    .Y(\u_cpu.ALU._0525_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1379_  (.A(\u_cpu.ALU._0524_ ),
    .B(\u_cpu.ALU._0525_ ),
    .Y(\u_cpu.ALU._0526_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1380_  (.A(\u_cpu.ALU._0526_ ),
    .Y(\u_cpu.ALU._0527_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._1381_  (.A1(\u_cpu.ALU._0517_ ),
    .A2(\u_cpu.ALU._0518_ ),
    .B1(\u_cpu.ALU._0523_ ),
    .C1(\u_cpu.ALU._0527_ ),
    .X(\u_cpu.ALU._0528_ ));
 sky130_fd_sc_hd__or4bb_2 \u_cpu.ALU._1382_  (.A(\u_cpu.ALU._0391_ ),
    .B(\u_cpu.ALU._0423_ ),
    .C_N(\u_cpu.ALU._0515_ ),
    .D_N(\u_cpu.ALU._0528_ ),
    .X(\u_cpu.ALU._0529_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU._1383_  (.A(\u_cpu.ALU.SrcA[19] ),
    .B(\u_cpu.ALU.SrcB[19] ),
    .X(\u_cpu.ALU._0530_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1384_  (.A(\u_cpu.ALU.SrcA[19] ),
    .B(\u_cpu.ALU.SrcB[19] ),
    .Y(\u_cpu.ALU._0531_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1385_  (.A(\u_cpu.ALU._0530_ ),
    .B(\u_cpu.ALU._0531_ ),
    .X(\u_cpu.ALU._0532_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1386_  (.A(\u_cpu.ALU.SrcA[18] ),
    .X(\u_cpu.ALU._0533_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1387_  (.A(\u_cpu.ALU.SrcB[18] ),
    .X(\u_cpu.ALU._0534_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu.ALU._1388_  (.A(\u_cpu.ALU._0533_ ),
    .B(\u_cpu.ALU._0534_ ),
    .Y(\u_cpu.ALU._0535_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1389_  (.A(\u_cpu.ALU.SrcA[17] ),
    .X(\u_cpu.ALU._0536_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1390_  (.A(\u_cpu.ALU.SrcB[17] ),
    .X(\u_cpu.ALU._0537_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1391_  (.A(\u_cpu.ALU._0537_ ),
    .Y(\u_cpu.ALU._0538_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1392_  (.A(\u_cpu.ALU.SrcA[17] ),
    .B(\u_cpu.ALU._0537_ ),
    .Y(\u_cpu.ALU._0539_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1393_  (.A(\u_cpu.ALU.SrcA[17] ),
    .B(\u_cpu.ALU._0537_ ),
    .X(\u_cpu.ALU._0540_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.ALU._1394_  (.A_N(\u_cpu.ALU.SrcA[16] ),
    .B(\u_cpu.ALU.SrcB[16] ),
    .X(\u_cpu.ALU._0541_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1395_  (.A1(\u_cpu.ALU._0539_ ),
    .A2(\u_cpu.ALU._0540_ ),
    .B1(\u_cpu.ALU._0541_ ),
    .Y(\u_cpu.ALU._0542_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1396_  (.A1(\u_cpu.ALU._0536_ ),
    .A2(\u_cpu.ALU._0538_ ),
    .B1(\u_cpu.ALU._0542_ ),
    .Y(\u_cpu.ALU._0543_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1397_  (.A(\u_cpu.ALU.SrcA[18] ),
    .Y(\u_cpu.ALU._0544_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1398_  (.A(\u_cpu.ALU._0544_ ),
    .B(\u_cpu.ALU._0534_ ),
    .X(\u_cpu.ALU._0545_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1399_  (.A1(\u_cpu.ALU._0535_ ),
    .A2(\u_cpu.ALU._0543_ ),
    .B1(\u_cpu.ALU._0545_ ),
    .Y(\u_cpu.ALU._0546_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1400_  (.A(\u_cpu.ALU.SrcA[19] ),
    .X(\u_cpu.ALU._0547_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.ALU._1401_  (.A(\u_cpu.ALU._0547_ ),
    .B_N(\u_cpu.ALU.SrcB[19] ),
    .X(\u_cpu.ALU._0548_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1402_  (.A1(\u_cpu.ALU._0532_ ),
    .A2(\u_cpu.ALU._0546_ ),
    .B1(\u_cpu.ALU._0548_ ),
    .Y(\u_cpu.ALU._0549_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1403_  (.A(\u_cpu.ALU.SrcA[21] ),
    .B(\u_cpu.ALU.SrcB[21] ),
    .X(\u_cpu.ALU._0550_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1404_  (.A(\u_cpu.ALU.SrcA[21] ),
    .B(\u_cpu.ALU.SrcB[21] ),
    .Y(\u_cpu.ALU._0551_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1405_  (.A(\u_cpu.ALU.SrcA[23] ),
    .Y(\u_cpu.ALU._0552_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1406_  (.A(\u_cpu.ALU.SrcB[23] ),
    .Y(\u_cpu.ALU._0553_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1407_  (.A(\u_cpu.ALU._0552_ ),
    .B(\u_cpu.ALU._0553_ ),
    .Y(\u_cpu.ALU._0554_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1408_  (.A(\u_cpu.ALU.SrcA[23] ),
    .X(\u_cpu.ALU._0555_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1409_  (.A(\u_cpu.ALU._0555_ ),
    .B(\u_cpu.ALU.SrcB[23] ),
    .Y(\u_cpu.ALU._0556_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1410_  (.A(\u_cpu.ALU.SrcB[20] ),
    .X(\u_cpu.ALU._0557_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1411_  (.A(\u_cpu.ALU.SrcA[20] ),
    .B(\u_cpu.ALU._0557_ ),
    .Y(\u_cpu.ALU._0558_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU._1412_  (.A(\u_cpu.ALU.SrcA[20] ),
    .B(\u_cpu.ALU._0557_ ),
    .X(\u_cpu.ALU._0559_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1413_  (.A(\u_cpu.ALU.SrcA[22] ),
    .X(\u_cpu.ALU._0560_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1414_  (.A(\u_cpu.ALU._0560_ ),
    .B(\u_cpu.ALU.SrcB[22] ),
    .Y(\u_cpu.ALU._0561_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1415_  (.A(\u_cpu.ALU.SrcA[22] ),
    .Y(\u_cpu.ALU._0562_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1416_  (.A(\u_cpu.ALU.SrcB[22] ),
    .Y(\u_cpu.ALU._0563_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1417_  (.A(\u_cpu.ALU._0562_ ),
    .B(\u_cpu.ALU._0563_ ),
    .Y(\u_cpu.ALU._0564_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU._1418_  (.A1_N(\u_cpu.ALU._0558_ ),
    .A2_N(\u_cpu.ALU._0559_ ),
    .B1(\u_cpu.ALU._0561_ ),
    .B2(\u_cpu.ALU._0564_ ),
    .X(\u_cpu.ALU._0565_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU._1419_  (.A1(\u_cpu.ALU._0550_ ),
    .A2(\u_cpu.ALU._0551_ ),
    .B1(\u_cpu.ALU._0554_ ),
    .B2(\u_cpu.ALU._0556_ ),
    .C1(\u_cpu.ALU._0565_ ),
    .X(\u_cpu.ALU._0566_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1420_  (.A(\u_cpu.ALU._0560_ ),
    .B(\u_cpu.ALU._0563_ ),
    .Y(\u_cpu.ALU._0567_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1421_  (.A(\u_cpu.ALU.SrcB[21] ),
    .Y(\u_cpu.ALU._0568_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU._1422_  (.A(\u_cpu.ALU.SrcA[21] ),
    .B(\u_cpu.ALU._0568_ ),
    .X(\u_cpu.ALU._0569_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1423_  (.A(\u_cpu.ALU.SrcA[20] ),
    .Y(\u_cpu.ALU._0570_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1424_  (.A1(\u_cpu.ALU._0550_ ),
    .A2(\u_cpu.ALU._0551_ ),
    .B1(\u_cpu.ALU._0570_ ),
    .C1(\u_cpu.ALU._0557_ ),
    .Y(\u_cpu.ALU._0571_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU._1425_  (.A1_N(\u_cpu.ALU._0561_ ),
    .A2_N(\u_cpu.ALU._0564_ ),
    .B1(\u_cpu.ALU._0569_ ),
    .B2(\u_cpu.ALU._0571_ ),
    .Y(\u_cpu.ALU._0572_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU._1426_  (.A1(\u_cpu.ALU._0554_ ),
    .A2(\u_cpu.ALU._0556_ ),
    .B1(\u_cpu.ALU._0567_ ),
    .B2(\u_cpu.ALU._0572_ ),
    .Y(\u_cpu.ALU._0573_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1427_  (.A1(\u_cpu.ALU._0555_ ),
    .A2(\u_cpu.ALU._0553_ ),
    .B1(\u_cpu.ALU._0573_ ),
    .Y(\u_cpu.ALU._0574_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1428_  (.A1(\u_cpu.ALU._0549_ ),
    .A2(\u_cpu.ALU._0566_ ),
    .B1(\u_cpu.ALU._0574_ ),
    .Y(\u_cpu.ALU._0575_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1429_  (.A(\u_cpu.ALU.SrcB[31] ),
    .Y(\u_cpu.ALU._0576_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1430_  (.A(\u_cpu.ALU.SrcA[31] ),
    .X(\u_cpu.ALU._0577_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.ALU._1431_  (.A(\u_cpu.ALU._0516_ ),
    .B_N(\u_cpu.ALU.SrcB[30] ),
    .X(\u_cpu.ALU._0578_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1432_  (.A(\u_cpu.ALU.SrcA[29] ),
    .X(\u_cpu.ALU._0579_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1433_  (.A(\u_cpu.ALU._0579_ ),
    .Y(\u_cpu.ALU._0580_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1434_  (.A(\u_cpu.ALU.SrcA[28] ),
    .X(\u_cpu.ALU._0581_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1435_  (.A(\u_cpu.ALU.SrcB[28] ),
    .X(\u_cpu.ALU._0582_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1436_  (.A1(\u_cpu.ALU._0521_ ),
    .A2(\u_cpu.ALU._0522_ ),
    .B1(\u_cpu.ALU._0582_ ),
    .Y(\u_cpu.ALU._0583_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU._1437_  (.A1_N(\u_cpu.ALU.SrcB[29] ),
    .A2_N(\u_cpu.ALU._0580_ ),
    .B1(\u_cpu.ALU._0581_ ),
    .B2(\u_cpu.ALU._0583_ ),
    .Y(\u_cpu.ALU._0584_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1438_  (.A1(\u_cpu.ALU._0517_ ),
    .A2(\u_cpu.ALU._0518_ ),
    .B1(\u_cpu.ALU._0584_ ),
    .Y(\u_cpu.ALU._0585_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.ALU._1439_  (.A1_N(\u_cpu.ALU._0524_ ),
    .A2_N(\u_cpu.ALU._0525_ ),
    .B1(\u_cpu.ALU._0578_ ),
    .B2(\u_cpu.ALU._0585_ ),
    .X(\u_cpu.ALU._0586_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1440_  (.A(\u_cpu.ALU._0338_ ),
    .B(\u_cpu.ALU._0370_ ),
    .Y(\u_cpu.ALU._0587_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1441_  (.A(\u_cpu.ALU.SrcA[26] ),
    .Y(\u_cpu.ALU._0588_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1442_  (.A(\u_cpu.ALU._0588_ ),
    .B(\u_cpu.ALU.SrcB[26] ),
    .Y(\u_cpu.ALU._0589_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.ALU._1443_  (.A_N(\u_cpu.ALU._0475_ ),
    .B(\u_cpu.ALU.SrcB[25] ),
    .X(\u_cpu.ALU._0590_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.ALU._1444_  (.A_N(\u_cpu.ALU.SrcA[24] ),
    .B(\u_cpu.ALU.SrcB[24] ),
    .X(\u_cpu.ALU._0591_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._1445_  (.A1(\u_cpu.ALU._0486_ ),
    .A2(\u_cpu.ALU._0496_ ),
    .B1(\u_cpu.ALU._0591_ ),
    .X(\u_cpu.ALU._0592_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU._1446_  (.A1(\u_cpu.ALU._0401_ ),
    .A2(\u_cpu.ALU._0412_ ),
    .B1(\u_cpu.ALU._0590_ ),
    .B2(\u_cpu.ALU._0592_ ),
    .Y(\u_cpu.ALU._0593_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU._1447_  (.A1_N(\u_cpu.ALU._0348_ ),
    .A2_N(\u_cpu.ALU._0380_ ),
    .B1(\u_cpu.ALU._0589_ ),
    .B2(\u_cpu.ALU._0593_ ),
    .Y(\u_cpu.ALU._0594_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1448_  (.A1(\u_cpu.ALU._0587_ ),
    .A2(\u_cpu.ALU._0594_ ),
    .B1(\u_cpu.ALU._0528_ ),
    .Y(\u_cpu.ALU._0595_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1449_  (.A1(\u_cpu.ALU._0576_ ),
    .A2(\u_cpu.ALU._0577_ ),
    .B1(\u_cpu.ALU._0586_ ),
    .C1(\u_cpu.ALU._0595_ ),
    .Y(\u_cpu.ALU._0596_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU._1450_  (.A1(\u_cpu.ALU._0529_ ),
    .A2(\u_cpu.ALU._0575_ ),
    .B1_N(\u_cpu.ALU._0596_ ),
    .Y(\u_cpu.ALU._0597_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1451_  (.A(\u_cpu.ALU.SrcA[7] ),
    .X(\u_cpu.ALU._0598_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1452_  (.A(\u_cpu.ALU.SrcB[7] ),
    .Y(\u_cpu.ALU._0599_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1453_  (.A(\u_cpu.ALU._0598_ ),
    .B(\u_cpu.ALU._0599_ ),
    .Y(\u_cpu.ALU._0600_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1454_  (.A(\u_cpu.ALU.SrcA[7] ),
    .B(\u_cpu.ALU.SrcB[7] ),
    .X(\u_cpu.ALU._0601_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU._1455_  (.A(\u_cpu.ALU.SrcA[7] ),
    .B(\u_cpu.ALU.SrcB[7] ),
    .X(\u_cpu.ALU._0602_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.ALU._1456_  (.A(\u_cpu.ALU._0601_ ),
    .B_N(\u_cpu.ALU._0602_ ),
    .X(\u_cpu.ALU._0603_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1457_  (.A(\u_cpu.ALU.SrcB[6] ),
    .Y(\u_cpu.ALU._0604_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1458_  (.A(\u_cpu.ALU.SrcA[6] ),
    .B(\u_cpu.ALU.SrcB[6] ),
    .Y(\u_cpu.ALU._0605_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1459_  (.A(\u_cpu.ALU.SrcA[6] ),
    .Y(\u_cpu.ALU._0606_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1460_  (.A(\u_cpu.ALU._0606_ ),
    .B(\u_cpu.ALU._0604_ ),
    .Y(\u_cpu.ALU._0607_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1461_  (.A(\u_cpu.ALU.SrcA[5] ),
    .X(\u_cpu.ALU._0608_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1462_  (.A(\u_cpu.ALU.SrcB[5] ),
    .X(\u_cpu.ALU._0609_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.ALU._1463_  (.A_N(\u_cpu.ALU._0608_ ),
    .B(\u_cpu.ALU._0609_ ),
    .X(\u_cpu.ALU._0610_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1464_  (.A(\u_cpu.ALU.SrcA[5] ),
    .B(\u_cpu.ALU._0609_ ),
    .Y(\u_cpu.ALU._0611_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1465_  (.A(\u_cpu.ALU.SrcA[5] ),
    .B(\u_cpu.ALU._0609_ ),
    .X(\u_cpu.ALU._0612_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1466_  (.A(\u_cpu.ALU.SrcB[4] ),
    .X(\u_cpu.ALU._0613_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.ALU._1467_  (.A_N(\u_cpu.ALU.SrcA[4] ),
    .B(\u_cpu.ALU._0613_ ),
    .X(\u_cpu.ALU._0614_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._1468_  (.A1(\u_cpu.ALU._0611_ ),
    .A2(\u_cpu.ALU._0612_ ),
    .B1(\u_cpu.ALU._0614_ ),
    .X(\u_cpu.ALU._0615_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU._1469_  (.A1(\u_cpu.ALU._0605_ ),
    .A2(\u_cpu.ALU._0607_ ),
    .B1(\u_cpu.ALU._0610_ ),
    .B2(\u_cpu.ALU._0615_ ),
    .Y(\u_cpu.ALU._0616_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1470_  (.A1(\u_cpu.ALU.SrcA[6] ),
    .A2(\u_cpu.ALU._0604_ ),
    .B1(\u_cpu.ALU._0616_ ),
    .Y(\u_cpu.ALU._0617_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1471_  (.A(\u_cpu.ALU.SrcA[4] ),
    .X(\u_cpu.ALU._0618_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1472_  (.A(\u_cpu.ALU._0613_ ),
    .B(\u_cpu.ALU._0618_ ),
    .Y(\u_cpu.ALU._0619_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1473_  (.A(\u_cpu.ALU._0613_ ),
    .B(\u_cpu.ALU.SrcA[4] ),
    .X(\u_cpu.ALU._0620_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU._1474_  (.A1(\u_cpu.ALU._0611_ ),
    .A2(\u_cpu.ALU._0612_ ),
    .B1(\u_cpu.ALU._0619_ ),
    .B2(\u_cpu.ALU._0620_ ),
    .X(\u_cpu.ALU._0621_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1475_  (.A1(\u_cpu.ALU._0605_ ),
    .A2(\u_cpu.ALU._0607_ ),
    .B1(\u_cpu.ALU._0621_ ),
    .C1(\u_cpu.ALU._0603_ ),
    .Y(\u_cpu.ALU._0622_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1476_  (.A(\u_cpu.ALU.SrcB[3] ),
    .X(\u_cpu.ALU._0623_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1477_  (.A(\u_cpu.ALU.SrcA[3] ),
    .X(\u_cpu.ALU._0624_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1478_  (.A(\u_cpu.ALU._0623_ ),
    .B(\u_cpu.ALU._0624_ ),
    .Y(\u_cpu.ALU._0625_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1479_  (.A(\u_cpu.ALU._0623_ ),
    .B(\u_cpu.ALU.SrcA[3] ),
    .X(\u_cpu.ALU._0626_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1480_  (.A(\u_cpu.ALU.SrcA[2] ),
    .X(\u_cpu.ALU._0627_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU._1481_  (.A(\u_cpu.ALU.SrcB[2] ),
    .B(\u_cpu.ALU._0627_ ),
    .X(\u_cpu.ALU._0628_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1482_  (.A(\u_cpu.ALU.SrcB[2] ),
    .X(\u_cpu.ALU._0629_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1483_  (.A(\u_cpu.ALU._0629_ ),
    .B(\u_cpu.ALU._0627_ ),
    .Y(\u_cpu.ALU._0630_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU._1484_  (.A1_N(\u_cpu.ALU._0625_ ),
    .A2_N(\u_cpu.ALU._0626_ ),
    .B1(\u_cpu.ALU._0628_ ),
    .B2(\u_cpu.ALU._0630_ ),
    .Y(\u_cpu.ALU._0631_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1485_  (.A(\u_cpu.ALU.SrcA[1] ),
    .X(\u_cpu.ALU._0632_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1486_  (.A(\u_cpu.ALU.SrcB[0] ),
    .X(\u_cpu.ALU._0633_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1487_  (.A(\u_cpu.ALU._0633_ ),
    .X(\u_cpu.ALU._0634_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1488_  (.A(\u_cpu.ALU._0634_ ),
    .X(\u_cpu.ALU._0635_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1489_  (.A(\u_cpu.ALU.SrcA[0] ),
    .Y(\u_cpu.ALU._0636_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1490_  (.A(\u_cpu.ALU.SrcB[1] ),
    .X(\u_cpu.ALU._0637_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1491_  (.A(\u_cpu.ALU._0637_ ),
    .X(\u_cpu.ALU._0638_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1492_  (.A1(\u_cpu.ALU._0635_ ),
    .A2(\u_cpu.ALU._0636_ ),
    .B1(\u_cpu.ALU._0638_ ),
    .Y(\u_cpu.ALU._0639_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1493_  (.A(\u_cpu.ALU.SrcB[0] ),
    .Y(\u_cpu.ALU._0640_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1494_  (.A(\u_cpu.ALU._0640_ ),
    .X(\u_cpu.ALU._0641_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1495_  (.A(\u_cpu.ALU._0637_ ),
    .Y(\u_cpu.ALU._0642_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1496_  (.A(\u_cpu.ALU._0642_ ),
    .X(\u_cpu.ALU._0643_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._1497_  (.A(\u_cpu.ALU._0641_ ),
    .B(\u_cpu.ALU._0643_ ),
    .C(\u_cpu.ALU.SrcA[0] ),
    .X(\u_cpu.ALU._0644_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1498_  (.A1(\u_cpu.ALU._0632_ ),
    .A2(\u_cpu.ALU._0639_ ),
    .B1(\u_cpu.ALU._0644_ ),
    .Y(\u_cpu.ALU._0645_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1499_  (.A(\u_cpu.ALU._0623_ ),
    .Y(\u_cpu.ALU._0646_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1500_  (.A(\u_cpu.ALU._0646_ ),
    .X(\u_cpu.ALU._0647_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1501_  (.A(\u_cpu.ALU.SrcA[2] ),
    .Y(\u_cpu.ALU._0648_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1502_  (.A1(\u_cpu.ALU._0625_ ),
    .A2(\u_cpu.ALU._0626_ ),
    .B1(\u_cpu.ALU._0629_ ),
    .C1(\u_cpu.ALU._0648_ ),
    .Y(\u_cpu.ALU._0649_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1503_  (.A1(\u_cpu.ALU._0647_ ),
    .A2(\u_cpu.ALU._0624_ ),
    .B1(\u_cpu.ALU._0649_ ),
    .Y(\u_cpu.ALU._0650_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1504_  (.A1(\u_cpu.ALU._0631_ ),
    .A2(\u_cpu.ALU._0645_ ),
    .B1(\u_cpu.ALU._0650_ ),
    .Y(\u_cpu.ALU._0651_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU._1505_  (.A1_N(\u_cpu.ALU._0603_ ),
    .A2_N(\u_cpu.ALU._0617_ ),
    .B1(\u_cpu.ALU._0622_ ),
    .B2(\u_cpu.ALU._0651_ ),
    .Y(\u_cpu.ALU._0652_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU._1506_  (.A(\u_cpu.ALU.SrcA[15] ),
    .B(\u_cpu.ALU.SrcB[15] ),
    .X(\u_cpu.ALU._0653_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1507_  (.A(\u_cpu.ALU.SrcB[14] ),
    .X(\u_cpu.ALU._0654_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1508_  (.A(\u_cpu.ALU.SrcA[14] ),
    .B(\u_cpu.ALU._0654_ ),
    .Y(\u_cpu.ALU._0655_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1509_  (.A(\u_cpu.ALU.SrcA[14] ),
    .B(\u_cpu.ALU._0654_ ),
    .Y(\u_cpu.ALU._0656_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.ALU._1510_  (.A_N(\u_cpu.ALU._0655_ ),
    .B(\u_cpu.ALU._0656_ ),
    .X(\u_cpu.ALU._0657_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1511_  (.A(\u_cpu.ALU.SrcB[13] ),
    .X(\u_cpu.ALU._0658_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu.ALU._1512_  (.A(\u_cpu.ALU.SrcA[13] ),
    .B(\u_cpu.ALU._0658_ ),
    .Y(\u_cpu.ALU._0659_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1513_  (.A(\u_cpu.ALU.SrcB[12] ),
    .X(\u_cpu.ALU._0660_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu.ALU._1514_  (.A(\u_cpu.ALU.SrcA[12] ),
    .B(\u_cpu.ALU._0660_ ),
    .Y(\u_cpu.ALU._0661_ ));
 sky130_fd_sc_hd__and4bb_2 \u_cpu.ALU._1515_  (.A_N(\u_cpu.ALU._0653_ ),
    .B_N(\u_cpu.ALU._0657_ ),
    .C(\u_cpu.ALU._0659_ ),
    .D(\u_cpu.ALU._0661_ ),
    .X(\u_cpu.ALU._0662_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1516_  (.A(\u_cpu.ALU.SrcA[8] ),
    .X(\u_cpu.ALU._0663_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1517_  (.A(\u_cpu.ALU.SrcB[8] ),
    .X(\u_cpu.ALU._0664_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu.ALU._1518_  (.A(\u_cpu.ALU._0663_ ),
    .B(\u_cpu.ALU._0664_ ),
    .Y(\u_cpu.ALU._0665_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1519_  (.A(\u_cpu.ALU.SrcA[10] ),
    .X(\u_cpu.ALU._0666_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1520_  (.A(\u_cpu.ALU.SrcB[10] ),
    .X(\u_cpu.ALU._0667_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu.ALU._1521_  (.A(\u_cpu.ALU._0666_ ),
    .B(\u_cpu.ALU._0667_ ),
    .Y(\u_cpu.ALU._0668_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1522_  (.A(\u_cpu.ALU.SrcA[9] ),
    .X(\u_cpu.ALU._0669_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1523_  (.A(\u_cpu.ALU._0669_ ),
    .B(\u_cpu.ALU.SrcB[9] ),
    .Y(\u_cpu.ALU._0670_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1524_  (.A(\u_cpu.ALU.SrcA[9] ),
    .B(\u_cpu.ALU.SrcB[9] ),
    .X(\u_cpu.ALU._0671_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU._1525_  (.A(\u_cpu.ALU.SrcA[11] ),
    .B(\u_cpu.ALU.SrcB[11] ),
    .X(\u_cpu.ALU._0672_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.ALU._1526_  (.A1(\u_cpu.ALU._0670_ ),
    .A2(\u_cpu.ALU._0671_ ),
    .B1_N(\u_cpu.ALU._0672_ ),
    .X(\u_cpu.ALU._0673_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU._1527_  (.A(\u_cpu.ALU._0662_ ),
    .B(\u_cpu.ALU._0665_ ),
    .C(\u_cpu.ALU._0668_ ),
    .D(\u_cpu.ALU._0673_ ),
    .X(\u_cpu.ALU._0674_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1528_  (.A1(\u_cpu.ALU._0600_ ),
    .A2(\u_cpu.ALU._0652_ ),
    .B1(\u_cpu.ALU._0674_ ),
    .Y(\u_cpu.ALU._0675_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1529_  (.A(\u_cpu.ALU.SrcA[12] ),
    .Y(\u_cpu.ALU._0676_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.ALU._1530_  (.A_N(\u_cpu.ALU.SrcA[13] ),
    .B(\u_cpu.ALU._0658_ ),
    .X(\u_cpu.ALU._0677_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU._1531_  (.A1(\u_cpu.ALU._0676_ ),
    .A2(\u_cpu.ALU._0659_ ),
    .A3(\u_cpu.ALU._0660_ ),
    .B1(\u_cpu.ALU._0677_ ),
    .Y(\u_cpu.ALU._0678_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1532_  (.A(\u_cpu.ALU.SrcA[14] ),
    .X(\u_cpu.ALU._0679_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1533_  (.A(\u_cpu.ALU._0679_ ),
    .Y(\u_cpu.ALU._0680_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1534_  (.A(\u_cpu.ALU._0680_ ),
    .B(\u_cpu.ALU._0654_ ),
    .Y(\u_cpu.ALU._0681_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._1535_  (.A1(\u_cpu.ALU._0657_ ),
    .A2(\u_cpu.ALU._0678_ ),
    .B1(\u_cpu.ALU._0681_ ),
    .X(\u_cpu.ALU._0682_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1536_  (.A(\u_cpu.ALU.SrcA[15] ),
    .Y(\u_cpu.ALU._0683_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1537_  (.A(\u_cpu.ALU._0683_ ),
    .B(\u_cpu.ALU.SrcB[15] ),
    .Y(\u_cpu.ALU._0684_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._1538_  (.A1(\u_cpu.ALU._0653_ ),
    .A2(\u_cpu.ALU._0682_ ),
    .B1(\u_cpu.ALU._0684_ ),
    .X(\u_cpu.ALU._0685_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1539_  (.A(\u_cpu.ALU.SrcA[11] ),
    .X(\u_cpu.ALU._0686_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1540_  (.A(\u_cpu.ALU.SrcB[11] ),
    .Y(\u_cpu.ALU._0687_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1541_  (.A(\u_cpu.ALU._0686_ ),
    .B(\u_cpu.ALU._0687_ ),
    .Y(\u_cpu.ALU._0688_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1542_  (.A(\u_cpu.ALU._0667_ ),
    .Y(\u_cpu.ALU._0689_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU._1543_  (.A(\u_cpu.ALU._0666_ ),
    .B(\u_cpu.ALU._0689_ ),
    .X(\u_cpu.ALU._0690_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1544_  (.A(\u_cpu.ALU.SrcB[9] ),
    .Y(\u_cpu.ALU._0691_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1545_  (.A(\u_cpu.ALU._0669_ ),
    .B(\u_cpu.ALU._0691_ ),
    .Y(\u_cpu.ALU._0692_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1546_  (.A(\u_cpu.ALU.SrcA[8] ),
    .Y(\u_cpu.ALU._0693_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._1547_  (.A1(\u_cpu.ALU._0670_ ),
    .A2(\u_cpu.ALU._0671_ ),
    .B1(\u_cpu.ALU._0693_ ),
    .C1(\u_cpu.ALU._0664_ ),
    .X(\u_cpu.ALU._0694_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1548_  (.A1(\u_cpu.ALU._0692_ ),
    .A2(\u_cpu.ALU._0694_ ),
    .B1(\u_cpu.ALU._0668_ ),
    .Y(\u_cpu.ALU._0695_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1549_  (.A1(\u_cpu.ALU._0690_ ),
    .A2(\u_cpu.ALU._0695_ ),
    .B1(\u_cpu.ALU._0672_ ),
    .Y(\u_cpu.ALU._0696_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1550_  (.A1(\u_cpu.ALU._0688_ ),
    .A2(\u_cpu.ALU._0696_ ),
    .B1(\u_cpu.ALU._0662_ ),
    .Y(\u_cpu.ALU._0697_ ));
 sky130_fd_sc_hd__and4bb_2 \u_cpu.ALU._1551_  (.A_N(\u_cpu.ALU._0391_ ),
    .B_N(\u_cpu.ALU._0423_ ),
    .C(\u_cpu.ALU._0515_ ),
    .D(\u_cpu.ALU._0528_ ),
    .X(\u_cpu.ALU._0698_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1552_  (.A(\u_cpu.ALU.SrcA[16] ),
    .X(\u_cpu.ALU._0699_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1553_  (.A(\u_cpu.ALU.SrcB[16] ),
    .X(\u_cpu.ALU._0700_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1554_  (.A(\u_cpu.ALU._0699_ ),
    .B(\u_cpu.ALU._0700_ ),
    .Y(\u_cpu.ALU._0701_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1555_  (.A(\u_cpu.ALU._0699_ ),
    .B(\u_cpu.ALU._0700_ ),
    .X(\u_cpu.ALU._0702_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU._1556_  (.A1_N(\u_cpu.ALU._0530_ ),
    .A2_N(\u_cpu.ALU._0531_ ),
    .B1(\u_cpu.ALU._0539_ ),
    .B2(\u_cpu.ALU._0540_ ),
    .X(\u_cpu.ALU._0703_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._1557_  (.A1(\u_cpu.ALU._0701_ ),
    .A2(\u_cpu.ALU._0702_ ),
    .B1(\u_cpu.ALU._0703_ ),
    .C1(\u_cpu.ALU._0535_ ),
    .D1(\u_cpu.ALU._0566_ ),
    .X(\u_cpu.ALU._0704_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1558_  (.A(\u_cpu.ALU._0698_ ),
    .B(\u_cpu.ALU._0704_ ),
    .Y(\u_cpu.ALU._0705_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU._1559_  (.A1(\u_cpu.ALU._0675_ ),
    .A2(\u_cpu.ALU._0685_ ),
    .A3(\u_cpu.ALU._0697_ ),
    .B1(\u_cpu.ALU._0705_ ),
    .Y(\u_cpu.ALU._0706_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.ALU._1560_  (.A(_71933_),
    .B_N(_71934_),
    .X(\u_cpu.ALU._0707_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1561_  (.A(\u_cpu.ALU._0707_ ),
    .X(\u_cpu.ALU._0708_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1562_  (.A(_71935_),
    .Y(\u_cpu.ALU._0709_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1563_  (.A(\u_cpu.ALU._0709_ ),
    .X(\u_cpu.ALU._0710_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1564_  (.A(\u_cpu.ALU._0710_ ),
    .X(\u_cpu.ALU._0711_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1565_  (.A(_71936_),
    .X(\u_cpu.ALU._0712_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1566_  (.A(\u_cpu.ALU._0711_ ),
    .B(\u_cpu.ALU._0712_ ),
    .Y(\u_cpu.ALU._0713_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._1567_  (.A1(\u_cpu.ALU._0708_ ),
    .A2(\u_cpu.ALU._0526_ ),
    .B1(\u_cpu.ALU._0713_ ),
    .X(\u_cpu.ALU._0714_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1568_  (.A1(\u_cpu.ALU._0597_ ),
    .A2(\u_cpu.ALU._0706_ ),
    .B1(\u_cpu.ALU._0714_ ),
    .Y(\u_cpu.ALU._0715_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._1569_  (.A1(\u_cpu.ALU._0549_ ),
    .A2(\u_cpu.ALU._0566_ ),
    .B1(\u_cpu.ALU._0574_ ),
    .X(\u_cpu.ALU._0716_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1570_  (.A1(\u_cpu.ALU._0716_ ),
    .A2(\u_cpu.ALU._0698_ ),
    .B1(\u_cpu.ALU._0596_ ),
    .Y(\u_cpu.ALU._0717_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._1571_  (.A1(\u_cpu.ALU._0675_ ),
    .A2(\u_cpu.ALU._0685_ ),
    .A3(\u_cpu.ALU._0697_ ),
    .B1(\u_cpu.ALU._0705_ ),
    .X(\u_cpu.ALU._0718_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1572_  (.A1(\u_cpu.ALU._0527_ ),
    .A2(\u_cpu.ALU._0708_ ),
    .B1(\u_cpu.ALU._0717_ ),
    .C1(\u_cpu.ALU._0718_ ),
    .Y(\u_cpu.ALU._0719_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1573_  (.A(\u_cpu.ALU.SrcB[0] ),
    .X(\u_cpu.ALU._0720_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1574_  (.A(\u_cpu.ALU._0720_ ),
    .X(\u_cpu.ALU._0721_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1575_  (.A(\u_cpu.ALU._0721_ ),
    .X(\u_cpu.ALU._0722_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1576_  (.A(\u_cpu.ALU._0722_ ),
    .X(\u_cpu.ALU._0723_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1577_  (.A(\u_cpu.ALU._0723_ ),
    .B(\u_cpu.ALU._0636_ ),
    .Y(\u_cpu.ALU._0724_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1578_  (.A(\u_cpu.ALU._0637_ ),
    .X(\u_cpu.ALU._0725_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1579_  (.A(\u_cpu.ALU._0725_ ),
    .X(\u_cpu.ALU._0726_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU._1580_  (.A(\u_cpu.ALU._0632_ ),
    .B(\u_cpu.ALU._0726_ ),
    .X(\u_cpu.ALU._0727_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1581_  (.A(\u_cpu.ALU._0637_ ),
    .X(\u_cpu.ALU._0728_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1582_  (.A(\u_cpu.ALU._0728_ ),
    .X(\u_cpu.ALU._0729_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1583_  (.A(\u_cpu.ALU._0632_ ),
    .B(\u_cpu.ALU._0729_ ),
    .Y(\u_cpu.ALU._0730_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1584_  (.A(\u_cpu.ALU._0727_ ),
    .B(\u_cpu.ALU._0730_ ),
    .Y(\u_cpu.ALU._0731_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1585_  (.A(\u_cpu.ALU._0636_ ),
    .B(\u_cpu.ALU._0721_ ),
    .Y(\u_cpu.ALU._0732_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.ALU._1586_  (.A_N(\u_cpu.ALU._0724_ ),
    .B(\u_cpu.ALU._0631_ ),
    .C(\u_cpu.ALU._0731_ ),
    .D(\u_cpu.ALU._0732_ ),
    .X(\u_cpu.ALU._0733_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU._1587_  (.A_N(\u_cpu.ALU._0622_ ),
    .B(\u_cpu.ALU._0674_ ),
    .C(\u_cpu.ALU._0733_ ),
    .Y(\u_cpu.ALU._0734_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1588_  (.A(_71937_),
    .X(\u_cpu.ALU._0735_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.ALU._1589_  (.A_N(\u_cpu.ALU._0735_ ),
    .B(_71938_),
    .X(\u_cpu.ALU._0736_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1590_  (.A(\u_cpu.ALU._0736_ ),
    .X(\u_cpu.ALU._0737_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1591_  (.A(\u_cpu.ALU._0737_ ),
    .X(\u_cpu.ALU._0738_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._1592_  (.A1(\u_cpu.ALU._0705_ ),
    .A2(\u_cpu.ALU._0734_ ),
    .B1(\u_cpu.ALU._0738_ ),
    .X(\u_cpu.ALU._0739_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._1593_  (.A(\u_cpu.ALU._0715_ ),
    .B(\u_cpu.ALU._0719_ ),
    .C(\u_cpu.ALU._0739_ ),
    .Y(\u_cpu.ALU._0740_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1594_  (.A(_71939_),
    .B(_71940_),
    .Y(\u_cpu.ALU._0741_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1595_  (.A(\u_cpu.ALU._0741_ ),
    .X(\u_cpu.ALU._0742_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._1596_  (.A(\u_cpu.ALU._0712_ ),
    .B(\u_cpu.ALU._0742_ ),
    .C(\u_cpu.ALU._0711_ ),
    .X(\u_cpu.ALU._0743_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1597_  (.A(\u_cpu.ALU._0743_ ),
    .X(\u_cpu.ALU._0744_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1598_  (.A(_71941_),
    .X(\u_cpu.ALU._0745_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1599_  (.A(\u_cpu.ALU._0745_ ),
    .X(\u_cpu.ALU._0746_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._1600_  (.A(\u_cpu.ALU._0712_ ),
    .B(\u_cpu.ALU._0746_ ),
    .C(\u_cpu.ALU._0742_ ),
    .X(\u_cpu.ALU._0747_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1601_  (.A(\u_cpu.ALU._0747_ ),
    .X(\u_cpu.ALU._0748_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1602_  (.A(\u_cpu.ALU._0748_ ),
    .X(\u_cpu.ALU._0749_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1603_  (.A(_71942_),
    .X(\u_cpu.ALU._0750_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1604_  (.A(\u_cpu.ALU._0735_ ),
    .X(\u_cpu.ALU._0751_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1605_  (.A(\u_cpu.ALU._0712_ ),
    .X(\u_cpu.ALU._0752_ ));
 sky130_fd_sc_hd__and4bb_2 \u_cpu.ALU._1606_  (.A_N(\u_cpu.ALU._0746_ ),
    .B_N(\u_cpu.ALU._0750_ ),
    .C(\u_cpu.ALU._0751_ ),
    .D(\u_cpu.ALU._0752_ ),
    .X(\u_cpu.ALU._0753_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1607_  (.A(\u_cpu.ALU._0753_ ),
    .X(\u_cpu.ALU._0754_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._1608_  (.A1(\u_cpu.ALU.SrcA[0] ),
    .A2(\u_cpu.ALU._0744_ ),
    .B1(\u_cpu.ALU._0749_ ),
    .C1(\u_cpu.ALU._0754_ ),
    .X(\u_cpu.ALU._0755_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1609_  (.A(\u_cpu.ALU._0755_ ),
    .B(\u_cpu.ALU._0723_ ),
    .Y(\u_cpu.ALU._0756_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1610_  (.A(\u_cpu.ALU._0613_ ),
    .X(\u_cpu.ALU._0757_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1611_  (.A(\u_cpu.ALU._0757_ ),
    .X(\u_cpu.ALU._0758_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1612_  (.A(\u_cpu.ALU._0758_ ),
    .X(\u_cpu.ALU._0759_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1613_  (.A(\u_cpu.ALU._0623_ ),
    .X(\u_cpu.ALU._0760_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1614_  (.A(\u_cpu.ALU._0760_ ),
    .X(\u_cpu.ALU._0761_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1615_  (.A0(\u_cpu.ALU.SrcA[28] ),
    .A1(\u_cpu.ALU._0579_ ),
    .A2(\u_cpu.ALU.SrcA[30] ),
    .A3(\u_cpu.ALU.SrcA[31] ),
    .S0(\u_cpu.ALU._0634_ ),
    .S1(\u_cpu.ALU._0725_ ),
    .X(\u_cpu.ALU._0762_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1616_  (.A0(\u_cpu.ALU._0433_ ),
    .A1(\u_cpu.ALU._0475_ ),
    .A2(\u_cpu.ALU.SrcA[26] ),
    .A3(\u_cpu.ALU._0338_ ),
    .S0(\u_cpu.ALU._0634_ ),
    .S1(\u_cpu.ALU._0725_ ),
    .X(\u_cpu.ALU._0763_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1617_  (.A(\u_cpu.ALU.SrcB[2] ),
    .Y(\u_cpu.ALU._0764_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1618_  (.A(\u_cpu.ALU._0764_ ),
    .X(\u_cpu.ALU._0765_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.ALU._1619_  (.A0(\u_cpu.ALU._0762_ ),
    .A1(\u_cpu.ALU._0763_ ),
    .S(\u_cpu.ALU._0765_ ),
    .X(\u_cpu.ALU._0766_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1620_  (.A0(\u_cpu.ALU.SrcA[20] ),
    .A1(\u_cpu.ALU.SrcA[21] ),
    .A2(\u_cpu.ALU._0560_ ),
    .A3(\u_cpu.ALU._0555_ ),
    .S0(\u_cpu.ALU._0720_ ),
    .S1(\u_cpu.ALU._0725_ ),
    .X(\u_cpu.ALU._0767_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1621_  (.A(\u_cpu.ALU._0764_ ),
    .X(\u_cpu.ALU._0768_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1622_  (.A(\u_cpu.ALU._0768_ ),
    .X(\u_cpu.ALU._0769_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1623_  (.A(\u_cpu.ALU._0647_ ),
    .X(\u_cpu.ALU._0770_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1624_  (.A(\u_cpu.ALU._0629_ ),
    .X(\u_cpu.ALU._0771_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1625_  (.A(\u_cpu.ALU._0637_ ),
    .X(\u_cpu.ALU._0772_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1626_  (.A(\u_cpu.ALU._0633_ ),
    .B(\u_cpu.ALU.SrcA[17] ),
    .X(\u_cpu.ALU._0773_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1627_  (.A1(\u_cpu.ALU._0641_ ),
    .A2(\u_cpu.ALU.SrcA[16] ),
    .B1(\u_cpu.ALU._0773_ ),
    .Y(\u_cpu.ALU._0774_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1628_  (.A(\u_cpu.ALU._0633_ ),
    .X(\u_cpu.ALU._0775_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1629_  (.A(\u_cpu.ALU._0720_ ),
    .B(\u_cpu.ALU.SrcA[19] ),
    .Y(\u_cpu.ALU._0776_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1630_  (.A1(\u_cpu.ALU._0775_ ),
    .A2(\u_cpu.ALU._0544_ ),
    .B1(\u_cpu.ALU._0776_ ),
    .Y(\u_cpu.ALU._0777_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1631_  (.A(\u_cpu.ALU._0777_ ),
    .B(\u_cpu.ALU._0638_ ),
    .Y(\u_cpu.ALU._0778_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1632_  (.A1(\u_cpu.ALU._0772_ ),
    .A2(\u_cpu.ALU._0774_ ),
    .B1(\u_cpu.ALU._0778_ ),
    .Y(\u_cpu.ALU._0779_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU._1633_  (.A(\u_cpu.ALU._0771_ ),
    .B(\u_cpu.ALU._0779_ ),
    .X(\u_cpu.ALU._0780_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._1634_  (.A1(\u_cpu.ALU._0767_ ),
    .A2(\u_cpu.ALU._0769_ ),
    .B1(\u_cpu.ALU._0770_ ),
    .C1(\u_cpu.ALU._0780_ ),
    .X(\u_cpu.ALU._0781_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1635_  (.A1(\u_cpu.ALU._0761_ ),
    .A2(\u_cpu.ALU._0766_ ),
    .B1(\u_cpu.ALU._0781_ ),
    .Y(\u_cpu.ALU._0782_ ));
 sky130_fd_sc_hd__or3b_2 \u_cpu.ALU._1636_  (.A(\u_cpu.ALU._0712_ ),
    .B(\u_cpu.ALU._0750_ ),
    .C_N(\u_cpu.ALU._0751_ ),
    .X(\u_cpu.ALU._0783_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1637_  (.A(\u_cpu.ALU._0783_ ),
    .X(\u_cpu.ALU._0784_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1638_  (.A(\u_cpu.ALU._0765_ ),
    .X(\u_cpu.ALU._0785_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1639_  (.A(\u_cpu.ALU._0785_ ),
    .X(\u_cpu.ALU._0786_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1640_  (.A(\u_cpu.ALU._0643_ ),
    .X(\u_cpu.ALU._0787_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1641_  (.A(\u_cpu.ALU._0634_ ),
    .B(\u_cpu.ALU.SrcA[3] ),
    .X(\u_cpu.ALU._0788_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._1642_  (.A1(\u_cpu.ALU._0641_ ),
    .A2(\u_cpu.ALU._0627_ ),
    .B1(\u_cpu.ALU._0787_ ),
    .C1(\u_cpu.ALU._0788_ ),
    .X(\u_cpu.ALU._0789_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1643_  (.A(\u_cpu.ALU._0772_ ),
    .X(\u_cpu.ALU._0790_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._1644_  (.A1(\u_cpu.ALU._0723_ ),
    .A2(\u_cpu.ALU._0632_ ),
    .B1(\u_cpu.ALU._0790_ ),
    .X(\u_cpu.ALU._0791_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1645_  (.A(\u_cpu.ALU._0721_ ),
    .B(\u_cpu.ALU._0608_ ),
    .X(\u_cpu.ALU._0792_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.ALU._1646_  (.A_N(\u_cpu.ALU._0634_ ),
    .B(\u_cpu.ALU.SrcA[4] ),
    .X(\u_cpu.ALU._0793_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1647_  (.A(\u_cpu.ALU._0775_ ),
    .X(\u_cpu.ALU._0794_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1648_  (.A(\u_cpu.ALU._0635_ ),
    .B(\u_cpu.ALU._0598_ ),
    .Y(\u_cpu.ALU._0795_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1649_  (.A1(\u_cpu.ALU._0794_ ),
    .A2(\u_cpu.ALU._0606_ ),
    .B1(\u_cpu.ALU._0795_ ),
    .C1(\u_cpu.ALU._0726_ ),
    .Y(\u_cpu.ALU._0796_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1650_  (.A(\u_cpu.ALU._0629_ ),
    .X(\u_cpu.ALU._0797_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU._1651_  (.A1(\u_cpu.ALU._0790_ ),
    .A2(\u_cpu.ALU._0792_ ),
    .A3(\u_cpu.ALU._0793_ ),
    .B1(\u_cpu.ALU._0796_ ),
    .C1(\u_cpu.ALU._0797_ ),
    .X(\u_cpu.ALU._0798_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU._1652_  (.A1(\u_cpu.ALU._0786_ ),
    .A2(\u_cpu.ALU._0789_ ),
    .A3(\u_cpu.ALU._0791_ ),
    .B1(\u_cpu.ALU._0798_ ),
    .Y(\u_cpu.ALU._0799_ ));
 sky130_fd_sc_hd__nor4_2 \u_cpu.ALU._1653_  (.A(\u_cpu.ALU.SrcB[0] ),
    .B(\u_cpu.ALU.SrcB[3] ),
    .C(\u_cpu.ALU.SrcB[2] ),
    .D(\u_cpu.ALU._0637_ ),
    .Y(\u_cpu.ALU._0800_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1654_  (.A(\u_cpu.ALU._0800_ ),
    .X(\u_cpu.ALU._0801_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1655_  (.A0(\u_cpu.ALU.SrcA[12] ),
    .A1(\u_cpu.ALU.SrcA[13] ),
    .A2(\u_cpu.ALU.SrcA[14] ),
    .A3(\u_cpu.ALU.SrcA[15] ),
    .S0(\u_cpu.ALU._0720_ ),
    .S1(\u_cpu.ALU._0725_ ),
    .X(\u_cpu.ALU._0802_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1656_  (.A0(\u_cpu.ALU.SrcA[8] ),
    .A1(\u_cpu.ALU.SrcA[9] ),
    .A2(\u_cpu.ALU.SrcA[10] ),
    .A3(\u_cpu.ALU.SrcA[11] ),
    .S0(\u_cpu.ALU._0720_ ),
    .S1(\u_cpu.ALU._0725_ ),
    .X(\u_cpu.ALU._0803_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.ALU._1657_  (.A0(\u_cpu.ALU._0802_ ),
    .A1(\u_cpu.ALU._0803_ ),
    .S(\u_cpu.ALU._0768_ ),
    .X(\u_cpu.ALU._0804_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1658_  (.A(\u_cpu.ALU._0623_ ),
    .X(\u_cpu.ALU._0805_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1659_  (.A(\u_cpu.ALU._0805_ ),
    .X(\u_cpu.ALU._0806_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.ALU._1660_  (.A1(\u_cpu.ALU.SrcA[0] ),
    .A2(\u_cpu.ALU._0801_ ),
    .B1(\u_cpu.ALU._0804_ ),
    .B2(\u_cpu.ALU._0806_ ),
    .C1(\u_cpu.ALU._0757_ ),
    .Y(\u_cpu.ALU._0807_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._1661_  (.A1(\u_cpu.ALU._0761_ ),
    .A2(\u_cpu.ALU._0799_ ),
    .B1(\u_cpu.ALU._0807_ ),
    .X(\u_cpu.ALU._0808_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._1662_  (.A1(\u_cpu.ALU._0759_ ),
    .A2(\u_cpu.ALU._0782_ ),
    .B1(\u_cpu.ALU._0784_ ),
    .C1(\u_cpu.ALU._0808_ ),
    .X(\u_cpu.ALU._0809_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1663_  (.A(_71943_),
    .Y(\u_cpu.ALU._0810_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1664_  (.A(\u_cpu.ALU._0810_ ),
    .X(\u_cpu.ALU._0811_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._1665_  (.A(\u_cpu.ALU._0737_ ),
    .B(\u_cpu.ALU._0711_ ),
    .C(\u_cpu.ALU._0811_ ),
    .X(\u_cpu.ALU._0812_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1666_  (.A(\u_cpu.ALU._0812_ ),
    .X(\u_cpu.ALU._0813_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU._1667_  (.A(_71944_),
    .B(_71945_),
    .C(\u_cpu.ALU._0735_ ),
    .Y(\u_cpu.ALU._0814_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1668_  (.A(\u_cpu.ALU.SrcA[0] ),
    .B(\u_cpu.ALU._0641_ ),
    .Y(\u_cpu.ALU._0815_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.ALU._1669_  (.A1(\u_cpu.ALU._0748_ ),
    .A2(\u_cpu.ALU._0813_ ),
    .A3(\u_cpu.ALU._0814_ ),
    .B1(\u_cpu.ALU._0815_ ),
    .B2(\u_cpu.ALU._0724_ ),
    .X(\u_cpu.ALU._0816_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1670_  (.A(\u_cpu.ALU._0613_ ),
    .Y(\u_cpu.ALU._0817_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU._1671_  (.A(\u_cpu.ALU._0817_ ),
    .B(\u_cpu.ALU._0736_ ),
    .C(\u_cpu.ALU._0712_ ),
    .D(\u_cpu.ALU._0746_ ),
    .X(\u_cpu.ALU._0818_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1672_  (.A(\u_cpu.ALU._0818_ ),
    .X(\u_cpu.ALU._0819_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.ALU._1673_  (.A_N(\u_cpu.ALU._0750_ ),
    .B(\u_cpu.ALU._0751_ ),
    .C(\u_cpu.ALU._0712_ ),
    .D(\u_cpu.ALU._0746_ ),
    .X(\u_cpu.ALU._0820_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1674_  (.A(\u_cpu.ALU._0820_ ),
    .X(\u_cpu.ALU._0821_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1675_  (.A(\u_cpu.ALU._0821_ ),
    .X(\u_cpu.ALU._0822_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU._1676_  (.A1(\u_cpu.ALU.SrcA[0] ),
    .A2(\u_cpu.ALU._0801_ ),
    .A3(\u_cpu.ALU._0819_ ),
    .B1(\u_cpu.ALU._0822_ ),
    .B2(\u_cpu.ALU.Product_Wallace[0] ),
    .X(\u_cpu.ALU._0823_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1677_  (.A(\u_cpu.ALU._0816_ ),
    .B(\u_cpu.ALU._0823_ ),
    .Y(\u_cpu.ALU._0824_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU._1678_  (.A(\u_cpu.ALU._0740_ ),
    .B(\u_cpu.ALU._0756_ ),
    .C(\u_cpu.ALU._0809_ ),
    .D(\u_cpu.ALU._0824_ ),
    .X(\u_cpu.ALU._0825_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1679_  (.A(\u_cpu.ALU._0825_ ),
    .Y(\u_cpu.ALU.ALUResult[0] ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1680_  (.A(\u_cpu.ALU._0725_ ),
    .X(\u_cpu.ALU._0826_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1681_  (.A(\u_cpu.ALU._0775_ ),
    .B(\u_cpu.ALU.SrcA[30] ),
    .Y(\u_cpu.ALU._0827_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._1682_  (.A1(\u_cpu.ALU._0721_ ),
    .A2(\u_cpu.ALU._0580_ ),
    .B1(\u_cpu.ALU._0827_ ),
    .X(\u_cpu.ALU._0828_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1683_  (.A(\u_cpu.ALU._0728_ ),
    .B(\u_cpu.ALU.SrcA[31] ),
    .Y(\u_cpu.ALU._0829_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1684_  (.A1(\u_cpu.ALU._0826_ ),
    .A2(\u_cpu.ALU._0828_ ),
    .B1(\u_cpu.ALU._0829_ ),
    .Y(\u_cpu.ALU._0830_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1685_  (.A(\u_cpu.ALU._0634_ ),
    .B(\u_cpu.ALU.SrcA[28] ),
    .X(\u_cpu.ALU._0831_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.ALU._1686_  (.A_N(\u_cpu.ALU._0634_ ),
    .B(\u_cpu.ALU.SrcA[27] ),
    .X(\u_cpu.ALU._0832_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.ALU._1687_  (.A(\u_cpu.ALU._0633_ ),
    .B_N(\u_cpu.ALU.SrcA[25] ),
    .X(\u_cpu.ALU._0833_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1688_  (.A1(\u_cpu.ALU._0641_ ),
    .A2(\u_cpu.ALU._0588_ ),
    .B1(\u_cpu.ALU._0833_ ),
    .C1(\u_cpu.ALU._0643_ ),
    .Y(\u_cpu.ALU._0834_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU._1689_  (.A1(\u_cpu.ALU._0787_ ),
    .A2(\u_cpu.ALU._0831_ ),
    .A3(\u_cpu.ALU._0832_ ),
    .B1(\u_cpu.ALU._0834_ ),
    .C1(\u_cpu.ALU._0765_ ),
    .X(\u_cpu.ALU._0835_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1690_  (.A1(\u_cpu.ALU._0830_ ),
    .A2(\u_cpu.ALU._0797_ ),
    .B1(\u_cpu.ALU._0835_ ),
    .Y(\u_cpu.ALU._0836_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1691_  (.A(\u_cpu.ALU.SrcA[20] ),
    .X(\u_cpu.ALU._0837_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1692_  (.A(\u_cpu.ALU._0720_ ),
    .X(\u_cpu.ALU._0838_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1693_  (.A0(\u_cpu.ALU._0536_ ),
    .A1(\u_cpu.ALU.SrcA[18] ),
    .A2(\u_cpu.ALU.SrcA[19] ),
    .A3(\u_cpu.ALU._0837_ ),
    .S0(\u_cpu.ALU._0838_ ),
    .S1(\u_cpu.ALU._0728_ ),
    .X(\u_cpu.ALU._0839_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1694_  (.A(\u_cpu.ALU._0633_ ),
    .X(\u_cpu.ALU._0840_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1695_  (.A(\u_cpu.ALU._0634_ ),
    .B(\u_cpu.ALU._0433_ ),
    .Y(\u_cpu.ALU._0841_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1696_  (.A1(\u_cpu.ALU._0840_ ),
    .A2(\u_cpu.ALU._0552_ ),
    .B1(\u_cpu.ALU._0841_ ),
    .Y(\u_cpu.ALU._0842_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.ALU._1697_  (.A(\u_cpu.ALU._0633_ ),
    .B_N(\u_cpu.ALU.SrcA[21] ),
    .X(\u_cpu.ALU._0843_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1698_  (.A(\u_cpu.ALU._0775_ ),
    .B(\u_cpu.ALU._0560_ ),
    .Y(\u_cpu.ALU._0844_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1699_  (.A1(\u_cpu.ALU._0843_ ),
    .A2(\u_cpu.ALU._0844_ ),
    .B1(\u_cpu.ALU._0638_ ),
    .Y(\u_cpu.ALU._0845_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._1700_  (.A1(\u_cpu.ALU._0726_ ),
    .A2(\u_cpu.ALU._0842_ ),
    .B1(\u_cpu.ALU._0765_ ),
    .C1(\u_cpu.ALU._0845_ ),
    .X(\u_cpu.ALU._0846_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1701_  (.A1(\u_cpu.ALU._0797_ ),
    .A2(\u_cpu.ALU._0839_ ),
    .B1(\u_cpu.ALU._0846_ ),
    .C1(\u_cpu.ALU._0770_ ),
    .Y(\u_cpu.ALU._0847_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1702_  (.A1(\u_cpu.ALU._0770_ ),
    .A2(\u_cpu.ALU._0836_ ),
    .B1(\u_cpu.ALU._0847_ ),
    .Y(\u_cpu.ALU._0848_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1703_  (.A(\u_cpu.ALU.SrcA[3] ),
    .Y(\u_cpu.ALU._0849_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1704_  (.A(\u_cpu.ALU._0721_ ),
    .B(\u_cpu.ALU._0618_ ),
    .Y(\u_cpu.ALU._0850_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1705_  (.A1(\u_cpu.ALU._0635_ ),
    .A2(\u_cpu.ALU._0849_ ),
    .B1(\u_cpu.ALU._0850_ ),
    .Y(\u_cpu.ALU._0851_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU._1706_  (.A1(\u_cpu.ALU._0838_ ),
    .A2(\u_cpu.ALU.SrcA[1] ),
    .B1_N(\u_cpu.ALU._0637_ ),
    .Y(\u_cpu.ALU._0852_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1707_  (.A1(\u_cpu.ALU._0648_ ),
    .A2(\u_cpu.ALU._0794_ ),
    .B1(\u_cpu.ALU._0852_ ),
    .Y(\u_cpu.ALU._0853_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1708_  (.A1(\u_cpu.ALU._0851_ ),
    .A2(\u_cpu.ALU._0826_ ),
    .B1(\u_cpu.ALU._0853_ ),
    .Y(\u_cpu.ALU._0854_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._1709_  (.A1(\u_cpu.ALU._0771_ ),
    .A2(\u_cpu.ALU._0854_ ),
    .B1(\u_cpu.ALU._0647_ ),
    .X(\u_cpu.ALU._0855_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1710_  (.A0(\u_cpu.ALU._0608_ ),
    .A1(\u_cpu.ALU.SrcA[6] ),
    .A2(\u_cpu.ALU._0598_ ),
    .A3(\u_cpu.ALU._0663_ ),
    .S0(\u_cpu.ALU._0721_ ),
    .S1(\u_cpu.ALU._0772_ ),
    .X(\u_cpu.ALU._0856_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1711_  (.A(\u_cpu.ALU._0797_ ),
    .B(\u_cpu.ALU._0856_ ),
    .Y(\u_cpu.ALU._0857_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1712_  (.A(\u_cpu.ALU.SrcA[11] ),
    .Y(\u_cpu.ALU._0858_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1713_  (.A(\u_cpu.ALU.SrcA[12] ),
    .X(\u_cpu.ALU._0859_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1714_  (.A(\u_cpu.ALU._0838_ ),
    .B(\u_cpu.ALU._0859_ ),
    .Y(\u_cpu.ALU._0860_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._1715_  (.A1(\u_cpu.ALU._0721_ ),
    .A2(\u_cpu.ALU._0858_ ),
    .B1(\u_cpu.ALU._0860_ ),
    .C1(\u_cpu.ALU._0638_ ),
    .X(\u_cpu.ALU._0861_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1716_  (.A(\u_cpu.ALU.SrcA[9] ),
    .Y(\u_cpu.ALU._0862_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1717_  (.A(\u_cpu.ALU._0838_ ),
    .B(\u_cpu.ALU.SrcA[10] ),
    .Y(\u_cpu.ALU._0863_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._1718_  (.A1(\u_cpu.ALU._0635_ ),
    .A2(\u_cpu.ALU._0862_ ),
    .B1(\u_cpu.ALU._0863_ ),
    .C1(\u_cpu.ALU._0643_ ),
    .X(\u_cpu.ALU._0864_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.ALU._1719_  (.A_N(\u_cpu.ALU._0775_ ),
    .B(\u_cpu.ALU.SrcA[13] ),
    .X(\u_cpu.ALU._0865_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1720_  (.A(\u_cpu.ALU._0775_ ),
    .B(\u_cpu.ALU.SrcA[14] ),
    .X(\u_cpu.ALU._0866_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1721_  (.A(\u_cpu.ALU._0840_ ),
    .B(\u_cpu.ALU.SrcA[16] ),
    .Y(\u_cpu.ALU._0867_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1722_  (.A1(\u_cpu.ALU._0721_ ),
    .A2(\u_cpu.ALU._0683_ ),
    .B1(\u_cpu.ALU._0867_ ),
    .C1(\u_cpu.ALU._0638_ ),
    .Y(\u_cpu.ALU._0868_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.ALU._1723_  (.A1(\u_cpu.ALU._0728_ ),
    .A2(\u_cpu.ALU._0865_ ),
    .A3(\u_cpu.ALU._0866_ ),
    .B1(\u_cpu.ALU._0868_ ),
    .C1(\u_cpu.ALU._0629_ ),
    .Y(\u_cpu.ALU._0869_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU._1724_  (.A1(\u_cpu.ALU._0771_ ),
    .A2(\u_cpu.ALU._0861_ ),
    .A3(\u_cpu.ALU._0864_ ),
    .B1(\u_cpu.ALU._0869_ ),
    .C1(\u_cpu.ALU._0805_ ),
    .X(\u_cpu.ALU._0870_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU._1725_  (.A1(\u_cpu.ALU._0855_ ),
    .A2(\u_cpu.ALU._0857_ ),
    .B1(\u_cpu.ALU._0757_ ),
    .C1(\u_cpu.ALU._0870_ ),
    .Y(\u_cpu.ALU._0871_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._1726_  (.A1(\u_cpu.ALU._0757_ ),
    .A2(\u_cpu.ALU._0848_ ),
    .B1(\u_cpu.ALU._0871_ ),
    .X(\u_cpu.ALU._0872_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1727_  (.A(\u_cpu.ALU._0711_ ),
    .X(\u_cpu.ALU._0873_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1728_  (.A(\u_cpu.ALU._0873_ ),
    .B(\u_cpu.ALU._0783_ ),
    .Y(\u_cpu.ALU._0874_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1729_  (.A(\u_cpu.ALU._0872_ ),
    .B(\u_cpu.ALU._0874_ ),
    .Y(\u_cpu.ALU._0875_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU._1730_  (.A1(\u_cpu.ALU._0829_ ),
    .A2(\u_cpu.ALU._0722_ ),
    .B1(\u_cpu.ALU._0826_ ),
    .B2(\u_cpu.ALU._0828_ ),
    .X(\u_cpu.ALU._0876_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU._1731_  (.A1(\u_cpu.ALU._0785_ ),
    .A2(\u_cpu.ALU._0876_ ),
    .B1_N(\u_cpu.ALU._0835_ ),
    .Y(\u_cpu.ALU._0877_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1732_  (.A(\u_cpu.ALU._0877_ ),
    .B(\u_cpu.ALU._0806_ ),
    .Y(\u_cpu.ALU._0878_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1733_  (.A(\u_cpu.ALU._0817_ ),
    .X(\u_cpu.ALU._0879_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1734_  (.A1(\u_cpu.ALU._0847_ ),
    .A2(\u_cpu.ALU._0878_ ),
    .B1(\u_cpu.ALU._0879_ ),
    .Y(\u_cpu.ALU._0880_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1735_  (.A(\u_cpu.ALU._0746_ ),
    .X(\u_cpu.ALU._0881_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1736_  (.A(\u_cpu.ALU._0881_ ),
    .B(\u_cpu.ALU._0783_ ),
    .Y(\u_cpu.ALU._0882_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1737_  (.A1(\u_cpu.ALU._0871_ ),
    .A2(\u_cpu.ALU._0880_ ),
    .B1(\u_cpu.ALU._0882_ ),
    .Y(\u_cpu.ALU._0883_ ));
 sky130_fd_sc_hd__nor4b_2 \u_cpu.ALU._1738_  (.A(_71946_),
    .B(_71947_),
    .C(\u_cpu.ALU._0735_ ),
    .D_N(_71948_),
    .Y(\u_cpu.ALU._0884_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU._1739_  (.A1(\u_cpu.ALU._0640_ ),
    .A2(\u_cpu.ALU._0884_ ),
    .B1_N(\u_cpu.ALU._0642_ ),
    .Y(\u_cpu.ALU._0885_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._1740_  (.A(\u_cpu.ALU._0741_ ),
    .B(\u_cpu.ALU._0810_ ),
    .C(\u_cpu.ALU._0745_ ),
    .Y(\u_cpu.ALU._0886_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._1741_  (.A(\u_cpu.ALU._0886_ ),
    .B(\u_cpu.ALU._0633_ ),
    .C(\u_cpu.ALU._0642_ ),
    .Y(\u_cpu.ALU._0887_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1742_  (.A1(\u_cpu.ALU._0885_ ),
    .A2(\u_cpu.ALU._0887_ ),
    .B1(\u_cpu.ALU.SrcA[1] ),
    .Y(\u_cpu.ALU._0888_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._1743_  (.A(\u_cpu.ALU._0885_ ),
    .B(\u_cpu.ALU._0887_ ),
    .C(\u_cpu.ALU._0632_ ),
    .X(\u_cpu.ALU._0889_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1744_  (.A(\u_cpu.ALU._0811_ ),
    .X(\u_cpu.ALU._0890_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU._1745_  (.A1(\u_cpu.ALU._0815_ ),
    .A2(\u_cpu.ALU._0888_ ),
    .A3(\u_cpu.ALU._0889_ ),
    .B1(\u_cpu.ALU._0742_ ),
    .C1(\u_cpu.ALU._0890_ ),
    .X(\u_cpu.ALU._0891_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1746_  (.A1(\u_cpu.ALU._0888_ ),
    .A2(\u_cpu.ALU._0889_ ),
    .B1(\u_cpu.ALU._0815_ ),
    .Y(\u_cpu.ALU._0892_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._1747_  (.A1(\u_cpu.ALU._0794_ ),
    .A2(\u_cpu.ALU._0632_ ),
    .B1(\u_cpu.ALU._0787_ ),
    .C1(\u_cpu.ALU._0732_ ),
    .X(\u_cpu.ALU._0893_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._1748_  (.A(\u_cpu.ALU._0893_ ),
    .B(\u_cpu.ALU._0768_ ),
    .C(\u_cpu.ALU._0647_ ),
    .X(\u_cpu.ALU._0894_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1749_  (.A(\u_cpu.ALU._0750_ ),
    .B(\u_cpu.ALU._0713_ ),
    .Y(\u_cpu.ALU._0895_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1750_  (.A(\u_cpu.ALU._0895_ ),
    .X(\u_cpu.ALU._0896_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._1751_  (.A1(\u_cpu.ALU._0751_ ),
    .A2(\u_cpu.ALU._0632_ ),
    .B1(\u_cpu.ALU._0790_ ),
    .C1(\u_cpu.ALU._0896_ ),
    .X(\u_cpu.ALU._0897_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._1752_  (.A1(\u_cpu.ALU.Product_Wallace[1] ),
    .A2(\u_cpu.ALU._0820_ ),
    .B1(\u_cpu.ALU._0894_ ),
    .B2(\u_cpu.ALU._0819_ ),
    .C1(\u_cpu.ALU._0897_ ),
    .X(\u_cpu.ALU._0898_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1753_  (.A(\u_cpu.ALU._0729_ ),
    .X(\u_cpu.ALU._0899_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1754_  (.A(\u_cpu.ALU._0711_ ),
    .X(\u_cpu.ALU._0900_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU._1755_  (.A(\u_cpu.ALU._0737_ ),
    .B(\u_cpu.ALU._0730_ ),
    .C(\u_cpu.ALU._0811_ ),
    .D(\u_cpu.ALU._0900_ ),
    .X(\u_cpu.ALU._0901_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU._1756_  (.A1(\u_cpu.ALU._0632_ ),
    .A2(\u_cpu.ALU._0899_ ),
    .B1(\u_cpu.ALU._0748_ ),
    .B2(\u_cpu.ALU._0901_ ),
    .X(\u_cpu.ALU._0902_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU._1757_  (.A1(\u_cpu.ALU._0891_ ),
    .A2(\u_cpu.ALU._0892_ ),
    .B1(\u_cpu.ALU._0898_ ),
    .C1(\u_cpu.ALU._0902_ ),
    .Y(\u_cpu.ALU._0903_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._1758_  (.A(\u_cpu.ALU._0875_ ),
    .B(\u_cpu.ALU._0883_ ),
    .C(\u_cpu.ALU._0903_ ),
    .X(\u_cpu.ALU._0904_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1759_  (.A(\u_cpu.ALU._0904_ ),
    .Y(\u_cpu.ALU.ALUResult[1] ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU._1760_  (.A1(\u_cpu.ALU._0741_ ),
    .A2(\u_cpu.ALU._0810_ ),
    .A3(\u_cpu.ALU._0745_ ),
    .B1(\u_cpu.ALU._0641_ ),
    .Y(\u_cpu.ALU._0905_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1761_  (.A1(\u_cpu.ALU._0642_ ),
    .A2(\u_cpu.ALU._0905_ ),
    .B1(\u_cpu.ALU.SrcA[1] ),
    .Y(\u_cpu.ALU._0906_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU._1762_  (.A1(_71949_),
    .A2(\u_cpu.ALU._0735_ ),
    .A3(\u_cpu.ALU._0707_ ),
    .B1(\u_cpu.ALU._0642_ ),
    .C1(\u_cpu.ALU._0633_ ),
    .X(\u_cpu.ALU._0907_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU._1763_  (.A1(\u_cpu.ALU._0906_ ),
    .A2(\u_cpu.ALU._0907_ ),
    .B1(\u_cpu.ALU._0815_ ),
    .B2(\u_cpu.ALU._0888_ ),
    .Y(\u_cpu.ALU._0908_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU._1764_  (.A(_71950_),
    .B(\u_cpu.ALU._0735_ ),
    .X(\u_cpu.ALU._0909_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU._1765_  (.A1(\u_cpu.ALU._0633_ ),
    .A2(\u_cpu.ALU._0637_ ),
    .B1(\u_cpu.ALU._0707_ ),
    .B2(\u_cpu.ALU._0909_ ),
    .C1(\u_cpu.ALU.SrcB[2] ),
    .Y(\u_cpu.ALU._0910_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1766_  (.A(\u_cpu.ALU.SrcB[0] ),
    .B(\u_cpu.ALU.SrcB[1] ),
    .Y(\u_cpu.ALU._0911_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._1767_  (.A1(\u_cpu.ALU._0741_ ),
    .A2(\u_cpu.ALU._0810_ ),
    .A3(\u_cpu.ALU._0745_ ),
    .B1(\u_cpu.ALU._0911_ ),
    .X(\u_cpu.ALU._0912_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1768_  (.A1(\u_cpu.ALU._0764_ ),
    .A2(\u_cpu.ALU._0912_ ),
    .B1(\u_cpu.ALU._0627_ ),
    .Y(\u_cpu.ALU._0913_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1769_  (.A(\u_cpu.ALU._0884_ ),
    .X(\u_cpu.ALU._0914_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1770_  (.A1(\u_cpu.ALU._0911_ ),
    .A2(\u_cpu.ALU._0914_ ),
    .B1(\u_cpu.ALU._0764_ ),
    .Y(\u_cpu.ALU._0915_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1771_  (.A1(\u_cpu.ALU._0915_ ),
    .A2(\u_cpu.ALU._0910_ ),
    .B1(\u_cpu.ALU._0648_ ),
    .Y(\u_cpu.ALU._0916_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1772_  (.A1(\u_cpu.ALU._0910_ ),
    .A2(\u_cpu.ALU._0913_ ),
    .B1(\u_cpu.ALU._0916_ ),
    .Y(\u_cpu.ALU._0917_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1773_  (.A(\u_cpu.ALU._0908_ ),
    .B(\u_cpu.ALU._0917_ ),
    .Y(\u_cpu.ALU._0918_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1774_  (.A(\u_cpu.ALU._0741_ ),
    .B(\u_cpu.ALU._0810_ ),
    .Y(\u_cpu.ALU._0919_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1775_  (.A(\u_cpu.ALU._0919_ ),
    .X(\u_cpu.ALU._0920_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1776_  (.A(\u_cpu.ALU._0920_ ),
    .X(\u_cpu.ALU._0921_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._1777_  (.A1(\u_cpu.ALU._0917_ ),
    .A2(\u_cpu.ALU._0908_ ),
    .B1(\u_cpu.ALU._0921_ ),
    .X(\u_cpu.ALU._0922_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1778_  (.A(\u_cpu.ALU._0720_ ),
    .B(\u_cpu.ALU.SrcA[27] ),
    .X(\u_cpu.ALU._0923_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.ALU._1779_  (.A_N(\u_cpu.ALU._0720_ ),
    .B(\u_cpu.ALU.SrcA[26] ),
    .X(\u_cpu.ALU._0924_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1780_  (.A(\u_cpu.ALU.SrcA[28] ),
    .Y(\u_cpu.ALU._0925_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1781_  (.A(\u_cpu.ALU._0634_ ),
    .B(\u_cpu.ALU._0579_ ),
    .Y(\u_cpu.ALU._0926_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1782_  (.A1(\u_cpu.ALU._0775_ ),
    .A2(\u_cpu.ALU._0925_ ),
    .B1(\u_cpu.ALU._0926_ ),
    .C1(\u_cpu.ALU._0725_ ),
    .Y(\u_cpu.ALU._0927_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.ALU._1783_  (.A1(\u_cpu.ALU._0826_ ),
    .A2(\u_cpu.ALU._0923_ ),
    .A3(\u_cpu.ALU._0924_ ),
    .B1(\u_cpu.ALU._0927_ ),
    .Y(\u_cpu.ALU._0928_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1784_  (.A(\u_cpu.ALU._0720_ ),
    .B(\u_cpu.ALU.SrcA[31] ),
    .X(\u_cpu.ALU._0929_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1785_  (.A1(\u_cpu.ALU._0641_ ),
    .A2(\u_cpu.ALU._0516_ ),
    .B1(\u_cpu.ALU._0929_ ),
    .Y(\u_cpu.ALU._0930_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU._1786_  (.A_N(\u_cpu.ALU._0930_ ),
    .B(\u_cpu.ALU._0771_ ),
    .C(\u_cpu.ALU._0787_ ),
    .Y(\u_cpu.ALU._0931_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1787_  (.A1(\u_cpu.ALU._0797_ ),
    .A2(\u_cpu.ALU._0928_ ),
    .B1(\u_cpu.ALU._0931_ ),
    .Y(\u_cpu.ALU._0932_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.ALU._1788_  (.A0(\u_cpu.ALU.SrcA[24] ),
    .A1(\u_cpu.ALU.SrcA[25] ),
    .S(\u_cpu.ALU._0720_ ),
    .X(\u_cpu.ALU._0933_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1789_  (.A(\u_cpu.ALU._0634_ ),
    .B(\u_cpu.ALU.SrcA[23] ),
    .Y(\u_cpu.ALU._0934_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1790_  (.A1(\u_cpu.ALU._0840_ ),
    .A2(\u_cpu.ALU._0562_ ),
    .B1(\u_cpu.ALU._0934_ ),
    .C1(\u_cpu.ALU._0643_ ),
    .Y(\u_cpu.ALU._0935_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1791_  (.A1(\u_cpu.ALU._0787_ ),
    .A2(\u_cpu.ALU._0933_ ),
    .B1(\u_cpu.ALU._0935_ ),
    .C1(\u_cpu.ALU._0629_ ),
    .Y(\u_cpu.ALU._0936_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1792_  (.A(\u_cpu.ALU._0840_ ),
    .B(\u_cpu.ALU.SrcA[21] ),
    .X(\u_cpu.ALU._0937_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1793_  (.A(\u_cpu.ALU._0635_ ),
    .B(\u_cpu.ALU._0570_ ),
    .Y(\u_cpu.ALU._0938_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1794_  (.A1(\u_cpu.ALU._0635_ ),
    .A2(\u_cpu.ALU._0544_ ),
    .B1(\u_cpu.ALU._0776_ ),
    .C1(\u_cpu.ALU._0643_ ),
    .Y(\u_cpu.ALU._0939_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.ALU._1795_  (.A1(\u_cpu.ALU._0787_ ),
    .A2(\u_cpu.ALU._0937_ ),
    .A3(\u_cpu.ALU._0938_ ),
    .B1(\u_cpu.ALU._0939_ ),
    .C1(\u_cpu.ALU._0765_ ),
    .Y(\u_cpu.ALU._0940_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1796_  (.A1(\u_cpu.ALU._0936_ ),
    .A2(\u_cpu.ALU._0940_ ),
    .B1(\u_cpu.ALU._0805_ ),
    .Y(\u_cpu.ALU._0941_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1797_  (.A1(\u_cpu.ALU._0760_ ),
    .A2(\u_cpu.ALU._0932_ ),
    .B1(\u_cpu.ALU._0941_ ),
    .Y(\u_cpu.ALU._0942_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1798_  (.A0(\u_cpu.ALU._0627_ ),
    .A1(\u_cpu.ALU._0624_ ),
    .A2(\u_cpu.ALU._0618_ ),
    .A3(\u_cpu.ALU._0608_ ),
    .S0(\u_cpu.ALU._0840_ ),
    .S1(\u_cpu.ALU._0728_ ),
    .X(\u_cpu.ALU._0943_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1799_  (.A(\u_cpu.ALU._0785_ ),
    .B(\u_cpu.ALU._0943_ ),
    .Y(\u_cpu.ALU._0944_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1800_  (.A0(\u_cpu.ALU.SrcA[6] ),
    .A1(\u_cpu.ALU._0598_ ),
    .A2(\u_cpu.ALU._0663_ ),
    .A3(\u_cpu.ALU._0669_ ),
    .S0(\u_cpu.ALU._0840_ ),
    .S1(\u_cpu.ALU._0728_ ),
    .X(\u_cpu.ALU._0945_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1801_  (.A(\u_cpu.ALU._0797_ ),
    .B(\u_cpu.ALU._0945_ ),
    .Y(\u_cpu.ALU._0946_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._1802_  (.A(\u_cpu.ALU._0770_ ),
    .B(\u_cpu.ALU._0944_ ),
    .C(\u_cpu.ALU._0946_ ),
    .Y(\u_cpu.ALU._0947_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1803_  (.A(\u_cpu.ALU.SrcA[15] ),
    .X(\u_cpu.ALU._0948_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1804_  (.A0(\u_cpu.ALU._0679_ ),
    .A1(\u_cpu.ALU._0948_ ),
    .A2(\u_cpu.ALU.SrcA[16] ),
    .A3(\u_cpu.ALU.SrcA[17] ),
    .S0(\u_cpu.ALU._0840_ ),
    .S1(\u_cpu.ALU._0638_ ),
    .X(\u_cpu.ALU._0949_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1805_  (.A(\u_cpu.ALU._0771_ ),
    .B(\u_cpu.ALU._0949_ ),
    .Y(\u_cpu.ALU._0950_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1806_  (.A0(\u_cpu.ALU.SrcA[10] ),
    .A1(\u_cpu.ALU._0686_ ),
    .A2(\u_cpu.ALU._0859_ ),
    .A3(\u_cpu.ALU.SrcA[13] ),
    .S0(\u_cpu.ALU._0840_ ),
    .S1(\u_cpu.ALU._0638_ ),
    .X(\u_cpu.ALU._0951_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1807_  (.A(\u_cpu.ALU._0951_ ),
    .B(\u_cpu.ALU._0768_ ),
    .Y(\u_cpu.ALU._0952_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._1808_  (.A(\u_cpu.ALU._0950_ ),
    .B(\u_cpu.ALU._0760_ ),
    .C(\u_cpu.ALU._0952_ ),
    .Y(\u_cpu.ALU._0953_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._1809_  (.A(\u_cpu.ALU._0817_ ),
    .B(\u_cpu.ALU._0947_ ),
    .C(\u_cpu.ALU._0953_ ),
    .Y(\u_cpu.ALU._0954_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1810_  (.A1(\u_cpu.ALU._0879_ ),
    .A2(\u_cpu.ALU._0942_ ),
    .B1(\u_cpu.ALU._0954_ ),
    .Y(\u_cpu.ALU._0955_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU._1811_  (.A1_N(\u_cpu.ALU._0918_ ),
    .A2_N(\u_cpu.ALU._0922_ ),
    .B1(\u_cpu.ALU._0882_ ),
    .B2(\u_cpu.ALU._0955_ ),
    .Y(\u_cpu.ALU._0956_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1812_  (.A(\u_cpu.ALU._0751_ ),
    .X(\u_cpu.ALU._0957_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1813_  (.A(\u_cpu.ALU._0629_ ),
    .X(\u_cpu.ALU._0958_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._1814_  (.A1(\u_cpu.ALU._0957_ ),
    .A2(\u_cpu.ALU._0627_ ),
    .B1(\u_cpu.ALU._0896_ ),
    .C1(\u_cpu.ALU._0958_ ),
    .X(\u_cpu.ALU._0959_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1815_  (.A(\u_cpu.ALU.SrcB[3] ),
    .B(\u_cpu.ALU.SrcB[2] ),
    .Y(\u_cpu.ALU._0960_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.ALU._1816_  (.A0(\u_cpu.ALU._0627_ ),
    .A1(\u_cpu.ALU._0632_ ),
    .S(\u_cpu.ALU._0838_ ),
    .X(\u_cpu.ALU._0961_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._1817_  (.A1(\u_cpu.ALU._0826_ ),
    .A2(\u_cpu.ALU._0961_ ),
    .B1(\u_cpu.ALU._0639_ ),
    .X(\u_cpu.ALU._0962_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1818_  (.A(\u_cpu.ALU._0752_ ),
    .X(\u_cpu.ALU._0963_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU._1819_  (.A1(\u_cpu.ALU._0963_ ),
    .A2(\u_cpu.ALU._0881_ ),
    .A3(\u_cpu.ALU._0742_ ),
    .B1(\u_cpu.ALU._0812_ ),
    .B2(\u_cpu.ALU._0630_ ),
    .X(\u_cpu.ALU._0964_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU._1820_  (.A1(\u_cpu.ALU._0960_ ),
    .A2(\u_cpu.ALU._0819_ ),
    .A3(\u_cpu.ALU._0962_ ),
    .B1(\u_cpu.ALU._0964_ ),
    .B2(\u_cpu.ALU._0628_ ),
    .X(\u_cpu.ALU._0965_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU._1821_  (.A1(\u_cpu.ALU.Product_Wallace[2] ),
    .A2(\u_cpu.ALU._0821_ ),
    .B1(\u_cpu.ALU._0959_ ),
    .C1(\u_cpu.ALU._0965_ ),
    .Y(\u_cpu.ALU._0966_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._1822_  (.A1(\u_cpu.ALU._0726_ ),
    .A2(\u_cpu.ALU._0930_ ),
    .B1(\u_cpu.ALU._0829_ ),
    .X(\u_cpu.ALU._0967_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU._1823_  (.A1(\u_cpu.ALU._0728_ ),
    .A2(\u_cpu.ALU._0923_ ),
    .A3(\u_cpu.ALU._0924_ ),
    .B1(\u_cpu.ALU._0927_ ),
    .X(\u_cpu.ALU._0968_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1824_  (.A(\u_cpu.ALU._0968_ ),
    .B(\u_cpu.ALU._0785_ ),
    .Y(\u_cpu.ALU._0969_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1825_  (.A1(\u_cpu.ALU._0785_ ),
    .A2(\u_cpu.ALU._0967_ ),
    .B1(\u_cpu.ALU._0969_ ),
    .Y(\u_cpu.ALU._0970_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1826_  (.A1(\u_cpu.ALU._0970_ ),
    .A2(\u_cpu.ALU._0806_ ),
    .B1(\u_cpu.ALU._0941_ ),
    .Y(\u_cpu.ALU._0971_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1827_  (.A1(\u_cpu.ALU._0879_ ),
    .A2(\u_cpu.ALU._0971_ ),
    .B1(\u_cpu.ALU._0954_ ),
    .Y(\u_cpu.ALU._0972_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1828_  (.A(\u_cpu.ALU._0972_ ),
    .B(\u_cpu.ALU._0874_ ),
    .Y(\u_cpu.ALU._0973_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._1829_  (.A(\u_cpu.ALU._0956_ ),
    .B(\u_cpu.ALU._0966_ ),
    .C(\u_cpu.ALU._0973_ ),
    .X(\u_cpu.ALU._0974_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1830_  (.A(\u_cpu.ALU._0974_ ),
    .Y(\u_cpu.ALU.ALUResult[2] ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1831_  (.A(\u_cpu.ALU._0814_ ),
    .X(\u_cpu.ALU._0975_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU._1832_  (.A(\u_cpu.ALU.SrcB[0] ),
    .B(\u_cpu.ALU.SrcB[2] ),
    .C(\u_cpu.ALU._0637_ ),
    .Y(\u_cpu.ALU._0976_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._1833_  (.A1(\u_cpu.ALU._0745_ ),
    .A2(\u_cpu.ALU._0741_ ),
    .A3(\u_cpu.ALU._0810_ ),
    .B1(\u_cpu.ALU._0976_ ),
    .X(\u_cpu.ALU._0977_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1834_  (.A1(\u_cpu.ALU._0646_ ),
    .A2(\u_cpu.ALU._0977_ ),
    .B1(\u_cpu.ALU.SrcA[3] ),
    .Y(\u_cpu.ALU._0978_ ));
 sky130_fd_sc_hd__a311o_2 \u_cpu.ALU._1835_  (.A1(\u_cpu.ALU._0741_ ),
    .A2(\u_cpu.ALU._0811_ ),
    .A3(\u_cpu.ALU._0745_ ),
    .B1(\u_cpu.ALU._0646_ ),
    .C1(\u_cpu.ALU._0976_ ),
    .X(\u_cpu.ALU._0979_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1836_  (.A(\u_cpu.ALU._0917_ ),
    .B(\u_cpu.ALU._0908_ ),
    .Y(\u_cpu.ALU._0980_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._1837_  (.A1(\u_cpu.ALU._0915_ ),
    .A2(\u_cpu.ALU._0910_ ),
    .B1(\u_cpu.ALU._0648_ ),
    .X(\u_cpu.ALU._0981_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1838_  (.A1(\u_cpu.ALU._0914_ ),
    .A2(\u_cpu.ALU._0976_ ),
    .B1(\u_cpu.ALU._0646_ ),
    .Y(\u_cpu.ALU._0982_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1839_  (.A1(\u_cpu.ALU._0982_ ),
    .A2(\u_cpu.ALU._0979_ ),
    .B1(\u_cpu.ALU._0849_ ),
    .Y(\u_cpu.ALU._0983_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._1840_  (.A1(\u_cpu.ALU._0978_ ),
    .A2(\u_cpu.ALU._0979_ ),
    .B1(\u_cpu.ALU._0980_ ),
    .B2(\u_cpu.ALU._0981_ ),
    .C1(\u_cpu.ALU._0983_ ),
    .X(\u_cpu.ALU._0984_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1841_  (.A(\u_cpu.ALU._0886_ ),
    .X(\u_cpu.ALU._0985_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1842_  (.A(\u_cpu.ALU._0911_ ),
    .B(\u_cpu.ALU._0764_ ),
    .Y(\u_cpu.ALU._0986_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1843_  (.A1(\u_cpu.ALU._0985_ ),
    .A2(\u_cpu.ALU._0986_ ),
    .B1(\u_cpu.ALU._0623_ ),
    .Y(\u_cpu.ALU._0987_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU._1844_  (.A1(\u_cpu.ALU._0633_ ),
    .A2(\u_cpu.ALU.SrcB[2] ),
    .A3(\u_cpu.ALU._0637_ ),
    .B1(\u_cpu.ALU._0623_ ),
    .C1(\u_cpu.ALU._0985_ ),
    .X(\u_cpu.ALU._0988_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1845_  (.A1(\u_cpu.ALU._0987_ ),
    .A2(\u_cpu.ALU._0988_ ),
    .B1(\u_cpu.ALU._0624_ ),
    .Y(\u_cpu.ALU._0989_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1846_  (.A1(\u_cpu.ALU._0646_ ),
    .A2(\u_cpu.ALU._0977_ ),
    .B1(\u_cpu.ALU._0978_ ),
    .Y(\u_cpu.ALU._0990_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._1847_  (.A1(\u_cpu.ALU._0989_ ),
    .A2(\u_cpu.ALU._0990_ ),
    .B1(\u_cpu.ALU._0917_ ),
    .B2(\u_cpu.ALU._0908_ ),
    .C1(\u_cpu.ALU._0916_ ),
    .X(\u_cpu.ALU._0991_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1848_  (.A1(\u_cpu.ALU._0641_ ),
    .A2(\u_cpu.ALU._0588_ ),
    .B1(\u_cpu.ALU._0833_ ),
    .C1(\u_cpu.ALU._0772_ ),
    .Y(\u_cpu.ALU._0992_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1849_  (.A1(\u_cpu.ALU._0826_ ),
    .A2(\u_cpu.ALU._0842_ ),
    .B1(\u_cpu.ALU._0992_ ),
    .Y(\u_cpu.ALU._0993_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1850_  (.A(\u_cpu.ALU.SrcA[31] ),
    .Y(\u_cpu.ALU._0994_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.ALU._1851_  (.A_N(\u_cpu.ALU._0838_ ),
    .B(\u_cpu.ALU.SrcA[19] ),
    .X(\u_cpu.ALU._0995_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1852_  (.A(\u_cpu.ALU._0838_ ),
    .B(\u_cpu.ALU._0837_ ),
    .X(\u_cpu.ALU._0996_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1853_  (.A1(\u_cpu.ALU._0641_ ),
    .A2(\u_cpu.ALU._0562_ ),
    .B1(\u_cpu.ALU._0843_ ),
    .C1(\u_cpu.ALU._0772_ ),
    .Y(\u_cpu.ALU._0997_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.ALU._1854_  (.A1(\u_cpu.ALU._0826_ ),
    .A2(\u_cpu.ALU._0995_ ),
    .A3(\u_cpu.ALU._0996_ ),
    .B1(\u_cpu.ALU._0997_ ),
    .Y(\u_cpu.ALU._0998_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1855_  (.A1(\u_cpu.ALU._0794_ ),
    .A2(\u_cpu.ALU._0580_ ),
    .B1(\u_cpu.ALU._0827_ ),
    .C1(\u_cpu.ALU._0772_ ),
    .Y(\u_cpu.ALU._0999_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.ALU._1856_  (.A1(\u_cpu.ALU._0726_ ),
    .A2(\u_cpu.ALU._0831_ ),
    .A3(\u_cpu.ALU._0832_ ),
    .B1(\u_cpu.ALU._0999_ ),
    .Y(\u_cpu.ALU._1000_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1857_  (.A0(\u_cpu.ALU._0993_ ),
    .A1(\u_cpu.ALU._0994_ ),
    .A2(\u_cpu.ALU._0998_ ),
    .A3(\u_cpu.ALU._1000_ ),
    .S0(\u_cpu.ALU._0805_ ),
    .S1(\u_cpu.ALU._0785_ ),
    .X(\u_cpu.ALU._1001_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU._1858_  (.A1(\u_cpu.ALU._0726_ ),
    .A2(\u_cpu.ALU._0995_ ),
    .A3(\u_cpu.ALU._0996_ ),
    .B1(\u_cpu.ALU._0997_ ),
    .X(\u_cpu.ALU._1002_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1859_  (.A(\u_cpu.ALU._0993_ ),
    .B(\u_cpu.ALU._0797_ ),
    .Y(\u_cpu.ALU._1003_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1860_  (.A1(\u_cpu.ALU._0797_ ),
    .A2(\u_cpu.ALU._1002_ ),
    .B1(\u_cpu.ALU._1003_ ),
    .C1(\u_cpu.ALU._0770_ ),
    .Y(\u_cpu.ALU._1004_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU._1861_  (.A1(\u_cpu.ALU._0722_ ),
    .A2(\u_cpu.ALU._0790_ ),
    .B1(\u_cpu.ALU._0797_ ),
    .B2(\u_cpu.ALU._1000_ ),
    .X(\u_cpu.ALU._1005_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1862_  (.A(\u_cpu.ALU._1004_ ),
    .B(\u_cpu.ALU._1005_ ),
    .Y(\u_cpu.ALU._1006_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1863_  (.A(\u_cpu.ALU._0900_ ),
    .B(\u_cpu.ALU._0757_ ),
    .Y(\u_cpu.ALU._1007_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU._1864_  (.A1_N(\u_cpu.ALU._0757_ ),
    .A2_N(\u_cpu.ALU._1001_ ),
    .B1(\u_cpu.ALU._1006_ ),
    .B2(\u_cpu.ALU._1007_ ),
    .Y(\u_cpu.ALU._1008_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1865_  (.A0(\u_cpu.ALU._0624_ ),
    .A1(\u_cpu.ALU._0618_ ),
    .A2(\u_cpu.ALU._0608_ ),
    .A3(\u_cpu.ALU.SrcA[6] ),
    .S0(\u_cpu.ALU._0635_ ),
    .S1(\u_cpu.ALU._0726_ ),
    .X(\u_cpu.ALU._1009_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1866_  (.A0(\u_cpu.ALU._0598_ ),
    .A1(\u_cpu.ALU._0663_ ),
    .A2(\u_cpu.ALU._0669_ ),
    .A3(\u_cpu.ALU._0666_ ),
    .S0(\u_cpu.ALU._0635_ ),
    .S1(\u_cpu.ALU._0772_ ),
    .X(\u_cpu.ALU._1010_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1867_  (.A0(\u_cpu.ALU._0686_ ),
    .A1(\u_cpu.ALU._0859_ ),
    .A2(\u_cpu.ALU.SrcA[13] ),
    .A3(\u_cpu.ALU._0679_ ),
    .S0(\u_cpu.ALU._0721_ ),
    .S1(\u_cpu.ALU._0772_ ),
    .X(\u_cpu.ALU._1011_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1868_  (.A0(\u_cpu.ALU._0948_ ),
    .A1(\u_cpu.ALU.SrcA[16] ),
    .A2(\u_cpu.ALU._0536_ ),
    .A3(\u_cpu.ALU.SrcA[18] ),
    .S0(\u_cpu.ALU._0721_ ),
    .S1(\u_cpu.ALU._0772_ ),
    .X(\u_cpu.ALU._1012_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1869_  (.A0(\u_cpu.ALU._1009_ ),
    .A1(\u_cpu.ALU._1010_ ),
    .A2(\u_cpu.ALU._1011_ ),
    .A3(\u_cpu.ALU._1012_ ),
    .S0(\u_cpu.ALU._0771_ ),
    .S1(\u_cpu.ALU._0760_ ),
    .X(\u_cpu.ALU._1013_ ));
 sky130_fd_sc_hd__nor3b_2 \u_cpu.ALU._1870_  (.A(\u_cpu.ALU._0752_ ),
    .B(\u_cpu.ALU._0750_ ),
    .C_N(\u_cpu.ALU._0751_ ),
    .Y(\u_cpu.ALU._1014_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1871_  (.A1(\u_cpu.ALU._0758_ ),
    .A2(\u_cpu.ALU._1013_ ),
    .B1(\u_cpu.ALU._1014_ ),
    .Y(\u_cpu.ALU._1015_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._1872_  (.A1(\u_cpu.ALU._0957_ ),
    .A2(\u_cpu.ALU._0624_ ),
    .B1(\u_cpu.ALU._0895_ ),
    .C1(\u_cpu.ALU._0805_ ),
    .X(\u_cpu.ALU._1016_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1873_  (.A0(\u_cpu.ALU._0624_ ),
    .A1(\u_cpu.ALU._0627_ ),
    .A2(\u_cpu.ALU._0632_ ),
    .A3(\u_cpu.ALU.SrcA[0] ),
    .S0(\u_cpu.ALU._0840_ ),
    .S1(\u_cpu.ALU._0638_ ),
    .X(\u_cpu.ALU._1017_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1874_  (.A(\u_cpu.ALU._0909_ ),
    .X(\u_cpu.ALU._1018_ ));
 sky130_fd_sc_hd__or4b_2 \u_cpu.ALU._1875_  (.A(_71951_),
    .B(\u_cpu.ALU._0745_ ),
    .C(\u_cpu.ALU._0735_ ),
    .D_N(_71952_),
    .X(\u_cpu.ALU._1019_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1876_  (.A(\u_cpu.ALU._1019_ ),
    .X(\u_cpu.ALU._1020_ ));
 sky130_fd_sc_hd__o32ai_2 \u_cpu.ALU._1877_  (.A1(\u_cpu.ALU._0811_ ),
    .A2(\u_cpu.ALU._0873_ ),
    .A3(\u_cpu.ALU._1018_ ),
    .B1(\u_cpu.ALU._0626_ ),
    .B2(\u_cpu.ALU._1020_ ),
    .Y(\u_cpu.ALU._1021_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU._1878_  (.A(\u_cpu.ALU._0623_ ),
    .B(\u_cpu.ALU._0624_ ),
    .X(\u_cpu.ALU._1022_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU._1879_  (.A1(\u_cpu.ALU._0960_ ),
    .A2(\u_cpu.ALU._0819_ ),
    .A3(\u_cpu.ALU._1017_ ),
    .B1(\u_cpu.ALU._1021_ ),
    .B2(\u_cpu.ALU._1022_ ),
    .X(\u_cpu.ALU._1023_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._1880_  (.A1(\u_cpu.ALU.Product_Wallace[3] ),
    .A2(\u_cpu.ALU._0821_ ),
    .B1(\u_cpu.ALU._1016_ ),
    .C1(\u_cpu.ALU._1023_ ),
    .X(\u_cpu.ALU._1024_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU._1881_  (.A1(\u_cpu.ALU._1008_ ),
    .A2(\u_cpu.ALU._1015_ ),
    .B1_N(\u_cpu.ALU._1024_ ),
    .Y(\u_cpu.ALU._1025_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU._1882_  (.A1(\u_cpu.ALU._0975_ ),
    .A2(\u_cpu.ALU._0984_ ),
    .A3(\u_cpu.ALU._0991_ ),
    .B1(\u_cpu.ALU._1025_ ),
    .Y(\u_cpu.ALU._1026_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1883_  (.A(\u_cpu.ALU._1026_ ),
    .Y(\u_cpu.ALU.ALUResult[3] ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU._1884_  (.A1(\u_cpu.ALU._0978_ ),
    .A2(\u_cpu.ALU._0979_ ),
    .B1(\u_cpu.ALU._0981_ ),
    .B2(\u_cpu.ALU._0989_ ),
    .Y(\u_cpu.ALU._1027_ ));
 sky130_fd_sc_hd__a41oi_2 \u_cpu.ALU._1885_  (.A1(\u_cpu.ALU._0917_ ),
    .A2(\u_cpu.ALU._0908_ ),
    .A3(\u_cpu.ALU._0989_ ),
    .A4(\u_cpu.ALU._0990_ ),
    .B1(\u_cpu.ALU._1027_ ),
    .Y(\u_cpu.ALU._1028_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1886_  (.A1(\u_cpu.ALU._0801_ ),
    .A2(\u_cpu.ALU._0914_ ),
    .B1(\u_cpu.ALU._0613_ ),
    .Y(\u_cpu.ALU._1029_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._1887_  (.A1(\u_cpu.ALU._0911_ ),
    .A2(\u_cpu.ALU._0960_ ),
    .B1(\u_cpu.ALU._0814_ ),
    .B2(\u_cpu.ALU._0745_ ),
    .C1(\u_cpu.ALU._0613_ ),
    .X(\u_cpu.ALU._1030_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._1888_  (.A1(\u_cpu.ALU._1029_ ),
    .A2(\u_cpu.ALU._1030_ ),
    .B1(\u_cpu.ALU._0618_ ),
    .X(\u_cpu.ALU._1031_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._1889_  (.A(\u_cpu.ALU._1030_ ),
    .B(\u_cpu.ALU._0618_ ),
    .C(\u_cpu.ALU._1029_ ),
    .Y(\u_cpu.ALU._1032_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1890_  (.A(\u_cpu.ALU._1031_ ),
    .B(\u_cpu.ALU._1032_ ),
    .Y(\u_cpu.ALU._1033_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1891_  (.A(\u_cpu.ALU._1028_ ),
    .B(\u_cpu.ALU._1033_ ),
    .Y(\u_cpu.ALU._1034_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._1892_  (.A(\u_cpu.ALU._0849_ ),
    .B(\u_cpu.ALU._0982_ ),
    .C(\u_cpu.ALU._0979_ ),
    .X(\u_cpu.ALU._1035_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1893_  (.A(\u_cpu.ALU._0916_ ),
    .B(\u_cpu.ALU._0983_ ),
    .Y(\u_cpu.ALU._1036_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU._1894_  (.A(\u_cpu.ALU._0917_ ),
    .B(\u_cpu.ALU._0908_ ),
    .C(\u_cpu.ALU._0989_ ),
    .D(\u_cpu.ALU._0990_ ),
    .Y(\u_cpu.ALU._1037_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1895_  (.A1(\u_cpu.ALU._1035_ ),
    .A2(\u_cpu.ALU._1036_ ),
    .B1(\u_cpu.ALU._1037_ ),
    .Y(\u_cpu.ALU._1038_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._1896_  (.A(\u_cpu.ALU._1031_ ),
    .B(\u_cpu.ALU._1032_ ),
    .C(\u_cpu.ALU._1038_ ),
    .Y(\u_cpu.ALU._1039_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU._1897_  (.A1(\u_cpu.ALU._0826_ ),
    .A2(\u_cpu.ALU._0792_ ),
    .A3(\u_cpu.ALU._0793_ ),
    .B1(\u_cpu.ALU._0796_ ),
    .C1(\u_cpu.ALU._0768_ ),
    .X(\u_cpu.ALU._1040_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1898_  (.A1(\u_cpu.ALU._0958_ ),
    .A2(\u_cpu.ALU._0803_ ),
    .B1(\u_cpu.ALU._1040_ ),
    .Y(\u_cpu.ALU._1041_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1899_  (.A1(\u_cpu.ALU._0729_ ),
    .A2(\u_cpu.ALU._0774_ ),
    .B1(\u_cpu.ALU._0771_ ),
    .C1(\u_cpu.ALU._0778_ ),
    .Y(\u_cpu.ALU._1042_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1900_  (.A1(\u_cpu.ALU._0958_ ),
    .A2(\u_cpu.ALU._0802_ ),
    .B1(\u_cpu.ALU._1042_ ),
    .C1(\u_cpu.ALU._0760_ ),
    .Y(\u_cpu.ALU._1043_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1901_  (.A1(\u_cpu.ALU._0806_ ),
    .A2(\u_cpu.ALU._1041_ ),
    .B1(\u_cpu.ALU._1043_ ),
    .Y(\u_cpu.ALU._1044_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1902_  (.A0(\u_cpu.ALU._0618_ ),
    .A1(\u_cpu.ALU._0624_ ),
    .A2(\u_cpu.ALU._0627_ ),
    .A3(\u_cpu.ALU.SrcA[1] ),
    .S0(\u_cpu.ALU._0775_ ),
    .S1(\u_cpu.ALU._0725_ ),
    .X(\u_cpu.ALU._1045_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._1903_  (.A1(\u_cpu.ALU._0641_ ),
    .A2(\u_cpu.ALU._0787_ ),
    .A3(\u_cpu.ALU.SrcA[0] ),
    .B1(\u_cpu.ALU._0768_ ),
    .X(\u_cpu.ALU._1046_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU._1904_  (.A(\u_cpu.ALU._0647_ ),
    .B(\u_cpu.ALU._0737_ ),
    .C(\u_cpu.ALU._0752_ ),
    .D(\u_cpu.ALU._0881_ ),
    .X(\u_cpu.ALU._1047_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._1905_  (.A1(\u_cpu.ALU._0958_ ),
    .A2(\u_cpu.ALU._1045_ ),
    .B1(\u_cpu.ALU._1046_ ),
    .C1(\u_cpu.ALU._1047_ ),
    .X(\u_cpu.ALU._1048_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1906_  (.A1(\u_cpu.ALU._1044_ ),
    .A2(\u_cpu.ALU._1014_ ),
    .B1(\u_cpu.ALU._1048_ ),
    .Y(\u_cpu.ALU._1049_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._1907_  (.A1(\u_cpu.ALU._0613_ ),
    .A2(\u_cpu.ALU._0618_ ),
    .B1(\u_cpu.ALU._0742_ ),
    .C1(\u_cpu.ALU._0746_ ),
    .D1(\u_cpu.ALU._0752_ ),
    .X(\u_cpu.ALU._1050_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._1908_  (.A1(\u_cpu.ALU._0620_ ),
    .A2(\u_cpu.ALU._0743_ ),
    .B1(\u_cpu.ALU._0820_ ),
    .B2(\u_cpu.ALU.Product_Wallace[4] ),
    .C1(\u_cpu.ALU._1050_ ),
    .X(\u_cpu.ALU._1051_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1909_  (.A1(\u_cpu.ALU._0757_ ),
    .A2(\u_cpu.ALU._0753_ ),
    .B1(\u_cpu.ALU._1051_ ),
    .Y(\u_cpu.ALU._1052_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU._1910_  (.A1(\u_cpu.ALU._0619_ ),
    .A2(\u_cpu.ALU._0620_ ),
    .A3(\u_cpu.ALU._1020_ ),
    .B1(\u_cpu.ALU._1052_ ),
    .X(\u_cpu.ALU._1053_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._1911_  (.A1(\u_cpu.ALU._0923_ ),
    .A2(\u_cpu.ALU._0924_ ),
    .B1(\u_cpu.ALU._0728_ ),
    .X(\u_cpu.ALU._1054_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._1912_  (.A1(\u_cpu.ALU._0787_ ),
    .A2(\u_cpu.ALU._0933_ ),
    .B1(\u_cpu.ALU._0765_ ),
    .C1(\u_cpu.ALU._1054_ ),
    .X(\u_cpu.ALU._1055_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1913_  (.A1(\u_cpu.ALU._0958_ ),
    .A2(\u_cpu.ALU._0767_ ),
    .B1(\u_cpu.ALU._1055_ ),
    .C1(\u_cpu.ALU._0770_ ),
    .Y(\u_cpu.ALU._1056_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1914_  (.A(\u_cpu.ALU._0629_ ),
    .B(\u_cpu.ALU._0647_ ),
    .Y(\u_cpu.ALU._1057_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.ALU._1915_  (.A(\u_cpu.ALU._0647_ ),
    .B(\u_cpu.ALU._0765_ ),
    .C(\u_cpu.ALU._0994_ ),
    .X(\u_cpu.ALU._1058_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU._1916_  (.A1_N(\u_cpu.ALU._0762_ ),
    .A2_N(\u_cpu.ALU._1057_ ),
    .B1(\u_cpu.ALU._1058_ ),
    .B2(\u_cpu.ALU._0900_ ),
    .X(\u_cpu.ALU._1059_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._1917_  (.A1(\u_cpu.ALU._1056_ ),
    .A2(\u_cpu.ALU._1059_ ),
    .B1(\u_cpu.ALU._0817_ ),
    .C1(\u_cpu.ALU._0784_ ),
    .X(\u_cpu.ALU._1060_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1918_  (.A1(\u_cpu.ALU._0758_ ),
    .A2(\u_cpu.ALU._1049_ ),
    .B1(\u_cpu.ALU._1053_ ),
    .C1(\u_cpu.ALU._1060_ ),
    .Y(\u_cpu.ALU._1061_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU._1919_  (.A1(\u_cpu.ALU._0975_ ),
    .A2(\u_cpu.ALU._1034_ ),
    .A3(\u_cpu.ALU._1039_ ),
    .B1(\u_cpu.ALU._1061_ ),
    .Y(\u_cpu.ALU._1062_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._1920_  (.A(\u_cpu.ALU._1062_ ),
    .Y(\u_cpu.ALU.ALUResult[4] ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1921_  (.A(\u_cpu.ALU.SrcB[4] ),
    .B(\u_cpu.ALU.SrcB[3] ),
    .Y(\u_cpu.ALU._1063_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._1922_  (.A(\u_cpu.ALU._0911_ ),
    .B(\u_cpu.ALU._1063_ ),
    .C(\u_cpu.ALU._0764_ ),
    .Y(\u_cpu.ALU._1064_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU._1923_  (.A1(_71953_),
    .A2(\u_cpu.ALU._0735_ ),
    .A3(\u_cpu.ALU._0708_ ),
    .B1(\u_cpu.ALU._1064_ ),
    .X(\u_cpu.ALU._1065_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU._1924_  (.A1(\u_cpu.ALU._0609_ ),
    .A2(\u_cpu.ALU._1065_ ),
    .B1_N(\u_cpu.ALU.SrcA[5] ),
    .Y(\u_cpu.ALU._1066_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU._1925_  (.A1(_71954_),
    .A2(\u_cpu.ALU._0735_ ),
    .A3(\u_cpu.ALU._0708_ ),
    .B1(\u_cpu.ALU._1064_ ),
    .C1(\u_cpu.ALU._0609_ ),
    .X(\u_cpu.ALU._1067_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1926_  (.A1(\u_cpu.ALU._0985_ ),
    .A2(\u_cpu.ALU._1064_ ),
    .B1(\u_cpu.ALU._0609_ ),
    .Y(\u_cpu.ALU._1068_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1927_  (.A1(\u_cpu.ALU._1068_ ),
    .A2(\u_cpu.ALU._1067_ ),
    .B1(\u_cpu.ALU._0608_ ),
    .Y(\u_cpu.ALU._1069_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1928_  (.A1(\u_cpu.ALU._1033_ ),
    .A2(\u_cpu.ALU._1028_ ),
    .B1(\u_cpu.ALU._1032_ ),
    .Y(\u_cpu.ALU._1070_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1929_  (.A1(\u_cpu.ALU._1066_ ),
    .A2(\u_cpu.ALU._1067_ ),
    .B1(\u_cpu.ALU._1069_ ),
    .C1(\u_cpu.ALU._1070_ ),
    .Y(\u_cpu.ALU._1071_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1930_  (.A1(\u_cpu.ALU._1067_ ),
    .A2(\u_cpu.ALU._1066_ ),
    .B1(\u_cpu.ALU._1069_ ),
    .Y(\u_cpu.ALU._1072_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1931_  (.A1(\u_cpu.ALU._1033_ ),
    .A2(\u_cpu.ALU._1028_ ),
    .B1(\u_cpu.ALU._1072_ ),
    .C1(\u_cpu.ALU._1032_ ),
    .Y(\u_cpu.ALU._1073_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._1932_  (.A(\u_cpu.ALU._1071_ ),
    .B(\u_cpu.ALU._1073_ ),
    .C(\u_cpu.ALU._0814_ ),
    .Y(\u_cpu.ALU._1074_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1933_  (.A(\u_cpu.ALU._0879_ ),
    .X(\u_cpu.ALU._1075_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1934_  (.A(\u_cpu.ALU._0770_ ),
    .X(\u_cpu.ALU._1076_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._1935_  (.A(\u_cpu.ALU._0963_ ),
    .B(\u_cpu.ALU._0881_ ),
    .C(\u_cpu.ALU._0737_ ),
    .X(\u_cpu.ALU._1077_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1936_  (.A0(\u_cpu.ALU._0608_ ),
    .A1(\u_cpu.ALU._0618_ ),
    .A2(\u_cpu.ALU._0624_ ),
    .A3(\u_cpu.ALU._0627_ ),
    .S0(\u_cpu.ALU._0838_ ),
    .S1(\u_cpu.ALU._0728_ ),
    .X(\u_cpu.ALU._1078_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.ALU._1937_  (.A0(\u_cpu.ALU._1078_ ),
    .A1(\u_cpu.ALU._0893_ ),
    .S(\u_cpu.ALU._0771_ ),
    .X(\u_cpu.ALU._1079_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1938_  (.A(\u_cpu.ALU._0861_ ),
    .B(\u_cpu.ALU._0864_ ),
    .Y(\u_cpu.ALU._1080_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU._1939_  (.A1(\u_cpu.ALU._0726_ ),
    .A2(\u_cpu.ALU._0865_ ),
    .A3(\u_cpu.ALU._0866_ ),
    .B1(\u_cpu.ALU._0868_ ),
    .X(\u_cpu.ALU._1081_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1940_  (.A0(\u_cpu.ALU._1080_ ),
    .A1(\u_cpu.ALU._0856_ ),
    .A2(\u_cpu.ALU._0839_ ),
    .A3(\u_cpu.ALU._1081_ ),
    .S0(\u_cpu.ALU._0768_ ),
    .S1(\u_cpu.ALU._0760_ ),
    .X(\u_cpu.ALU._1082_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU._1941_  (.A1(\u_cpu.ALU._1076_ ),
    .A2(\u_cpu.ALU._1077_ ),
    .A3(\u_cpu.ALU._1079_ ),
    .B1(\u_cpu.ALU._1082_ ),
    .B2(\u_cpu.ALU._1014_ ),
    .X(\u_cpu.ALU._1083_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1942_  (.A(\u_cpu.ALU._1075_ ),
    .B(\u_cpu.ALU._1083_ ),
    .Y(\u_cpu.ALU._1084_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._1943_  (.A1(\u_cpu.ALU._0772_ ),
    .A2(\u_cpu.ALU._0842_ ),
    .B1(\u_cpu.ALU._0845_ ),
    .X(\u_cpu.ALU._1085_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU._1944_  (.A1(\u_cpu.ALU._0643_ ),
    .A2(\u_cpu.ALU._0831_ ),
    .A3(\u_cpu.ALU._0832_ ),
    .B1(\u_cpu.ALU._0834_ ),
    .X(\u_cpu.ALU._1086_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1945_  (.A0(\u_cpu.ALU._1085_ ),
    .A1(\u_cpu.ALU._1086_ ),
    .A2(\u_cpu.ALU._0830_ ),
    .A3(\u_cpu.ALU.SrcA[31] ),
    .S0(\u_cpu.ALU._0771_ ),
    .S1(\u_cpu.ALU._0805_ ),
    .X(\u_cpu.ALU._1087_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._1946_  (.A(\u_cpu.ALU._0647_ ),
    .X(\u_cpu.ALU._1088_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.ALU._1947_  (.A0(\u_cpu.ALU._1085_ ),
    .A1(\u_cpu.ALU._1086_ ),
    .S(\u_cpu.ALU._0771_ ),
    .X(\u_cpu.ALU._1089_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1948_  (.A(\u_cpu.ALU._0765_ ),
    .B(\u_cpu.ALU._0623_ ),
    .Y(\u_cpu.ALU._1090_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU._1949_  (.A1_N(\u_cpu.ALU._1088_ ),
    .A2_N(\u_cpu.ALU._1089_ ),
    .B1(\u_cpu.ALU._0876_ ),
    .B2(\u_cpu.ALU._1090_ ),
    .Y(\u_cpu.ALU._1091_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU._1950_  (.A1(\u_cpu.ALU._0874_ ),
    .A2(\u_cpu.ALU._1087_ ),
    .B1(\u_cpu.ALU._1091_ ),
    .B2(\u_cpu.ALU._0882_ ),
    .X(\u_cpu.ALU._1092_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._1951_  (.A(\u_cpu.ALU._0608_ ),
    .B(\u_cpu.ALU._0609_ ),
    .C(\u_cpu.ALU._0744_ ),
    .X(\u_cpu.ALU._1093_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1952_  (.A(\u_cpu.ALU._0611_ ),
    .B(\u_cpu.ALU._0612_ ),
    .Y(\u_cpu.ALU._1094_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._1953_  (.A1(\u_cpu.ALU._0608_ ),
    .A2(\u_cpu.ALU._0609_ ),
    .B1(\u_cpu.ALU._0742_ ),
    .C1(\u_cpu.ALU._0881_ ),
    .D1(\u_cpu.ALU._0752_ ),
    .X(\u_cpu.ALU._1095_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._1954_  (.A1(\u_cpu.ALU._0609_ ),
    .A2(\u_cpu.ALU._0753_ ),
    .B1(\u_cpu.ALU._0812_ ),
    .B2(\u_cpu.ALU._1094_ ),
    .C1(\u_cpu.ALU._1095_ ),
    .X(\u_cpu.ALU._1096_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._1955_  (.A1(\u_cpu.ALU.Product_Wallace[5] ),
    .A2(\u_cpu.ALU._0821_ ),
    .B1(\u_cpu.ALU._1093_ ),
    .C1(\u_cpu.ALU._1096_ ),
    .X(\u_cpu.ALU._1097_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1956_  (.A1(\u_cpu.ALU._1092_ ),
    .A2(\u_cpu.ALU._0759_ ),
    .B1(\u_cpu.ALU._1097_ ),
    .Y(\u_cpu.ALU._1098_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._1957_  (.A(\u_cpu.ALU._1074_ ),
    .B(\u_cpu.ALU._1084_ ),
    .C(\u_cpu.ALU._1098_ ),
    .Y(\u_cpu.ALU.ALUResult[5] ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1958_  (.A(\u_cpu.ALU.SrcB[4] ),
    .B(\u_cpu.ALU.SrcB[5] ),
    .Y(\u_cpu.ALU._1099_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU._1959_  (.A(\u_cpu.ALU._0960_ ),
    .B(\u_cpu.ALU._1099_ ),
    .C(\u_cpu.ALU._0640_ ),
    .D(\u_cpu.ALU._0642_ ),
    .Y(\u_cpu.ALU._1100_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._1960_  (.A1(\u_cpu.ALU._0985_ ),
    .A2(\u_cpu.ALU._1100_ ),
    .B1(\u_cpu.ALU.SrcB[6] ),
    .X(\u_cpu.ALU._1101_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1961_  (.A1(\u_cpu.ALU._0708_ ),
    .A2(\u_cpu.ALU._1018_ ),
    .B1(\u_cpu.ALU._1100_ ),
    .C1(\u_cpu.ALU.SrcB[6] ),
    .Y(\u_cpu.ALU._1102_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._1962_  (.A1(\u_cpu.ALU._1101_ ),
    .A2(\u_cpu.ALU._1102_ ),
    .B1(\u_cpu.ALU._0606_ ),
    .X(\u_cpu.ALU._1103_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._1963_  (.A(\u_cpu.ALU._0606_ ),
    .B(\u_cpu.ALU._1101_ ),
    .C(\u_cpu.ALU._1102_ ),
    .Y(\u_cpu.ALU._1104_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1964_  (.A(\u_cpu.ALU._1103_ ),
    .B(\u_cpu.ALU._1104_ ),
    .X(\u_cpu.ALU._1105_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1965_  (.A1(\u_cpu.ALU._0609_ ),
    .A2(\u_cpu.ALU._1065_ ),
    .B1(\u_cpu.ALU._1066_ ),
    .Y(\u_cpu.ALU._1106_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._1966_  (.A(\u_cpu.ALU._1032_ ),
    .B(\u_cpu.ALU._1069_ ),
    .X(\u_cpu.ALU._1107_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU._1967_  (.A1(\u_cpu.ALU._1067_ ),
    .A2(\u_cpu.ALU._1066_ ),
    .B1(\u_cpu.ALU._1069_ ),
    .C1(\u_cpu.ALU._1031_ ),
    .D1(\u_cpu.ALU._1032_ ),
    .Y(\u_cpu.ALU._1108_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU._1968_  (.A1(\u_cpu.ALU._1106_ ),
    .A2(\u_cpu.ALU._1107_ ),
    .B1(\u_cpu.ALU._1108_ ),
    .B2(\u_cpu.ALU._1028_ ),
    .Y(\u_cpu.ALU._1109_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1969_  (.A1(\u_cpu.ALU._1109_ ),
    .A2(\u_cpu.ALU._1105_ ),
    .B1(\u_cpu.ALU._0921_ ),
    .Y(\u_cpu.ALU._1110_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1970_  (.A1(\u_cpu.ALU._1105_ ),
    .A2(\u_cpu.ALU._1109_ ),
    .B1(\u_cpu.ALU._1110_ ),
    .Y(\u_cpu.ALU._1111_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1971_  (.A(\u_cpu.ALU._0775_ ),
    .B(\u_cpu.ALU.SrcA[5] ),
    .Y(\u_cpu.ALU._1112_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._1972_  (.A1(\u_cpu.ALU._0838_ ),
    .A2(\u_cpu.ALU._0606_ ),
    .B1(\u_cpu.ALU._1112_ ),
    .C1(\u_cpu.ALU._0643_ ),
    .Y(\u_cpu.ALU._1113_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU._1973_  (.A1(\u_cpu.ALU._0787_ ),
    .A2(\u_cpu.ALU._0788_ ),
    .A3(\u_cpu.ALU._0793_ ),
    .B1(\u_cpu.ALU._1113_ ),
    .X(\u_cpu.ALU._1114_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.ALU._1974_  (.A0(\u_cpu.ALU._0962_ ),
    .A1(\u_cpu.ALU._1114_ ),
    .S(\u_cpu.ALU._0785_ ),
    .X(\u_cpu.ALU._1115_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU._1975_  (.A1(\u_cpu.ALU._0787_ ),
    .A2(\u_cpu.ALU._0937_ ),
    .A3(\u_cpu.ALU._0938_ ),
    .B1(\u_cpu.ALU._0939_ ),
    .X(\u_cpu.ALU._1116_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._1976_  (.A0(\u_cpu.ALU._1116_ ),
    .A1(\u_cpu.ALU._0951_ ),
    .A2(\u_cpu.ALU._0949_ ),
    .A3(\u_cpu.ALU._0945_ ),
    .S0(\u_cpu.ALU._0647_ ),
    .S1(\u_cpu.ALU._0769_ ),
    .X(\u_cpu.ALU._1117_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU._1977_  (.A1(\u_cpu.ALU._1076_ ),
    .A2(\u_cpu.ALU._1077_ ),
    .A3(\u_cpu.ALU._1115_ ),
    .B1(\u_cpu.ALU._1117_ ),
    .B2(\u_cpu.ALU._1014_ ),
    .X(\u_cpu.ALU._1118_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1978_  (.A(\u_cpu.ALU._1075_ ),
    .B(\u_cpu.ALU._1118_ ),
    .Y(\u_cpu.ALU._1119_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._1979_  (.A1(\u_cpu.ALU._0643_ ),
    .A2(\u_cpu.ALU._0933_ ),
    .B1(\u_cpu.ALU._0935_ ),
    .X(\u_cpu.ALU._1120_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU._1980_  (.A1(\u_cpu.ALU._0725_ ),
    .A2(\u_cpu.ALU._0923_ ),
    .A3(\u_cpu.ALU._0924_ ),
    .B1(\u_cpu.ALU._0927_ ),
    .C1(\u_cpu.ALU._0629_ ),
    .X(\u_cpu.ALU._1121_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1981_  (.A1(\u_cpu.ALU._1120_ ),
    .A2(\u_cpu.ALU._0765_ ),
    .B1(\u_cpu.ALU._1121_ ),
    .Y(\u_cpu.ALU._1122_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.ALU._1982_  (.A1(\u_cpu.ALU._0790_ ),
    .A2(\u_cpu.ALU._0930_ ),
    .A3(\u_cpu.ALU._1090_ ),
    .B1(\u_cpu.ALU._0805_ ),
    .B2(\u_cpu.ALU._1122_ ),
    .X(\u_cpu.ALU._1123_ ));
 sky130_fd_sc_hd__or4b_2 \u_cpu.ALU._1983_  (.A(\u_cpu.ALU._0752_ ),
    .B(\u_cpu.ALU._0881_ ),
    .C(\u_cpu.ALU._0750_ ),
    .D_N(\u_cpu.ALU._0751_ ),
    .X(\u_cpu.ALU._1124_ ));
 sky130_fd_sc_hd__or4b_2 \u_cpu.ALU._1984_  (.A(\u_cpu.ALU._0752_ ),
    .B(\u_cpu.ALU._0873_ ),
    .C(\u_cpu.ALU._0750_ ),
    .D_N(\u_cpu.ALU._0751_ ),
    .X(\u_cpu.ALU._1125_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU._1985_  (.A1(\u_cpu.ALU._1090_ ),
    .A2(\u_cpu.ALU._0967_ ),
    .B1(\u_cpu.ALU._0805_ ),
    .B2(\u_cpu.ALU._1122_ ),
    .C1(\u_cpu.ALU._1058_ ),
    .X(\u_cpu.ALU._1126_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU._1986_  (.A1(\u_cpu.ALU._1123_ ),
    .A2(\u_cpu.ALU._1124_ ),
    .B1(\u_cpu.ALU._1125_ ),
    .B2(\u_cpu.ALU._1126_ ),
    .X(\u_cpu.ALU._1127_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._1987_  (.A(\u_cpu.ALU._0605_ ),
    .B(\u_cpu.ALU._0607_ ),
    .Y(\u_cpu.ALU._1128_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._1988_  (.A1(\u_cpu.ALU.SrcA[6] ),
    .A2(\u_cpu.ALU.SrcB[6] ),
    .B1(\u_cpu.ALU._0742_ ),
    .C1(\u_cpu.ALU._0746_ ),
    .D1(\u_cpu.ALU._0752_ ),
    .X(\u_cpu.ALU._1129_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._1989_  (.A1(\u_cpu.ALU._0607_ ),
    .A2(\u_cpu.ALU._0743_ ),
    .B1(\u_cpu.ALU._0820_ ),
    .B2(\u_cpu.ALU.Product_Wallace[6] ),
    .C1(\u_cpu.ALU._1129_ ),
    .X(\u_cpu.ALU._1130_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._1990_  (.A1(\u_cpu.ALU.SrcB[6] ),
    .A2(\u_cpu.ALU._0754_ ),
    .B1(\u_cpu.ALU._0812_ ),
    .B2(\u_cpu.ALU._1128_ ),
    .C1(\u_cpu.ALU._1130_ ),
    .X(\u_cpu.ALU._1131_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.ALU._1991_  (.A1(\u_cpu.ALU._0879_ ),
    .A2(\u_cpu.ALU._1127_ ),
    .B1_N(\u_cpu.ALU._1131_ ),
    .X(\u_cpu.ALU._1132_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._1992_  (.A(\u_cpu.ALU._1111_ ),
    .B(\u_cpu.ALU._1119_ ),
    .C(\u_cpu.ALU._1132_ ),
    .Y(\u_cpu.ALU.ALUResult[6] ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._1993_  (.A(\u_cpu.ALU._1109_ ),
    .B(\u_cpu.ALU._1105_ ),
    .Y(\u_cpu.ALU._1133_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU._1994_  (.A(\u_cpu.ALU._0911_ ),
    .B(\u_cpu.ALU._0960_ ),
    .C(\u_cpu.ALU._1099_ ),
    .D(\u_cpu.ALU._0604_ ),
    .Y(\u_cpu.ALU._1134_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._1995_  (.A1(\u_cpu.ALU._0985_ ),
    .A2(\u_cpu.ALU._1134_ ),
    .B1(\u_cpu.ALU.SrcB[7] ),
    .Y(\u_cpu.ALU._1135_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU._1996_  (.A1(_71955_),
    .A2(\u_cpu.ALU._0709_ ),
    .A3(\u_cpu.ALU._0909_ ),
    .B1(\u_cpu.ALU._1134_ ),
    .C1(\u_cpu.ALU.SrcB[7] ),
    .X(\u_cpu.ALU._1136_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._1997_  (.A1(\u_cpu.ALU._1135_ ),
    .A2(\u_cpu.ALU._1136_ ),
    .B1(\u_cpu.ALU._0598_ ),
    .Y(\u_cpu.ALU._1137_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._1998_  (.A1(\u_cpu.ALU._0985_ ),
    .A2(\u_cpu.ALU._1134_ ),
    .B1(\u_cpu.ALU.SrcB[7] ),
    .X(\u_cpu.ALU._1138_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU._1999_  (.A1(\u_cpu.ALU._0710_ ),
    .A2(\u_cpu.ALU._0919_ ),
    .B1(\u_cpu.ALU.SrcB[6] ),
    .B2(\u_cpu.ALU._1100_ ),
    .C1(\u_cpu.ALU.SrcB[7] ),
    .Y(\u_cpu.ALU._1139_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU._2000_  (.A_N(\u_cpu.ALU.SrcA[7] ),
    .B(\u_cpu.ALU._1138_ ),
    .C(\u_cpu.ALU._1139_ ),
    .Y(\u_cpu.ALU._1140_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2001_  (.A(\u_cpu.ALU._1137_ ),
    .B(\u_cpu.ALU._1140_ ),
    .Y(\u_cpu.ALU._1141_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2002_  (.A1(\u_cpu.ALU._1103_ ),
    .A2(\u_cpu.ALU._1133_ ),
    .B1(\u_cpu.ALU._1141_ ),
    .X(\u_cpu.ALU._1142_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._2003_  (.A(\u_cpu.ALU._1103_ ),
    .B(\u_cpu.ALU._1133_ ),
    .C(\u_cpu.ALU._1141_ ),
    .Y(\u_cpu.ALU._1143_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2004_  (.A(\u_cpu.ALU._0758_ ),
    .X(\u_cpu.ALU._1144_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2005_  (.A(\u_cpu.ALU._0958_ ),
    .X(\u_cpu.ALU._1145_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2006_  (.A1(\u_cpu.ALU._0790_ ),
    .A2(\u_cpu.ALU._0842_ ),
    .B1(\u_cpu.ALU._0992_ ),
    .X(\u_cpu.ALU._1146_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2007_  (.A(\u_cpu.ALU._0958_ ),
    .B(\u_cpu.ALU._1146_ ),
    .Y(\u_cpu.ALU._1147_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._2008_  (.A1(\u_cpu.ALU._1000_ ),
    .A2(\u_cpu.ALU._1145_ ),
    .B1(\u_cpu.ALU._0806_ ),
    .C1(\u_cpu.ALU._1147_ ),
    .X(\u_cpu.ALU._1148_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2009_  (.A(\u_cpu.ALU._0900_ ),
    .X(\u_cpu.ALU._1149_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._2010_  (.A1(\u_cpu.ALU._1149_ ),
    .A2(\u_cpu.ALU._0986_ ),
    .B1(\u_cpu.ALU._0994_ ),
    .C1(\u_cpu.ALU._1076_ ),
    .X(\u_cpu.ALU._1150_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2011_  (.A1(\u_cpu.ALU._1148_ ),
    .A2(\u_cpu.ALU._1150_ ),
    .B1(\u_cpu.ALU._0784_ ),
    .Y(\u_cpu.ALU._1151_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2012_  (.A(\u_cpu.ALU._1020_ ),
    .B(\u_cpu.ALU._0603_ ),
    .Y(\u_cpu.ALU._1152_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2013_  (.A1(\u_cpu.ALU._0602_ ),
    .A2(\u_cpu.ALU._0748_ ),
    .B1(\u_cpu.ALU._0820_ ),
    .B2(\u_cpu.ALU.Product_Wallace[7] ),
    .C1(\u_cpu.ALU._1152_ ),
    .X(\u_cpu.ALU._1153_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2014_  (.A1(\u_cpu.ALU._0601_ ),
    .A2(\u_cpu.ALU._0744_ ),
    .B1(\u_cpu.ALU._0754_ ),
    .B2(\u_cpu.ALU.SrcB[7] ),
    .C1(\u_cpu.ALU._1153_ ),
    .X(\u_cpu.ALU._1154_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2015_  (.A0(\u_cpu.ALU._0598_ ),
    .A1(\u_cpu.ALU.SrcA[6] ),
    .A2(\u_cpu.ALU._0608_ ),
    .A3(\u_cpu.ALU._0618_ ),
    .S0(\u_cpu.ALU._0794_ ),
    .S1(\u_cpu.ALU._0729_ ),
    .X(\u_cpu.ALU._1155_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.ALU._2016_  (.A0(\u_cpu.ALU._1017_ ),
    .A1(\u_cpu.ALU._1155_ ),
    .S(\u_cpu.ALU._0769_ ),
    .X(\u_cpu.ALU._1156_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2017_  (.A0(\u_cpu.ALU._1002_ ),
    .A1(\u_cpu.ALU._1012_ ),
    .A2(\u_cpu.ALU._1011_ ),
    .A3(\u_cpu.ALU._1010_ ),
    .S0(\u_cpu.ALU._0785_ ),
    .S1(\u_cpu.ALU._1088_ ),
    .X(\u_cpu.ALU._1157_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2018_  (.A(\u_cpu.ALU._1014_ ),
    .X(\u_cpu.ALU._1158_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU._2019_  (.A1(\u_cpu.ALU._1047_ ),
    .A2(\u_cpu.ALU._1156_ ),
    .B1(\u_cpu.ALU._1157_ ),
    .B2(\u_cpu.ALU._1158_ ),
    .Y(\u_cpu.ALU._1159_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2020_  (.A(\u_cpu.ALU._0759_ ),
    .B(\u_cpu.ALU._1159_ ),
    .Y(\u_cpu.ALU._1160_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._2021_  (.A1(\u_cpu.ALU._1144_ ),
    .A2(\u_cpu.ALU._1151_ ),
    .B1(\u_cpu.ALU._1154_ ),
    .C1(\u_cpu.ALU._1160_ ),
    .X(\u_cpu.ALU._1161_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU._2022_  (.A1(\u_cpu.ALU._1142_ ),
    .A2(\u_cpu.ALU._1143_ ),
    .A3(\u_cpu.ALU._0975_ ),
    .B1(\u_cpu.ALU._1161_ ),
    .Y(\u_cpu.ALU._1162_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._2023_  (.A(\u_cpu.ALU._1162_ ),
    .Y(\u_cpu.ALU.ALUResult[7] ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._2024_  (.A(\u_cpu.ALU._0664_ ),
    .Y(\u_cpu.ALU._1163_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._2025_  (.A(\u_cpu.ALU._1099_ ),
    .B(\u_cpu.ALU._0604_ ),
    .C(\u_cpu.ALU._0599_ ),
    .Y(\u_cpu.ALU._1164_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2026_  (.A(\u_cpu.ALU._0911_ ),
    .B(\u_cpu.ALU._0960_ ),
    .Y(\u_cpu.ALU._1165_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU._2027_  (.A1(\u_cpu.ALU._0709_ ),
    .A2(\u_cpu.ALU._0919_ ),
    .B1(\u_cpu.ALU._1164_ ),
    .B2(\u_cpu.ALU._1165_ ),
    .Y(\u_cpu.ALU._1166_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2028_  (.A(\u_cpu.ALU._1163_ ),
    .B(\u_cpu.ALU._1166_ ),
    .Y(\u_cpu.ALU._1167_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU._2029_  (.A1(\u_cpu.ALU._0710_ ),
    .A2(\u_cpu.ALU._0919_ ),
    .B1(\u_cpu.ALU._1164_ ),
    .B2(\u_cpu.ALU._1165_ ),
    .C1(\u_cpu.ALU._0664_ ),
    .Y(\u_cpu.ALU._1168_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._2030_  (.A(\u_cpu.ALU._0693_ ),
    .B(\u_cpu.ALU._1167_ ),
    .C(\u_cpu.ALU._1168_ ),
    .Y(\u_cpu.ALU._1169_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2031_  (.A1(\u_cpu.ALU._1166_ ),
    .A2(\u_cpu.ALU._0664_ ),
    .B1(\u_cpu.ALU._0693_ ),
    .Y(\u_cpu.ALU._1170_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2032_  (.A1(\u_cpu.ALU._0664_ ),
    .A2(\u_cpu.ALU._1166_ ),
    .B1(\u_cpu.ALU._1170_ ),
    .Y(\u_cpu.ALU._1171_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2033_  (.A(\u_cpu.ALU._1169_ ),
    .B(\u_cpu.ALU._1171_ ),
    .Y(\u_cpu.ALU._1172_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2034_  (.A1(\u_cpu.ALU._1067_ ),
    .A2(\u_cpu.ALU._1066_ ),
    .B1(\u_cpu.ALU._1069_ ),
    .C1(\u_cpu.ALU._1031_ ),
    .D1(\u_cpu.ALU._1032_ ),
    .X(\u_cpu.ALU._1173_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU._2035_  (.A(\u_cpu.ALU._1103_ ),
    .B(\u_cpu.ALU._1104_ ),
    .C(\u_cpu.ALU._1137_ ),
    .D(\u_cpu.ALU._1140_ ),
    .X(\u_cpu.ALU._1174_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU._2036_  (.A1_N(\u_cpu.ALU._1032_ ),
    .A2_N(\u_cpu.ALU._1069_ ),
    .B1(\u_cpu.ALU._1066_ ),
    .B2(\u_cpu.ALU._1067_ ),
    .Y(\u_cpu.ALU._1175_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU._2037_  (.A(\u_cpu.ALU._1103_ ),
    .B(\u_cpu.ALU._1104_ ),
    .C(\u_cpu.ALU._1137_ ),
    .D(\u_cpu.ALU._1140_ ),
    .Y(\u_cpu.ALU._1176_ ));
 sky130_fd_sc_hd__a21bo_2 \u_cpu.ALU._2038_  (.A1(\u_cpu.ALU._1103_ ),
    .A2(\u_cpu.ALU._1137_ ),
    .B1_N(\u_cpu.ALU._1140_ ),
    .X(\u_cpu.ALU._1177_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2039_  (.A1(\u_cpu.ALU._1175_ ),
    .A2(\u_cpu.ALU._1176_ ),
    .B1(\u_cpu.ALU._1177_ ),
    .Y(\u_cpu.ALU._1178_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU._2040_  (.A1(\u_cpu.ALU._1038_ ),
    .A2(\u_cpu.ALU._1173_ ),
    .A3(\u_cpu.ALU._1174_ ),
    .B1(\u_cpu.ALU._1178_ ),
    .Y(\u_cpu.ALU._1179_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2041_  (.A(\u_cpu.ALU._1172_ ),
    .B(\u_cpu.ALU._1179_ ),
    .Y(\u_cpu.ALU._1180_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._2042_  (.A(\u_cpu.ALU._1169_ ),
    .B(\u_cpu.ALU._1171_ ),
    .X(\u_cpu.ALU._1181_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2043_  (.A1(\u_cpu.ALU._1175_ ),
    .A2(\u_cpu.ALU._1176_ ),
    .B1(\u_cpu.ALU._1177_ ),
    .X(\u_cpu.ALU._1182_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.ALU._2044_  (.A1(\u_cpu.ALU._1108_ ),
    .A2(\u_cpu.ALU._1176_ ),
    .A3(\u_cpu.ALU._1028_ ),
    .B1(\u_cpu.ALU._1182_ ),
    .Y(\u_cpu.ALU._1183_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2045_  (.A1(\u_cpu.ALU._1181_ ),
    .A2(\u_cpu.ALU._1183_ ),
    .B1(\u_cpu.ALU._0975_ ),
    .Y(\u_cpu.ALU._1184_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2046_  (.A(\u_cpu.ALU._0647_ ),
    .B(\u_cpu.ALU._0994_ ),
    .Y(\u_cpu.ALU._1185_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU._2047_  (.A1(\u_cpu.ALU._0881_ ),
    .A2(\u_cpu.ALU._1185_ ),
    .B1(\u_cpu.ALU._0766_ ),
    .B2(\u_cpu.ALU._0770_ ),
    .Y(\u_cpu.ALU._1186_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2048_  (.A0(\u_cpu.ALU._0802_ ),
    .A1(\u_cpu.ALU._0803_ ),
    .A2(\u_cpu.ALU._0767_ ),
    .A3(\u_cpu.ALU._0779_ ),
    .S0(\u_cpu.ALU._0765_ ),
    .S1(\u_cpu.ALU._0623_ ),
    .X(\u_cpu.ALU._1187_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2049_  (.A(\u_cpu.ALU._0817_ ),
    .B(\u_cpu.ALU._1187_ ),
    .Y(\u_cpu.ALU._1188_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2050_  (.A1(\u_cpu.ALU._0817_ ),
    .A2(\u_cpu.ALU._1186_ ),
    .B1(\u_cpu.ALU._1188_ ),
    .X(\u_cpu.ALU._1189_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2051_  (.A1(\u_cpu.ALU._0693_ ),
    .A2(\u_cpu.ALU._1163_ ),
    .B1(\u_cpu.ALU._0737_ ),
    .C1(\u_cpu.ALU._0900_ ),
    .D1(\u_cpu.ALU._0811_ ),
    .X(\u_cpu.ALU._1190_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU._2052_  (.A1(\u_cpu.ALU._0663_ ),
    .A2(\u_cpu.ALU._0664_ ),
    .B1(\u_cpu.ALU._0748_ ),
    .B2(\u_cpu.ALU._1190_ ),
    .X(\u_cpu.ALU._1191_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._2053_  (.A1(\u_cpu.ALU._0957_ ),
    .A2(\u_cpu.ALU._0663_ ),
    .B1(\u_cpu.ALU._0664_ ),
    .C1(\u_cpu.ALU._0896_ ),
    .X(\u_cpu.ALU._1192_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU._2054_  (.A1(\u_cpu.ALU.Product_Wallace[8] ),
    .A2(\u_cpu.ALU._0821_ ),
    .B1(\u_cpu.ALU._1191_ ),
    .C1(\u_cpu.ALU._1192_ ),
    .Y(\u_cpu.ALU._1193_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2055_  (.A0(\u_cpu.ALU._0663_ ),
    .A1(\u_cpu.ALU._0598_ ),
    .A2(\u_cpu.ALU.SrcA[6] ),
    .A3(\u_cpu.ALU.SrcA[5] ),
    .S0(\u_cpu.ALU._0775_ ),
    .S1(\u_cpu.ALU._0638_ ),
    .X(\u_cpu.ALU._1194_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.ALU._2056_  (.A0(\u_cpu.ALU._1045_ ),
    .A1(\u_cpu.ALU._1194_ ),
    .S(\u_cpu.ALU._0768_ ),
    .X(\u_cpu.ALU._1195_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU._2057_  (.A1(\u_cpu.ALU.SrcA[0] ),
    .A2(\u_cpu.ALU._0911_ ),
    .A3(\u_cpu.ALU._1057_ ),
    .B1(\u_cpu.ALU._1195_ ),
    .B2(\u_cpu.ALU._1088_ ),
    .X(\u_cpu.ALU._1196_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._2058_  (.A(\u_cpu.ALU._0879_ ),
    .B(\u_cpu.ALU._1196_ ),
    .C(\u_cpu.ALU._1077_ ),
    .Y(\u_cpu.ALU._1197_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._2059_  (.A1(\u_cpu.ALU._0784_ ),
    .A2(\u_cpu.ALU._1189_ ),
    .B1(\u_cpu.ALU._1193_ ),
    .C1(\u_cpu.ALU._1197_ ),
    .X(\u_cpu.ALU._1198_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2060_  (.A1(\u_cpu.ALU._1180_ ),
    .A2(\u_cpu.ALU._1184_ ),
    .B1(\u_cpu.ALU._1198_ ),
    .Y(\u_cpu.ALU.ALUResult[8] ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2061_  (.A(\u_cpu.ALU._1183_ ),
    .B(\u_cpu.ALU._1181_ ),
    .Y(\u_cpu.ALU._1199_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2062_  (.A(\u_cpu.ALU._0914_ ),
    .X(\u_cpu.ALU._1200_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._2063_  (.A1(\u_cpu.ALU._1200_ ),
    .A2(\u_cpu.ALU._1163_ ),
    .B1(\u_cpu.ALU._0691_ ),
    .C1(\u_cpu.ALU._1166_ ),
    .X(\u_cpu.ALU._1201_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU._2064_  (.A(\u_cpu.ALU._0613_ ),
    .B(\u_cpu.ALU.SrcB[7] ),
    .C(\u_cpu.ALU.SrcB[5] ),
    .Y(\u_cpu.ALU._1202_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU._2065_  (.A(\u_cpu.ALU._0911_ ),
    .B(\u_cpu.ALU._0960_ ),
    .C(\u_cpu.ALU._1202_ ),
    .D(\u_cpu.ALU._0604_ ),
    .Y(\u_cpu.ALU._1203_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU._2066_  (.A1(\u_cpu.ALU._0710_ ),
    .A2(\u_cpu.ALU._0919_ ),
    .B1(\u_cpu.ALU._0664_ ),
    .B2(\u_cpu.ALU._1203_ ),
    .C1(\u_cpu.ALU.SrcB[9] ),
    .Y(\u_cpu.ALU._1204_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2067_  (.A(\u_cpu.ALU._0862_ ),
    .B(\u_cpu.ALU._1204_ ),
    .Y(\u_cpu.ALU._1205_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._2068_  (.A1(\u_cpu.ALU._0914_ ),
    .A2(\u_cpu.ALU._1163_ ),
    .B1(\u_cpu.ALU._0691_ ),
    .C1(\u_cpu.ALU._1166_ ),
    .Y(\u_cpu.ALU._1206_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2069_  (.A1(\u_cpu.ALU._1204_ ),
    .A2(\u_cpu.ALU._1206_ ),
    .B1(\u_cpu.ALU._0862_ ),
    .X(\u_cpu.ALU._1207_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2070_  (.A1(\u_cpu.ALU._1201_ ),
    .A2(\u_cpu.ALU._1205_ ),
    .B1(\u_cpu.ALU._1207_ ),
    .Y(\u_cpu.ALU._1208_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2071_  (.A1(\u_cpu.ALU._1171_ ),
    .A2(\u_cpu.ALU._1199_ ),
    .B1(\u_cpu.ALU._1208_ ),
    .X(\u_cpu.ALU._1209_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU._2072_  (.A1(\u_cpu.ALU._1171_ ),
    .A2(\u_cpu.ALU._1199_ ),
    .A3(\u_cpu.ALU._1208_ ),
    .B1(\u_cpu.ALU._0921_ ),
    .Y(\u_cpu.ALU._1210_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2073_  (.A(\u_cpu.ALU._1209_ ),
    .B(\u_cpu.ALU._1210_ ),
    .Y(\u_cpu.ALU._1211_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2074_  (.A(\u_cpu.ALU._1076_ ),
    .X(\u_cpu.ALU._1212_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU._2075_  (.A1(\u_cpu.ALU._0761_ ),
    .A2(\u_cpu.ALU._0836_ ),
    .B1_N(\u_cpu.ALU._1185_ ),
    .Y(\u_cpu.ALU._1213_ ));
 sky130_fd_sc_hd__a32oi_2 \u_cpu.ALU._2076_  (.A1(\u_cpu.ALU._1212_ ),
    .A2(\u_cpu.ALU._0877_ ),
    .A3(\u_cpu.ALU._0882_ ),
    .B1(\u_cpu.ALU._1213_ ),
    .B2(\u_cpu.ALU._0874_ ),
    .Y(\u_cpu.ALU._1214_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2077_  (.A1(\u_cpu.ALU._0862_ ),
    .A2(\u_cpu.ALU._0691_ ),
    .B1(\u_cpu.ALU._0737_ ),
    .C1(\u_cpu.ALU._0900_ ),
    .D1(\u_cpu.ALU._0890_ ),
    .X(\u_cpu.ALU._1215_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU._2078_  (.A1(\u_cpu.ALU._0669_ ),
    .A2(\u_cpu.ALU.SrcB[9] ),
    .B1(\u_cpu.ALU._0749_ ),
    .B2(\u_cpu.ALU._1215_ ),
    .X(\u_cpu.ALU._1216_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._2079_  (.A1(\u_cpu.ALU._0957_ ),
    .A2(\u_cpu.ALU._0669_ ),
    .B1(\u_cpu.ALU.SrcB[9] ),
    .C1(\u_cpu.ALU._0896_ ),
    .X(\u_cpu.ALU._1217_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU._2080_  (.A1(\u_cpu.ALU.Product_Wallace[9] ),
    .A2(\u_cpu.ALU._0822_ ),
    .B1(\u_cpu.ALU._1216_ ),
    .C1(\u_cpu.ALU._1217_ ),
    .Y(\u_cpu.ALU._1218_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2081_  (.A(\u_cpu.ALU._1088_ ),
    .X(\u_cpu.ALU._1219_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2082_  (.A1(\u_cpu.ALU._1145_ ),
    .A2(\u_cpu.ALU._0839_ ),
    .B1(\u_cpu.ALU._0846_ ),
    .X(\u_cpu.ALU._1220_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.ALU._2083_  (.A1(\u_cpu.ALU._1145_ ),
    .A2(\u_cpu.ALU._0861_ ),
    .A3(\u_cpu.ALU._0864_ ),
    .B1(\u_cpu.ALU._0869_ ),
    .C1(\u_cpu.ALU._1076_ ),
    .Y(\u_cpu.ALU._1221_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._2084_  (.A1(\u_cpu.ALU._1219_ ),
    .A2(\u_cpu.ALU._1220_ ),
    .B1(\u_cpu.ALU._1221_ ),
    .C1(\u_cpu.ALU._1158_ ),
    .X(\u_cpu.ALU._1222_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2085_  (.A0(\u_cpu.ALU._0669_ ),
    .A1(\u_cpu.ALU._0663_ ),
    .A2(\u_cpu.ALU._0598_ ),
    .A3(\u_cpu.ALU.SrcA[6] ),
    .S0(\u_cpu.ALU._0838_ ),
    .S1(\u_cpu.ALU._0728_ ),
    .X(\u_cpu.ALU._1223_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.ALU._2086_  (.A0(\u_cpu.ALU._1078_ ),
    .A1(\u_cpu.ALU._1223_ ),
    .S(\u_cpu.ALU._0768_ ),
    .X(\u_cpu.ALU._1224_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU._2087_  (.A1(\u_cpu.ALU._0893_ ),
    .A2(\u_cpu.ALU._1057_ ),
    .B1(\u_cpu.ALU._1224_ ),
    .B2(\u_cpu.ALU._1088_ ),
    .X(\u_cpu.ALU._1225_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2088_  (.A(\u_cpu.ALU._0881_ ),
    .X(\u_cpu.ALU._1226_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU._2089_  (.A(\u_cpu.ALU._1225_ ),
    .B(\u_cpu.ALU._0738_ ),
    .C(\u_cpu.ALU._1226_ ),
    .D(\u_cpu.ALU._0963_ ),
    .X(\u_cpu.ALU._1227_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2090_  (.A1(\u_cpu.ALU._1222_ ),
    .A2(\u_cpu.ALU._1227_ ),
    .B1(\u_cpu.ALU._1075_ ),
    .Y(\u_cpu.ALU._1228_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._2091_  (.A1(\u_cpu.ALU._1075_ ),
    .A2(\u_cpu.ALU._1214_ ),
    .B1(\u_cpu.ALU._1218_ ),
    .C1(\u_cpu.ALU._1228_ ),
    .X(\u_cpu.ALU._1229_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2092_  (.A(\u_cpu.ALU._1211_ ),
    .B(\u_cpu.ALU._1229_ ),
    .Y(\u_cpu.ALU.ALUResult[9] ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2093_  (.A1(\u_cpu.ALU._1205_ ),
    .A2(\u_cpu.ALU._1201_ ),
    .B1(\u_cpu.ALU._1171_ ),
    .C1(\u_cpu.ALU._1169_ ),
    .D1(\u_cpu.ALU._1207_ ),
    .X(\u_cpu.ALU._1230_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._2094_  (.A(\u_cpu.ALU._1230_ ),
    .Y(\u_cpu.ALU._1231_ ));
 sky130_fd_sc_hd__nor4_2 \u_cpu.ALU._2095_  (.A(\u_cpu.ALU.SrcB[4] ),
    .B(\u_cpu.ALU.SrcB[7] ),
    .C(\u_cpu.ALU.SrcB[6] ),
    .D(\u_cpu.ALU.SrcB[5] ),
    .Y(\u_cpu.ALU._1232_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2096_  (.A(\u_cpu.ALU.SrcB[9] ),
    .B(\u_cpu.ALU._0664_ ),
    .Y(\u_cpu.ALU._1233_ ));
 sky130_fd_sc_hd__a311o_2 \u_cpu.ALU._2097_  (.A1(\u_cpu.ALU._0801_ ),
    .A2(\u_cpu.ALU._1232_ ),
    .A3(\u_cpu.ALU._1233_ ),
    .B1(\u_cpu.ALU._0914_ ),
    .C1(\u_cpu.ALU._0667_ ),
    .X(\u_cpu.ALU._1234_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._2098_  (.A1(\u_cpu.ALU._0914_ ),
    .A2(\u_cpu.ALU._1233_ ),
    .B1(\u_cpu.ALU._0667_ ),
    .C1(\u_cpu.ALU._1166_ ),
    .Y(\u_cpu.ALU._1235_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._2099_  (.A(\u_cpu.ALU._1234_ ),
    .B(\u_cpu.ALU._1235_ ),
    .C(\u_cpu.ALU._0666_ ),
    .Y(\u_cpu.ALU._1236_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU._2100_  (.A1(\u_cpu.ALU._0801_ ),
    .A2(\u_cpu.ALU._1232_ ),
    .A3(\u_cpu.ALU._1233_ ),
    .B1(\u_cpu.ALU._0914_ ),
    .Y(\u_cpu.ALU._1237_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2101_  (.A1(\u_cpu.ALU._1237_ ),
    .A2(\u_cpu.ALU._0667_ ),
    .B1(\u_cpu.ALU.SrcA[10] ),
    .Y(\u_cpu.ALU._1238_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2102_  (.A1(\u_cpu.ALU._0667_ ),
    .A2(\u_cpu.ALU._1237_ ),
    .B1(\u_cpu.ALU._1238_ ),
    .Y(\u_cpu.ALU._1239_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2103_  (.A(\u_cpu.ALU._1236_ ),
    .B(\u_cpu.ALU._1239_ ),
    .Y(\u_cpu.ALU._1240_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2104_  (.A1(\u_cpu.ALU._1167_ ),
    .A2(\u_cpu.ALU._1168_ ),
    .B1(\u_cpu.ALU._0693_ ),
    .Y(\u_cpu.ALU._1241_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2105_  (.A1(\u_cpu.ALU._1204_ ),
    .A2(\u_cpu.ALU._1206_ ),
    .B1(\u_cpu.ALU._0862_ ),
    .Y(\u_cpu.ALU._1242_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU._2106_  (.A1(\u_cpu.ALU._1205_ ),
    .A2(\u_cpu.ALU._1201_ ),
    .B1(\u_cpu.ALU._1241_ ),
    .B2(\u_cpu.ALU._1242_ ),
    .Y(\u_cpu.ALU._1243_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._2107_  (.A1(\u_cpu.ALU._1231_ ),
    .A2(\u_cpu.ALU._1179_ ),
    .B1(\u_cpu.ALU._1240_ ),
    .C1(\u_cpu.ALU._1243_ ),
    .Y(\u_cpu.ALU._1244_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2108_  (.A1(\u_cpu.ALU._1231_ ),
    .A2(\u_cpu.ALU._1179_ ),
    .B1(\u_cpu.ALU._1243_ ),
    .Y(\u_cpu.ALU._1245_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._2109_  (.A(\u_cpu.ALU._1236_ ),
    .B(\u_cpu.ALU._1239_ ),
    .X(\u_cpu.ALU._1246_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2110_  (.A(\u_cpu.ALU._1245_ ),
    .B(\u_cpu.ALU._1246_ ),
    .Y(\u_cpu.ALU._1247_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2111_  (.A1(\u_cpu.ALU._1088_ ),
    .A2(\u_cpu.ALU._0970_ ),
    .B1(\u_cpu.ALU._1185_ ),
    .X(\u_cpu.ALU._1248_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU._2112_  (.A1(\u_cpu.ALU._1219_ ),
    .A2(\u_cpu.ALU._0882_ ),
    .A3(\u_cpu.ALU._0932_ ),
    .B1(\u_cpu.ALU._1248_ ),
    .B2(\u_cpu.ALU._0874_ ),
    .X(\u_cpu.ALU._1249_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2113_  (.A1(\u_cpu.ALU._0666_ ),
    .A2(\u_cpu.ALU._0667_ ),
    .B1(\u_cpu.ALU._1020_ ),
    .Y(\u_cpu.ALU._1250_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU._2114_  (.A1(\u_cpu.ALU._0666_ ),
    .A2(\u_cpu.ALU._0667_ ),
    .B1(\u_cpu.ALU._0748_ ),
    .B2(\u_cpu.ALU._1250_ ),
    .X(\u_cpu.ALU._1251_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._2115_  (.A1(\u_cpu.ALU._0957_ ),
    .A2(\u_cpu.ALU._0666_ ),
    .B1(\u_cpu.ALU._0667_ ),
    .C1(\u_cpu.ALU._0896_ ),
    .X(\u_cpu.ALU._1252_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._2116_  (.A1(\u_cpu.ALU.Product_Wallace[10] ),
    .A2(\u_cpu.ALU._0821_ ),
    .B1(\u_cpu.ALU._1251_ ),
    .C1(\u_cpu.ALU._1252_ ),
    .X(\u_cpu.ALU._1253_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._2117_  (.A(\u_cpu.ALU._0940_ ),
    .B(\u_cpu.ALU._0805_ ),
    .C(\u_cpu.ALU._0936_ ),
    .X(\u_cpu.ALU._1254_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._2118_  (.A(\u_cpu.ALU._1088_ ),
    .B(\u_cpu.ALU._0952_ ),
    .C(\u_cpu.ALU._0950_ ),
    .Y(\u_cpu.ALU._1255_ ));
 sky130_fd_sc_hd__or3b_2 \u_cpu.ALU._2119_  (.A(\u_cpu.ALU._1254_ ),
    .B(\u_cpu.ALU._0783_ ),
    .C_N(\u_cpu.ALU._1255_ ),
    .X(\u_cpu.ALU._1256_ ));
 sky130_fd_sc_hd__or4b_2 \u_cpu.ALU._2120_  (.A(\u_cpu.ALU._0811_ ),
    .B(\u_cpu.ALU._0873_ ),
    .C(\u_cpu.ALU._0751_ ),
    .D_N(\u_cpu.ALU._0750_ ),
    .X(\u_cpu.ALU._1257_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2121_  (.A0(\u_cpu.ALU.SrcA[10] ),
    .A1(\u_cpu.ALU._0669_ ),
    .A2(\u_cpu.ALU._0663_ ),
    .A3(\u_cpu.ALU._0598_ ),
    .S0(\u_cpu.ALU._0840_ ),
    .S1(\u_cpu.ALU._0638_ ),
    .X(\u_cpu.ALU._1258_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU._2122_  (.A1(\u_cpu.ALU._0643_ ),
    .A2(\u_cpu.ALU._0788_ ),
    .A3(\u_cpu.ALU._0793_ ),
    .B1(\u_cpu.ALU._1113_ ),
    .C1(\u_cpu.ALU._0629_ ),
    .X(\u_cpu.ALU._1259_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2123_  (.A1(\u_cpu.ALU._1258_ ),
    .A2(\u_cpu.ALU._0768_ ),
    .B1(\u_cpu.ALU._1259_ ),
    .Y(\u_cpu.ALU._1260_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU._2124_  (.A1_N(\u_cpu.ALU._0962_ ),
    .A2_N(\u_cpu.ALU._1057_ ),
    .B1(\u_cpu.ALU._0760_ ),
    .B2(\u_cpu.ALU._1260_ ),
    .X(\u_cpu.ALU._1261_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU._2125_  (.A(\u_cpu.ALU._1257_ ),
    .B(\u_cpu.ALU._1261_ ),
    .X(\u_cpu.ALU._1262_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2126_  (.A1(\u_cpu.ALU._1256_ ),
    .A2(\u_cpu.ALU._1262_ ),
    .B1(\u_cpu.ALU._0759_ ),
    .Y(\u_cpu.ALU._1263_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._2127_  (.A1(\u_cpu.ALU._1144_ ),
    .A2(\u_cpu.ALU._1249_ ),
    .B1(\u_cpu.ALU._1253_ ),
    .C1(\u_cpu.ALU._1263_ ),
    .X(\u_cpu.ALU._1264_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._2128_  (.A1(\u_cpu.ALU._0975_ ),
    .A2(\u_cpu.ALU._1244_ ),
    .A3(\u_cpu.ALU._1247_ ),
    .B1(\u_cpu.ALU._1264_ ),
    .X(\u_cpu.ALU.ALUResult[10] ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._2129_  (.A(\u_cpu.ALU._1234_ ),
    .B(\u_cpu.ALU._1235_ ),
    .C(\u_cpu.ALU.SrcA[10] ),
    .X(\u_cpu.ALU._1265_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._2130_  (.A1(\u_cpu.ALU._0741_ ),
    .A2(\u_cpu.ALU._0811_ ),
    .A3(\u_cpu.ALU._0745_ ),
    .B1(\u_cpu.ALU._1233_ ),
    .X(\u_cpu.ALU._1266_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU._2131_  (.A1(\u_cpu.ALU._0914_ ),
    .A2(\u_cpu.ALU._0689_ ),
    .B1(\u_cpu.ALU._0687_ ),
    .C1(\u_cpu.ALU._1266_ ),
    .D1(\u_cpu.ALU._1166_ ),
    .Y(\u_cpu.ALU._1267_ ));
 sky130_fd_sc_hd__a41oi_2 \u_cpu.ALU._2132_  (.A1(\u_cpu.ALU._0801_ ),
    .A2(\u_cpu.ALU._1232_ ),
    .A3(\u_cpu.ALU._1233_ ),
    .A4(\u_cpu.ALU._0689_ ),
    .B1(\u_cpu.ALU._0914_ ),
    .Y(\u_cpu.ALU._1268_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2133_  (.A1(\u_cpu.ALU._1268_ ),
    .A2(\u_cpu.ALU.SrcB[11] ),
    .B1(\u_cpu.ALU._0686_ ),
    .Y(\u_cpu.ALU._1269_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2134_  (.A(\u_cpu.ALU._1268_ ),
    .B(\u_cpu.ALU.SrcB[11] ),
    .Y(\u_cpu.ALU._1270_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2135_  (.A1(\u_cpu.ALU._1270_ ),
    .A2(\u_cpu.ALU._1267_ ),
    .B1(\u_cpu.ALU._0858_ ),
    .Y(\u_cpu.ALU._1271_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2136_  (.A1(\u_cpu.ALU._1267_ ),
    .A2(\u_cpu.ALU._1269_ ),
    .B1(\u_cpu.ALU._1271_ ),
    .Y(\u_cpu.ALU._1272_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU._2137_  (.A1(\u_cpu.ALU._1245_ ),
    .A2(\u_cpu.ALU._1246_ ),
    .B1(\u_cpu.ALU._1265_ ),
    .C1(\u_cpu.ALU._1272_ ),
    .Y(\u_cpu.ALU._1273_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.ALU._2138_  (.A1(\u_cpu.ALU._1269_ ),
    .A2(\u_cpu.ALU._1267_ ),
    .B1(\u_cpu.ALU._1247_ ),
    .B2(\u_cpu.ALU._1236_ ),
    .C1(\u_cpu.ALU._1271_ ),
    .Y(\u_cpu.ALU._1274_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2139_  (.A(\u_cpu.ALU._1075_ ),
    .X(\u_cpu.ALU._1275_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2140_  (.A0(\u_cpu.ALU._0686_ ),
    .A1(\u_cpu.ALU._0666_ ),
    .A2(\u_cpu.ALU._0669_ ),
    .A3(\u_cpu.ALU._0663_ ),
    .S0(\u_cpu.ALU._0722_ ),
    .S1(\u_cpu.ALU._0729_ ),
    .X(\u_cpu.ALU._1276_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.ALU._2141_  (.A0(\u_cpu.ALU._1155_ ),
    .A1(\u_cpu.ALU._1276_ ),
    .S(\u_cpu.ALU._0769_ ),
    .X(\u_cpu.ALU._1277_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU._2142_  (.A1(\u_cpu.ALU._1017_ ),
    .A2(\u_cpu.ALU._1057_ ),
    .B1(\u_cpu.ALU._1277_ ),
    .B2(\u_cpu.ALU._1219_ ),
    .Y(\u_cpu.ALU._1278_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2143_  (.A(\u_cpu.ALU._0786_ ),
    .X(\u_cpu.ALU._1279_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2144_  (.A0(\u_cpu.ALU._1146_ ),
    .A1(\u_cpu.ALU._1012_ ),
    .A2(\u_cpu.ALU._1002_ ),
    .A3(\u_cpu.ALU._1011_ ),
    .S0(\u_cpu.ALU._1076_ ),
    .S1(\u_cpu.ALU._1279_ ),
    .X(\u_cpu.ALU._1280_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.ALU._2145_  (.A1_N(\u_cpu.ALU._1257_ ),
    .A2_N(\u_cpu.ALU._1278_ ),
    .B1(\u_cpu.ALU._1280_ ),
    .B2(\u_cpu.ALU._1158_ ),
    .X(\u_cpu.ALU._1281_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2146_  (.A(\u_cpu.ALU._1275_ ),
    .B(\u_cpu.ALU._1281_ ),
    .Y(\u_cpu.ALU._1282_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2147_  (.A(\u_cpu.ALU._1144_ ),
    .X(\u_cpu.ALU._1283_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU._2148_  (.A1(\u_cpu.ALU._0729_ ),
    .A2(\u_cpu.ALU._0831_ ),
    .A3(\u_cpu.ALU._0832_ ),
    .B1(\u_cpu.ALU._0999_ ),
    .X(\u_cpu.ALU._1284_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.ALU._2149_  (.A0(\u_cpu.ALU._1284_ ),
    .A1(\u_cpu.ALU._0577_ ),
    .S(\u_cpu.ALU._0958_ ),
    .X(\u_cpu.ALU._1285_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU._2150_  (.A1(\u_cpu.ALU._0874_ ),
    .A2(\u_cpu.ALU._1185_ ),
    .B1(\u_cpu.ALU._1285_ ),
    .B2(\u_cpu.ALU._1212_ ),
    .Y(\u_cpu.ALU._1286_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU._2151_  (.A1(\u_cpu.ALU._1149_ ),
    .A2(\u_cpu.ALU._1005_ ),
    .B1(\u_cpu.ALU._0784_ ),
    .C1(\u_cpu.ALU._1286_ ),
    .Y(\u_cpu.ALU._1287_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._2152_  (.A1(\u_cpu.ALU._0957_ ),
    .A2(\u_cpu.ALU._0686_ ),
    .B1(\u_cpu.ALU.SrcB[11] ),
    .C1(\u_cpu.ALU._0896_ ),
    .X(\u_cpu.ALU._1288_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2153_  (.A1(\u_cpu.ALU._0858_ ),
    .A2(\u_cpu.ALU._0687_ ),
    .B1(\u_cpu.ALU._0737_ ),
    .C1(\u_cpu.ALU._1149_ ),
    .D1(\u_cpu.ALU._0890_ ),
    .X(\u_cpu.ALU._1289_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU._2154_  (.A1(\u_cpu.ALU._0686_ ),
    .A2(\u_cpu.ALU.SrcB[11] ),
    .B1(\u_cpu.ALU._0749_ ),
    .B2(\u_cpu.ALU._1289_ ),
    .X(\u_cpu.ALU._1290_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._2155_  (.A1(\u_cpu.ALU.Product_Wallace[11] ),
    .A2(\u_cpu.ALU._0822_ ),
    .B1(\u_cpu.ALU._1288_ ),
    .C1(\u_cpu.ALU._1290_ ),
    .X(\u_cpu.ALU._1291_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2156_  (.A1(\u_cpu.ALU._1283_ ),
    .A2(\u_cpu.ALU._1287_ ),
    .B1(\u_cpu.ALU._1291_ ),
    .Y(\u_cpu.ALU._1292_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.ALU._2157_  (.A1(\u_cpu.ALU._1273_ ),
    .A2(\u_cpu.ALU._0921_ ),
    .A3(\u_cpu.ALU._1274_ ),
    .B1(\u_cpu.ALU._1282_ ),
    .C1(\u_cpu.ALU._1292_ ),
    .Y(\u_cpu.ALU.ALUResult[11] ));
 sky130_fd_sc_hd__nor4_2 \u_cpu.ALU._2158_  (.A(\u_cpu.ALU.SrcB[11] ),
    .B(\u_cpu.ALU.SrcB[10] ),
    .C(\u_cpu.ALU.SrcB[9] ),
    .D(\u_cpu.ALU.SrcB[8] ),
    .Y(\u_cpu.ALU._1293_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._2159_  (.A1(\u_cpu.ALU._0801_ ),
    .A2(\u_cpu.ALU._1232_ ),
    .A3(\u_cpu.ALU._1293_ ),
    .B1(\u_cpu.ALU._0660_ ),
    .X(\u_cpu.ALU._1294_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2160_  (.A1(\u_cpu.ALU._0746_ ),
    .A2(\u_cpu.ALU._0814_ ),
    .B1(\u_cpu.ALU._1294_ ),
    .Y(\u_cpu.ALU._1295_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2161_  (.A(\u_cpu.ALU.SrcB[11] ),
    .B(\u_cpu.ALU._0667_ ),
    .Y(\u_cpu.ALU._1296_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU._2162_  (.A(\u_cpu.ALU._1202_ ),
    .B(\u_cpu.ALU._1233_ ),
    .C(\u_cpu.ALU._1296_ ),
    .D(\u_cpu.ALU._0604_ ),
    .Y(\u_cpu.ALU._1297_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2163_  (.A1(\u_cpu.ALU._1165_ ),
    .A2(\u_cpu.ALU._1297_ ),
    .B1(\u_cpu.ALU._0985_ ),
    .Y(\u_cpu.ALU._1298_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2164_  (.A1(\u_cpu.ALU._1298_ ),
    .A2(\u_cpu.ALU._0660_ ),
    .B1(\u_cpu.ALU._0676_ ),
    .X(\u_cpu.ALU._1299_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2165_  (.A(\u_cpu.ALU._1298_ ),
    .B(\u_cpu.ALU._0660_ ),
    .Y(\u_cpu.ALU._1300_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2166_  (.A1(\u_cpu.ALU._1200_ ),
    .A2(\u_cpu.ALU._1294_ ),
    .B1(\u_cpu.ALU._1300_ ),
    .Y(\u_cpu.ALU._1301_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2167_  (.A(\u_cpu.ALU._1301_ ),
    .B(\u_cpu.ALU._0676_ ),
    .Y(\u_cpu.ALU._1302_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2168_  (.A1(\u_cpu.ALU._1295_ ),
    .A2(\u_cpu.ALU._1299_ ),
    .B1(\u_cpu.ALU._1302_ ),
    .Y(\u_cpu.ALU._1303_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2169_  (.A1(\u_cpu.ALU.SrcB[11] ),
    .A2(\u_cpu.ALU._1268_ ),
    .B1(\u_cpu.ALU._1269_ ),
    .Y(\u_cpu.ALU._1304_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2170_  (.A(\u_cpu.ALU._1265_ ),
    .B(\u_cpu.ALU._1271_ ),
    .Y(\u_cpu.ALU._1305_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2171_  (.A1(\u_cpu.ALU._1240_ ),
    .A2(\u_cpu.ALU._1243_ ),
    .B1(\u_cpu.ALU._1305_ ),
    .Y(\u_cpu.ALU._1306_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._2172_  (.A(\u_cpu.ALU._1246_ ),
    .B(\u_cpu.ALU._1230_ ),
    .C(\u_cpu.ALU._1272_ ),
    .X(\u_cpu.ALU._1307_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU._2173_  (.A1(\u_cpu.ALU._1304_ ),
    .A2(\u_cpu.ALU._1306_ ),
    .B1(\u_cpu.ALU._1183_ ),
    .B2(\u_cpu.ALU._1307_ ),
    .Y(\u_cpu.ALU._1308_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2174_  (.A(\u_cpu.ALU._1303_ ),
    .B(\u_cpu.ALU._1308_ ),
    .Y(\u_cpu.ALU._1309_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2175_  (.A1(\u_cpu.ALU._1308_ ),
    .A2(\u_cpu.ALU._1303_ ),
    .B1(\u_cpu.ALU._0921_ ),
    .X(\u_cpu.ALU._1310_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2176_  (.A1(\u_cpu.ALU._0958_ ),
    .A2(\u_cpu.ALU._0802_ ),
    .B1(\u_cpu.ALU._1042_ ),
    .X(\u_cpu.ALU._1311_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2177_  (.A1(\u_cpu.ALU._0797_ ),
    .A2(\u_cpu.ALU._0767_ ),
    .B1(\u_cpu.ALU._1055_ ),
    .Y(\u_cpu.ALU._1312_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2178_  (.A1(\u_cpu.ALU._1312_ ),
    .A2(\u_cpu.ALU._0760_ ),
    .B1(\u_cpu.ALU._0757_ ),
    .Y(\u_cpu.ALU._1313_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2179_  (.A1(\u_cpu.ALU._0806_ ),
    .A2(\u_cpu.ALU._1311_ ),
    .B1(\u_cpu.ALU._1313_ ),
    .X(\u_cpu.ALU._1314_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._2180_  (.A1(\u_cpu.ALU._0758_ ),
    .A2(\u_cpu.ALU._0960_ ),
    .A3(\u_cpu.ALU._0762_ ),
    .B1(\u_cpu.ALU._1314_ ),
    .X(\u_cpu.ALU._1315_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._2181_  (.A(\u_cpu.ALU._0762_ ),
    .B(\u_cpu.ALU._0785_ ),
    .C(\u_cpu.ALU._0770_ ),
    .X(\u_cpu.ALU._1316_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2182_  (.A1(\u_cpu.ALU._0760_ ),
    .A2(\u_cpu.ALU._0958_ ),
    .B1(\u_cpu.ALU._0577_ ),
    .X(\u_cpu.ALU._1317_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2183_  (.A1(\u_cpu.ALU._1316_ ),
    .A2(\u_cpu.ALU._1317_ ),
    .B1(\u_cpu.ALU._0757_ ),
    .X(\u_cpu.ALU._1318_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._2184_  (.A1(\u_cpu.ALU._1314_ ),
    .A2(\u_cpu.ALU._1318_ ),
    .B1(\u_cpu.ALU._1226_ ),
    .C1(\u_cpu.ALU._1158_ ),
    .X(\u_cpu.ALU._1319_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2185_  (.A1(\u_cpu.ALU._0859_ ),
    .A2(\u_cpu.ALU._0660_ ),
    .B1(\u_cpu.ALU._0749_ ),
    .Y(\u_cpu.ALU._1320_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2186_  (.A0(\u_cpu.ALU._0859_ ),
    .A1(\u_cpu.ALU._0686_ ),
    .A2(\u_cpu.ALU._0666_ ),
    .A3(\u_cpu.ALU._0669_ ),
    .S0(\u_cpu.ALU._0794_ ),
    .S1(\u_cpu.ALU._0826_ ),
    .X(\u_cpu.ALU._1321_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2187_  (.A0(\u_cpu.ALU._1194_ ),
    .A1(\u_cpu.ALU._0644_ ),
    .A2(\u_cpu.ALU._1321_ ),
    .A3(\u_cpu.ALU._1045_ ),
    .S0(\u_cpu.ALU._0805_ ),
    .S1(\u_cpu.ALU._0769_ ),
    .X(\u_cpu.ALU._1322_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU._2188_  (.A1(\u_cpu.ALU._0859_ ),
    .A2(\u_cpu.ALU._0660_ ),
    .A3(\u_cpu.ALU._0744_ ),
    .B1(\u_cpu.ALU._0821_ ),
    .B2(\u_cpu.ALU.Product_Wallace[12] ),
    .X(\u_cpu.ALU._1323_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.ALU._2189_  (.A1(\u_cpu.ALU._0660_ ),
    .A2(\u_cpu.ALU._0754_ ),
    .B1(\u_cpu.ALU._1322_ ),
    .B2(\u_cpu.ALU._0819_ ),
    .C1(\u_cpu.ALU._1323_ ),
    .Y(\u_cpu.ALU._1324_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._2190_  (.A1(\u_cpu.ALU._0661_ ),
    .A2(\u_cpu.ALU._1020_ ),
    .B1(\u_cpu.ALU._1320_ ),
    .C1(\u_cpu.ALU._1324_ ),
    .Y(\u_cpu.ALU._1325_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU._2191_  (.A1(\u_cpu.ALU._0882_ ),
    .A2(\u_cpu.ALU._1315_ ),
    .B1(\u_cpu.ALU._1319_ ),
    .C1(\u_cpu.ALU._1325_ ),
    .Y(\u_cpu.ALU._1326_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2192_  (.A1(\u_cpu.ALU._1309_ ),
    .A2(\u_cpu.ALU._1310_ ),
    .B1(\u_cpu.ALU._1326_ ),
    .Y(\u_cpu.ALU.ALUResult[12] ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2193_  (.A0(\u_cpu.ALU._1085_ ),
    .A1(\u_cpu.ALU._1086_ ),
    .A2(\u_cpu.ALU._1081_ ),
    .A3(\u_cpu.ALU._0839_ ),
    .S0(\u_cpu.ALU._1145_ ),
    .S1(\u_cpu.ALU._1212_ ),
    .X(\u_cpu.ALU._1327_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2194_  (.A(\u_cpu.ALU.SrcA[13] ),
    .X(\u_cpu.ALU._1328_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2195_  (.A0(\u_cpu.ALU._1328_ ),
    .A1(\u_cpu.ALU._0859_ ),
    .A2(\u_cpu.ALU._0686_ ),
    .A3(\u_cpu.ALU._0666_ ),
    .S0(\u_cpu.ALU._0635_ ),
    .S1(\u_cpu.ALU._0726_ ),
    .X(\u_cpu.ALU._1329_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2196_  (.A0(\u_cpu.ALU._1223_ ),
    .A1(\u_cpu.ALU._0893_ ),
    .A2(\u_cpu.ALU._1329_ ),
    .A3(\u_cpu.ALU._1078_ ),
    .S0(\u_cpu.ALU._0806_ ),
    .S1(\u_cpu.ALU._1279_ ),
    .X(\u_cpu.ALU._1330_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2197_  (.A(\u_cpu.ALU._1226_ ),
    .X(\u_cpu.ALU._1331_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2198_  (.A(\u_cpu.ALU._0963_ ),
    .X(\u_cpu.ALU._1332_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU._2199_  (.A(\u_cpu.ALU._1330_ ),
    .B(\u_cpu.ALU._0738_ ),
    .C(\u_cpu.ALU._1331_ ),
    .D(\u_cpu.ALU._1332_ ),
    .X(\u_cpu.ALU._1333_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2200_  (.A1(\u_cpu.ALU._1158_ ),
    .A2(\u_cpu.ALU._1327_ ),
    .B1(\u_cpu.ALU._1333_ ),
    .Y(\u_cpu.ALU._1334_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU._2201_  (.A1(\u_cpu.ALU._1219_ ),
    .A2(\u_cpu.ALU._1279_ ),
    .A3(\u_cpu.ALU._0830_ ),
    .B1(\u_cpu.ALU._1317_ ),
    .Y(\u_cpu.ALU._1335_ ));
 sky130_fd_sc_hd__or4_2 \u_cpu.ALU._2202_  (.A(\u_cpu.ALU._1226_ ),
    .B(\u_cpu.ALU._0806_ ),
    .C(\u_cpu.ALU._1145_ ),
    .D(\u_cpu.ALU._0783_ ),
    .X(\u_cpu.ALU._1336_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.ALU._2203_  (.A1(\u_cpu.ALU._1149_ ),
    .A2(\u_cpu.ALU._0784_ ),
    .A3(\u_cpu.ALU._1335_ ),
    .B1(\u_cpu.ALU._1336_ ),
    .B2(\u_cpu.ALU._0876_ ),
    .X(\u_cpu.ALU._1337_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2204_  (.A(\u_cpu.ALU._0822_ ),
    .X(\u_cpu.ALU._1338_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2205_  (.A1(\u_cpu.ALU._1328_ ),
    .A2(\u_cpu.ALU._0658_ ),
    .B1(\u_cpu.ALU._1020_ ),
    .Y(\u_cpu.ALU._1339_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU._2206_  (.A1(\u_cpu.ALU._1328_ ),
    .A2(\u_cpu.ALU._0658_ ),
    .B1(\u_cpu.ALU._0749_ ),
    .B2(\u_cpu.ALU._1339_ ),
    .X(\u_cpu.ALU._1340_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._2207_  (.A1(\u_cpu.ALU._0957_ ),
    .A2(\u_cpu.ALU._1328_ ),
    .B1(\u_cpu.ALU._0658_ ),
    .C1(\u_cpu.ALU._0896_ ),
    .X(\u_cpu.ALU._1341_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU._2208_  (.A1(\u_cpu.ALU.Product_Wallace[13] ),
    .A2(\u_cpu.ALU._1338_ ),
    .B1(\u_cpu.ALU._1340_ ),
    .C1(\u_cpu.ALU._1341_ ),
    .Y(\u_cpu.ALU._1342_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2209_  (.A1(\u_cpu.ALU._1275_ ),
    .A2(\u_cpu.ALU._1337_ ),
    .B1(\u_cpu.ALU._1342_ ),
    .X(\u_cpu.ALU._1343_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU._2210_  (.A_N(\u_cpu.ALU._0660_ ),
    .B(\u_cpu.ALU._0800_ ),
    .C(\u_cpu.ALU._1232_ ),
    .D(\u_cpu.ALU._1293_ ),
    .Y(\u_cpu.ALU._1344_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU._2211_  (.A1(\u_cpu.ALU._0712_ ),
    .A2(\u_cpu.ALU._0710_ ),
    .A3(\u_cpu.ALU._1018_ ),
    .B1(\u_cpu.ALU._0658_ ),
    .C1(\u_cpu.ALU._1344_ ),
    .X(\u_cpu.ALU._1345_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2212_  (.A(\u_cpu.ALU._0985_ ),
    .X(\u_cpu.ALU._1346_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2213_  (.A1(\u_cpu.ALU._1346_ ),
    .A2(\u_cpu.ALU._1344_ ),
    .B1(\u_cpu.ALU._0658_ ),
    .Y(\u_cpu.ALU._1347_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2214_  (.A1(\u_cpu.ALU._1345_ ),
    .A2(\u_cpu.ALU._1347_ ),
    .B1(\u_cpu.ALU._1328_ ),
    .Y(\u_cpu.ALU._1348_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._2215_  (.A1(\u_cpu.ALU._0711_ ),
    .A2(\u_cpu.ALU._0920_ ),
    .B1(\u_cpu.ALU._0658_ ),
    .C1(\u_cpu.ALU._1344_ ),
    .Y(\u_cpu.ALU._1349_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2216_  (.A1(\u_cpu.ALU._0708_ ),
    .A2(\u_cpu.ALU._1018_ ),
    .B1(\u_cpu.ALU._0660_ ),
    .Y(\u_cpu.ALU._1350_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU._2217_  (.A_N(\u_cpu.ALU._0658_ ),
    .B(\u_cpu.ALU._1298_ ),
    .C(\u_cpu.ALU._1350_ ),
    .Y(\u_cpu.ALU._0000_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU._2218_  (.A_N(\u_cpu.ALU._1328_ ),
    .B(\u_cpu.ALU._1349_ ),
    .C(\u_cpu.ALU._0000_ ),
    .Y(\u_cpu.ALU._0001_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._2219_  (.A(\u_cpu.ALU._1348_ ),
    .B(\u_cpu.ALU._0001_ ),
    .X(\u_cpu.ALU._0002_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU._2220_  (.A1(\u_cpu.ALU._1295_ ),
    .A2(\u_cpu.ALU._1299_ ),
    .B1(\u_cpu.ALU._1303_ ),
    .B2(\u_cpu.ALU._1308_ ),
    .Y(\u_cpu.ALU._0003_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2221_  (.A1(\u_cpu.ALU._0003_ ),
    .A2(\u_cpu.ALU._0002_ ),
    .B1(\u_cpu.ALU._0921_ ),
    .Y(\u_cpu.ALU._0004_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2222_  (.A1(\u_cpu.ALU._0002_ ),
    .A2(\u_cpu.ALU._0003_ ),
    .B1(\u_cpu.ALU._0004_ ),
    .Y(\u_cpu.ALU._0005_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._2223_  (.A1(\u_cpu.ALU._1283_ ),
    .A2(\u_cpu.ALU._1334_ ),
    .B1(\u_cpu.ALU._1343_ ),
    .C1(\u_cpu.ALU._0005_ ),
    .Y(\u_cpu.ALU.ALUResult[13] ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2224_  (.A(\u_cpu.ALU.SrcB[13] ),
    .B(\u_cpu.ALU.SrcB[12] ),
    .Y(\u_cpu.ALU._0006_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU._2225_  (.A(\u_cpu.ALU._0800_ ),
    .B(\u_cpu.ALU._1232_ ),
    .C(\u_cpu.ALU._1293_ ),
    .D(\u_cpu.ALU._0006_ ),
    .Y(\u_cpu.ALU._0007_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU._2226_  (.A1(\u_cpu.ALU._0712_ ),
    .A2(\u_cpu.ALU._0710_ ),
    .A3(\u_cpu.ALU._1018_ ),
    .B1(\u_cpu.ALU._0654_ ),
    .C1(\u_cpu.ALU._0007_ ),
    .X(\u_cpu.ALU._0008_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2227_  (.A1(\u_cpu.ALU._1346_ ),
    .A2(\u_cpu.ALU._0007_ ),
    .B1(\u_cpu.ALU._0654_ ),
    .Y(\u_cpu.ALU._0009_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2228_  (.A1(\u_cpu.ALU._0008_ ),
    .A2(\u_cpu.ALU._0009_ ),
    .B1(\u_cpu.ALU._0679_ ),
    .Y(\u_cpu.ALU._0010_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._2229_  (.A1(\u_cpu.ALU._0711_ ),
    .A2(\u_cpu.ALU._0919_ ),
    .B1(\u_cpu.ALU._0654_ ),
    .C1(\u_cpu.ALU._0007_ ),
    .Y(\u_cpu.ALU._0011_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2230_  (.A1(\u_cpu.ALU._0985_ ),
    .A2(\u_cpu.ALU._0007_ ),
    .B1(\u_cpu.ALU._0654_ ),
    .X(\u_cpu.ALU._0012_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._2231_  (.A(\u_cpu.ALU._0680_ ),
    .B(\u_cpu.ALU._0011_ ),
    .C(\u_cpu.ALU._0012_ ),
    .Y(\u_cpu.ALU._0013_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._2232_  (.A(\u_cpu.ALU._0010_ ),
    .B(\u_cpu.ALU._0013_ ),
    .X(\u_cpu.ALU._0014_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU._2233_  (.A1(\u_cpu.ALU._1295_ ),
    .A2(\u_cpu.ALU._1299_ ),
    .B1(\u_cpu.ALU._1348_ ),
    .C1(\u_cpu.ALU._0001_ ),
    .D1(\u_cpu.ALU._1302_ ),
    .Y(\u_cpu.ALU._0015_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._2234_  (.A1(\u_cpu.ALU._1200_ ),
    .A2(\u_cpu.ALU._1294_ ),
    .B1(\u_cpu.ALU._0859_ ),
    .C1(\u_cpu.ALU._1300_ ),
    .X(\u_cpu.ALU._0016_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU._2235_  (.A1(\u_cpu.ALU._1349_ ),
    .A2(\u_cpu.ALU._0000_ ),
    .B1_N(\u_cpu.ALU._1328_ ),
    .Y(\u_cpu.ALU._0017_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2236_  (.A1(\u_cpu.ALU._0016_ ),
    .A2(\u_cpu.ALU._0017_ ),
    .B1(\u_cpu.ALU._0001_ ),
    .Y(\u_cpu.ALU._0018_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2237_  (.A1(\u_cpu.ALU._0015_ ),
    .A2(\u_cpu.ALU._1308_ ),
    .B1(\u_cpu.ALU._0018_ ),
    .Y(\u_cpu.ALU._0019_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2238_  (.A1(\u_cpu.ALU._0014_ ),
    .A2(\u_cpu.ALU._0019_ ),
    .B1(\u_cpu.ALU._0975_ ),
    .Y(\u_cpu.ALU._0020_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._2239_  (.A(\u_cpu.ALU._0019_ ),
    .B(\u_cpu.ALU._0010_ ),
    .C(\u_cpu.ALU._0013_ ),
    .X(\u_cpu.ALU._0021_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2240_  (.A0(\u_cpu.ALU._1116_ ),
    .A1(\u_cpu.ALU._0968_ ),
    .A2(\u_cpu.ALU._0949_ ),
    .A3(\u_cpu.ALU._1120_ ),
    .S0(\u_cpu.ALU._0806_ ),
    .S1(\u_cpu.ALU._1279_ ),
    .X(\u_cpu.ALU._0022_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2241_  (.A0(\u_cpu.ALU._0679_ ),
    .A1(\u_cpu.ALU._1328_ ),
    .A2(\u_cpu.ALU._0859_ ),
    .A3(\u_cpu.ALU._0686_ ),
    .S0(\u_cpu.ALU._0794_ ),
    .S1(\u_cpu.ALU._0729_ ),
    .X(\u_cpu.ALU._0023_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.ALU._2242_  (.A0(\u_cpu.ALU._1258_ ),
    .A1(\u_cpu.ALU._0023_ ),
    .S(\u_cpu.ALU._0769_ ),
    .X(\u_cpu.ALU._0024_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.ALU._2243_  (.A0(\u_cpu.ALU._1115_ ),
    .A1(\u_cpu.ALU._0024_ ),
    .S(\u_cpu.ALU._1219_ ),
    .X(\u_cpu.ALU._0025_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2244_  (.A(\u_cpu.ALU._1077_ ),
    .X(\u_cpu.ALU._0026_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU._2245_  (.A1(\u_cpu.ALU._0022_ ),
    .A2(\u_cpu.ALU._1158_ ),
    .B1(\u_cpu.ALU._0025_ ),
    .B2(\u_cpu.ALU._0026_ ),
    .Y(\u_cpu.ALU._0027_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2246_  (.A1(\u_cpu.ALU._0813_ ),
    .A2(\u_cpu.ALU._0656_ ),
    .B1(\u_cpu.ALU._0749_ ),
    .Y(\u_cpu.ALU._0028_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._2247_  (.A1(\u_cpu.ALU._0957_ ),
    .A2(\u_cpu.ALU._0679_ ),
    .B1(\u_cpu.ALU._0654_ ),
    .C1(\u_cpu.ALU._0896_ ),
    .X(\u_cpu.ALU._0029_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2248_  (.A1(\u_cpu.ALU.Product_Wallace[14] ),
    .A2(\u_cpu.ALU._1338_ ),
    .B1(\u_cpu.ALU._0029_ ),
    .Y(\u_cpu.ALU._0030_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU._2249_  (.A1(\u_cpu.ALU._1283_ ),
    .A2(\u_cpu.ALU._0027_ ),
    .B1(\u_cpu.ALU._0028_ ),
    .B2(\u_cpu.ALU._0655_ ),
    .C1(\u_cpu.ALU._0030_ ),
    .X(\u_cpu.ALU._0031_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2250_  (.A1(\u_cpu.ALU._0761_ ),
    .A2(\u_cpu.ALU._1145_ ),
    .B1(\u_cpu.ALU._0577_ ),
    .Y(\u_cpu.ALU._0032_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU._2251_  (.A1(\u_cpu.ALU._0761_ ),
    .A2(\u_cpu.ALU._1145_ ),
    .A3(\u_cpu.ALU._0967_ ),
    .B1(\u_cpu.ALU._0032_ ),
    .X(\u_cpu.ALU._0033_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.ALU._2252_  (.A1(\u_cpu.ALU._0899_ ),
    .A2(\u_cpu.ALU._0930_ ),
    .A3(\u_cpu.ALU._1336_ ),
    .B1(\u_cpu.ALU._0033_ ),
    .B2(\u_cpu.ALU._1125_ ),
    .X(\u_cpu.ALU._0034_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU._2253_  (.A(\u_cpu.ALU._1275_ ),
    .B(\u_cpu.ALU._0034_ ),
    .X(\u_cpu.ALU._0035_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._2254_  (.A1(\u_cpu.ALU._0020_ ),
    .A2(\u_cpu.ALU._0021_ ),
    .B1(\u_cpu.ALU._0031_ ),
    .C1(\u_cpu.ALU._0035_ ),
    .Y(\u_cpu.ALU.ALUResult[14] ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2255_  (.A(\u_cpu.ALU._0019_ ),
    .B(\u_cpu.ALU._0014_ ),
    .Y(\u_cpu.ALU._0036_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU._2256_  (.A(\u_cpu.ALU._0654_ ),
    .B(\u_cpu.ALU._0658_ ),
    .C(\u_cpu.ALU.SrcB[12] ),
    .Y(\u_cpu.ALU._0037_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU._2257_  (.A(\u_cpu.ALU._0800_ ),
    .B(\u_cpu.ALU._1232_ ),
    .C(\u_cpu.ALU._1293_ ),
    .D(\u_cpu.ALU._0037_ ),
    .Y(\u_cpu.ALU._0038_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU._2258_  (.A1(\u_cpu.ALU._0712_ ),
    .A2(\u_cpu.ALU._0710_ ),
    .A3(\u_cpu.ALU._1018_ ),
    .B1(\u_cpu.ALU.SrcB[15] ),
    .C1(\u_cpu.ALU._0038_ ),
    .X(\u_cpu.ALU._0039_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2259_  (.A1(\u_cpu.ALU._1346_ ),
    .A2(\u_cpu.ALU._0038_ ),
    .B1(\u_cpu.ALU.SrcB[15] ),
    .Y(\u_cpu.ALU._0040_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2260_  (.A1(\u_cpu.ALU._0039_ ),
    .A2(\u_cpu.ALU._0040_ ),
    .B1(\u_cpu.ALU._0948_ ),
    .Y(\u_cpu.ALU._0041_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._2261_  (.A1(\u_cpu.ALU._0710_ ),
    .A2(\u_cpu.ALU._0919_ ),
    .B1(\u_cpu.ALU.SrcB[15] ),
    .C1(\u_cpu.ALU._0038_ ),
    .Y(\u_cpu.ALU._0042_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._2262_  (.A(\u_cpu.ALU._0654_ ),
    .Y(\u_cpu.ALU._0043_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._2263_  (.A(\u_cpu.ALU.SrcB[15] ),
    .Y(\u_cpu.ALU._0044_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._2264_  (.A1(\u_cpu.ALU._0741_ ),
    .A2(\u_cpu.ALU._0811_ ),
    .A3(\u_cpu.ALU._0745_ ),
    .B1(\u_cpu.ALU._0006_ ),
    .X(\u_cpu.ALU._0045_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU._2265_  (.A1(\u_cpu.ALU._1200_ ),
    .A2(\u_cpu.ALU._0043_ ),
    .B1(\u_cpu.ALU._0044_ ),
    .C1(\u_cpu.ALU._0045_ ),
    .D1(\u_cpu.ALU._1298_ ),
    .Y(\u_cpu.ALU._0046_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._2266_  (.A(\u_cpu.ALU._0683_ ),
    .B(\u_cpu.ALU._0042_ ),
    .C(\u_cpu.ALU._0046_ ),
    .Y(\u_cpu.ALU._0047_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2267_  (.A(\u_cpu.ALU._0041_ ),
    .B(\u_cpu.ALU._0047_ ),
    .Y(\u_cpu.ALU._0048_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2268_  (.A1(\u_cpu.ALU._0010_ ),
    .A2(\u_cpu.ALU._0036_ ),
    .B1(\u_cpu.ALU._0048_ ),
    .Y(\u_cpu.ALU._0049_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._2269_  (.A1(\u_cpu.ALU._0010_ ),
    .A2(\u_cpu.ALU._0036_ ),
    .A3(\u_cpu.ALU._0048_ ),
    .B1(\u_cpu.ALU._0921_ ),
    .X(\u_cpu.ALU._0050_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2270_  (.A0(\u_cpu.ALU._0948_ ),
    .A1(\u_cpu.ALU._0679_ ),
    .A2(\u_cpu.ALU._1328_ ),
    .A3(\u_cpu.ALU._0859_ ),
    .S0(\u_cpu.ALU._0722_ ),
    .S1(\u_cpu.ALU._0729_ ),
    .X(\u_cpu.ALU._0051_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.ALU._2271_  (.A0(\u_cpu.ALU._1276_ ),
    .A1(\u_cpu.ALU._0051_ ),
    .S(\u_cpu.ALU._0769_ ),
    .X(\u_cpu.ALU._0052_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.ALU._2272_  (.A0(\u_cpu.ALU._1156_ ),
    .A1(\u_cpu.ALU._0052_ ),
    .S(\u_cpu.ALU._1219_ ),
    .X(\u_cpu.ALU._0053_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2273_  (.A0(\u_cpu.ALU._1146_ ),
    .A1(\u_cpu.ALU._1012_ ),
    .A2(\u_cpu.ALU._1284_ ),
    .A3(\u_cpu.ALU._1002_ ),
    .S0(\u_cpu.ALU._1076_ ),
    .S1(\u_cpu.ALU._1145_ ),
    .X(\u_cpu.ALU._0054_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU._2274_  (.A1(\u_cpu.ALU._0053_ ),
    .A2(\u_cpu.ALU._0026_ ),
    .B1(\u_cpu.ALU._1158_ ),
    .B2(\u_cpu.ALU._0054_ ),
    .X(\u_cpu.ALU._0055_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._2275_  (.A(\u_cpu.ALU._0881_ ),
    .B(\u_cpu.ALU.SrcA[31] ),
    .C(\u_cpu.ALU._1014_ ),
    .X(\u_cpu.ALU._0056_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._2276_  (.A1(\u_cpu.ALU._0577_ ),
    .A2(\u_cpu.ALU._0801_ ),
    .A3(\u_cpu.ALU._0882_ ),
    .B1(\u_cpu.ALU._0056_ ),
    .X(\u_cpu.ALU._0057_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2277_  (.A(\u_cpu.ALU._0744_ ),
    .X(\u_cpu.ALU._0058_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU._2278_  (.A1(\u_cpu.ALU._0948_ ),
    .A2(\u_cpu.ALU.SrcB[15] ),
    .A3(\u_cpu.ALU._0058_ ),
    .B1(\u_cpu.ALU._0822_ ),
    .B2(\u_cpu.ALU.Product_Wallace[15] ),
    .X(\u_cpu.ALU._0059_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2279_  (.A(\u_cpu.ALU._0754_ ),
    .X(\u_cpu.ALU._0060_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2280_  (.A(\u_cpu.ALU._0742_ ),
    .X(\u_cpu.ALU._0061_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2281_  (.A1(\u_cpu.ALU._0948_ ),
    .A2(\u_cpu.ALU.SrcB[15] ),
    .B1(\u_cpu.ALU._0061_ ),
    .C1(\u_cpu.ALU._1226_ ),
    .D1(\u_cpu.ALU._0963_ ),
    .X(\u_cpu.ALU._0062_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2282_  (.A1(\u_cpu.ALU.SrcB[15] ),
    .A2(\u_cpu.ALU._0060_ ),
    .B1(\u_cpu.ALU._0813_ ),
    .B2(\u_cpu.ALU._0653_ ),
    .C1(\u_cpu.ALU._0062_ ),
    .X(\u_cpu.ALU._0063_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._2283_  (.A1(\u_cpu.ALU._0057_ ),
    .A2(\u_cpu.ALU._1144_ ),
    .B1(\u_cpu.ALU._0059_ ),
    .C1(\u_cpu.ALU._0063_ ),
    .X(\u_cpu.ALU._0064_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2284_  (.A1(\u_cpu.ALU._1275_ ),
    .A2(\u_cpu.ALU._0055_ ),
    .B1(\u_cpu.ALU._0064_ ),
    .Y(\u_cpu.ALU._0065_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2285_  (.A1(\u_cpu.ALU._0049_ ),
    .A2(\u_cpu.ALU._0050_ ),
    .B1(\u_cpu.ALU._0065_ ),
    .Y(\u_cpu.ALU.ALUResult[15] ));
 sky130_fd_sc_hd__nor4_2 \u_cpu.ALU._2286_  (.A(\u_cpu.ALU.SrcB[15] ),
    .B(\u_cpu.ALU.SrcB[14] ),
    .C(\u_cpu.ALU.SrcB[13] ),
    .D(\u_cpu.ALU.SrcB[12] ),
    .Y(\u_cpu.ALU._0066_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU._2287_  (.A(\u_cpu.ALU._0800_ ),
    .B(\u_cpu.ALU._1232_ ),
    .C(\u_cpu.ALU._1293_ ),
    .D(\u_cpu.ALU._0066_ ),
    .Y(\u_cpu.ALU._0067_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2288_  (.A1(\u_cpu.ALU._0710_ ),
    .A2(\u_cpu.ALU._0919_ ),
    .B1(\u_cpu.ALU._0067_ ),
    .Y(\u_cpu.ALU._0068_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2289_  (.A(\u_cpu.ALU._0700_ ),
    .B(\u_cpu.ALU._0068_ ),
    .Y(\u_cpu.ALU._0069_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2290_  (.A(\u_cpu.ALU._0068_ ),
    .B(\u_cpu.ALU._0700_ ),
    .Y(\u_cpu.ALU._0070_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2291_  (.A(\u_cpu.ALU._0070_ ),
    .B(\u_cpu.ALU._0699_ ),
    .Y(\u_cpu.ALU._0071_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2292_  (.A(\u_cpu.ALU._0067_ ),
    .X(\u_cpu.ALU._0072_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU._2293_  (.A_N(\u_cpu.ALU._0700_ ),
    .B(\u_cpu.ALU._1346_ ),
    .C(\u_cpu.ALU._0072_ ),
    .Y(\u_cpu.ALU._0073_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2294_  (.A1(\u_cpu.ALU._0070_ ),
    .A2(\u_cpu.ALU._0073_ ),
    .B1(\u_cpu.ALU._0699_ ),
    .X(\u_cpu.ALU._0074_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2295_  (.A1(\u_cpu.ALU._0069_ ),
    .A2(\u_cpu.ALU._0071_ ),
    .B1(\u_cpu.ALU._0074_ ),
    .X(\u_cpu.ALU._0075_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU._2296_  (.A(\u_cpu.ALU._1230_ ),
    .B(\u_cpu.ALU._1272_ ),
    .C(\u_cpu.ALU._1236_ ),
    .D(\u_cpu.ALU._1239_ ),
    .Y(\u_cpu.ALU._0076_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2297_  (.A1(\u_cpu.ALU._1295_ ),
    .A2(\u_cpu.ALU._1299_ ),
    .B1(\u_cpu.ALU._1348_ ),
    .C1(\u_cpu.ALU._0001_ ),
    .D1(\u_cpu.ALU._1302_ ),
    .X(\u_cpu.ALU._0077_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU._2298_  (.A(\u_cpu.ALU._0010_ ),
    .B(\u_cpu.ALU._0013_ ),
    .C(\u_cpu.ALU._0041_ ),
    .D(\u_cpu.ALU._0047_ ),
    .X(\u_cpu.ALU._0078_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2299_  (.A(\u_cpu.ALU._0077_ ),
    .B(\u_cpu.ALU._0078_ ),
    .Y(\u_cpu.ALU._0079_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._2300_  (.A(\u_cpu.ALU._0683_ ),
    .B(\u_cpu.ALU._0042_ ),
    .C(\u_cpu.ALU._0046_ ),
    .X(\u_cpu.ALU._0080_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2301_  (.A(\u_cpu.ALU._0042_ ),
    .B(\u_cpu.ALU._0046_ ),
    .Y(\u_cpu.ALU._0081_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2302_  (.A(\u_cpu.ALU._0011_ ),
    .B(\u_cpu.ALU._0012_ ),
    .Y(\u_cpu.ALU._0082_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU._2303_  (.A1(\u_cpu.ALU._0081_ ),
    .A2(\u_cpu.ALU._0948_ ),
    .B1(\u_cpu.ALU._0082_ ),
    .B2(\u_cpu.ALU._0679_ ),
    .Y(\u_cpu.ALU._0083_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU._2304_  (.A(\u_cpu.ALU._0010_ ),
    .B(\u_cpu.ALU._0013_ ),
    .C(\u_cpu.ALU._0041_ ),
    .D(\u_cpu.ALU._0047_ ),
    .Y(\u_cpu.ALU._0084_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU._2305_  (.A1(\u_cpu.ALU._0080_ ),
    .A2(\u_cpu.ALU._0083_ ),
    .B1(\u_cpu.ALU._0084_ ),
    .B2(\u_cpu.ALU._0018_ ),
    .Y(\u_cpu.ALU._0085_ ));
 sky130_fd_sc_hd__a41oi_2 \u_cpu.ALU._2306_  (.A1(\u_cpu.ALU._1304_ ),
    .A2(\u_cpu.ALU._1306_ ),
    .A3(\u_cpu.ALU._0077_ ),
    .A4(\u_cpu.ALU._0078_ ),
    .B1(\u_cpu.ALU._0085_ ),
    .Y(\u_cpu.ALU._0086_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.ALU._2307_  (.A1(\u_cpu.ALU._0076_ ),
    .A2(\u_cpu.ALU._0079_ ),
    .A3(\u_cpu.ALU._1179_ ),
    .B1(\u_cpu.ALU._0086_ ),
    .Y(\u_cpu.ALU._0087_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2308_  (.A1(\u_cpu.ALU._0075_ ),
    .A2(\u_cpu.ALU._0087_ ),
    .B1(\u_cpu.ALU._0975_ ),
    .Y(\u_cpu.ALU._0088_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._2309_  (.A1(\u_cpu.ALU._0071_ ),
    .A2(\u_cpu.ALU._0069_ ),
    .B1(\u_cpu.ALU._0074_ ),
    .C1(\u_cpu.ALU._0087_ ),
    .X(\u_cpu.ALU._0089_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2310_  (.A0(\u_cpu.ALU._0699_ ),
    .A1(\u_cpu.ALU._0948_ ),
    .A2(\u_cpu.ALU._0679_ ),
    .A3(\u_cpu.ALU._1328_ ),
    .S0(\u_cpu.ALU._0794_ ),
    .S1(\u_cpu.ALU._0729_ ),
    .X(\u_cpu.ALU._0090_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2311_  (.A0(\u_cpu.ALU._1045_ ),
    .A1(\u_cpu.ALU._1194_ ),
    .A2(\u_cpu.ALU._1321_ ),
    .A3(\u_cpu.ALU._0090_ ),
    .S0(\u_cpu.ALU._0769_ ),
    .S1(\u_cpu.ALU._1088_ ),
    .X(\u_cpu.ALU._0091_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU._2312_  (.A1_N(\u_cpu.ALU._0026_ ),
    .A2_N(\u_cpu.ALU._0091_ ),
    .B1(\u_cpu.ALU._0784_ ),
    .B2(\u_cpu.ALU._0782_ ),
    .X(\u_cpu.ALU._0092_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._2313_  (.A1(\u_cpu.ALU.SrcA[0] ),
    .A2(\u_cpu.ALU._0801_ ),
    .A3(\u_cpu.ALU._1077_ ),
    .B1(\u_cpu.ALU._0056_ ),
    .X(\u_cpu.ALU._0093_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2314_  (.A1(\u_cpu.ALU._0699_ ),
    .A2(\u_cpu.ALU._0700_ ),
    .B1(\u_cpu.ALU._1020_ ),
    .Y(\u_cpu.ALU._0094_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU._2315_  (.A1(\u_cpu.ALU._0699_ ),
    .A2(\u_cpu.ALU._0700_ ),
    .B1(\u_cpu.ALU._0748_ ),
    .B2(\u_cpu.ALU._0094_ ),
    .X(\u_cpu.ALU._0095_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2316_  (.A1(\u_cpu.ALU._0702_ ),
    .A2(\u_cpu.ALU._0744_ ),
    .B1(\u_cpu.ALU._0821_ ),
    .B2(\u_cpu.ALU.Product_Wallace[16] ),
    .C1(\u_cpu.ALU._0095_ ),
    .X(\u_cpu.ALU._0096_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2317_  (.A1(\u_cpu.ALU._0700_ ),
    .A2(\u_cpu.ALU._0754_ ),
    .B1(\u_cpu.ALU._0093_ ),
    .B2(\u_cpu.ALU._0758_ ),
    .C1(\u_cpu.ALU._0096_ ),
    .X(\u_cpu.ALU._0097_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.ALU._2318_  (.A1(\u_cpu.ALU._1144_ ),
    .A2(\u_cpu.ALU._0092_ ),
    .B1_N(\u_cpu.ALU._0097_ ),
    .X(\u_cpu.ALU._0098_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2319_  (.A1(\u_cpu.ALU._0088_ ),
    .A2(\u_cpu.ALU._0089_ ),
    .B1(\u_cpu.ALU._0098_ ),
    .Y(\u_cpu.ALU.ALUResult[16] ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU._2320_  (.A1(\u_cpu.ALU._0710_ ),
    .A2(\u_cpu.ALU._0919_ ),
    .B1(\u_cpu.ALU._0700_ ),
    .B2(\u_cpu.ALU._0067_ ),
    .C1(\u_cpu.ALU._0537_ ),
    .X(\u_cpu.ALU._0099_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU._2321_  (.A1(\u_cpu.ALU._0750_ ),
    .A2(\u_cpu.ALU._0735_ ),
    .A3(\u_cpu.ALU._0708_ ),
    .B1(\u_cpu.ALU.SrcB[16] ),
    .X(\u_cpu.ALU._0100_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU._2322_  (.A1(\u_cpu.ALU._1346_ ),
    .A2(\u_cpu.ALU._0072_ ),
    .B1(\u_cpu.ALU._0100_ ),
    .C1(\u_cpu.ALU._0537_ ),
    .Y(\u_cpu.ALU._0101_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2323_  (.A1(\u_cpu.ALU._0099_ ),
    .A2(\u_cpu.ALU._0101_ ),
    .B1(\u_cpu.ALU._0536_ ),
    .Y(\u_cpu.ALU._0102_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2324_  (.A1(\u_cpu.ALU._1346_ ),
    .A2(\u_cpu.ALU._0067_ ),
    .B1(\u_cpu.ALU._0537_ ),
    .Y(\u_cpu.ALU._0103_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2325_  (.A1(\u_cpu.ALU._0708_ ),
    .A2(\u_cpu.ALU._1018_ ),
    .B1(\u_cpu.ALU._0700_ ),
    .Y(\u_cpu.ALU._0104_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._2326_  (.A1(\u_cpu.ALU._0103_ ),
    .A2(\u_cpu.ALU._0104_ ),
    .B1(\u_cpu.ALU._0536_ ),
    .C1(\u_cpu.ALU._0099_ ),
    .X(\u_cpu.ALU._0105_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._2327_  (.A(\u_cpu.ALU._0102_ ),
    .B(\u_cpu.ALU._0105_ ),
    .X(\u_cpu.ALU._0106_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU._2328_  (.A1_N(\u_cpu.ALU._0075_ ),
    .A2_N(\u_cpu.ALU._0087_ ),
    .B1(\u_cpu.ALU._0069_ ),
    .B2(\u_cpu.ALU._0071_ ),
    .Y(\u_cpu.ALU._0107_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2329_  (.A1(\u_cpu.ALU._0106_ ),
    .A2(\u_cpu.ALU._0107_ ),
    .B1(\u_cpu.ALU._0975_ ),
    .X(\u_cpu.ALU._0108_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2330_  (.A(\u_cpu.ALU._0107_ ),
    .B(\u_cpu.ALU._0106_ ),
    .Y(\u_cpu.ALU._0109_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2331_  (.A0(\u_cpu.ALU._0536_ ),
    .A1(\u_cpu.ALU._0699_ ),
    .A2(\u_cpu.ALU._0948_ ),
    .A3(\u_cpu.ALU._0679_ ),
    .S0(\u_cpu.ALU._0635_ ),
    .S1(\u_cpu.ALU._0726_ ),
    .X(\u_cpu.ALU._0110_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2332_  (.A0(\u_cpu.ALU._1078_ ),
    .A1(\u_cpu.ALU._1223_ ),
    .A2(\u_cpu.ALU._1329_ ),
    .A3(\u_cpu.ALU._0110_ ),
    .S0(\u_cpu.ALU._0785_ ),
    .S1(\u_cpu.ALU._0770_ ),
    .X(\u_cpu.ALU._0111_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU._2333_  (.A(\u_cpu.ALU._0758_ ),
    .B(\u_cpu.ALU._0111_ ),
    .X(\u_cpu.ALU._0112_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._2334_  (.A1(\u_cpu.ALU._1075_ ),
    .A2(\u_cpu.ALU._0894_ ),
    .B1(\u_cpu.ALU._0026_ ),
    .C1(\u_cpu.ALU._0112_ ),
    .X(\u_cpu.ALU._0113_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._2335_  (.A(\u_cpu.ALU._0613_ ),
    .B(\u_cpu.ALU._0577_ ),
    .C(\u_cpu.ALU._0874_ ),
    .X(\u_cpu.ALU._0114_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2336_  (.A(\u_cpu.ALU._0114_ ),
    .X(\u_cpu.ALU._0115_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._2337_  (.A1(\u_cpu.ALU._1075_ ),
    .A2(\u_cpu.ALU._0848_ ),
    .A3(\u_cpu.ALU._0874_ ),
    .B1(\u_cpu.ALU._0115_ ),
    .X(\u_cpu.ALU._0116_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2338_  (.A(\u_cpu.ALU._0539_ ),
    .B(\u_cpu.ALU._0540_ ),
    .Y(\u_cpu.ALU._0117_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2339_  (.A1(\u_cpu.ALU._0536_ ),
    .A2(\u_cpu.ALU._0537_ ),
    .B1(\u_cpu.ALU._0742_ ),
    .C1(\u_cpu.ALU._0881_ ),
    .D1(\u_cpu.ALU._0963_ ),
    .X(\u_cpu.ALU._0118_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2340_  (.A1(\u_cpu.ALU._0537_ ),
    .A2(\u_cpu.ALU._0754_ ),
    .B1(\u_cpu.ALU._0812_ ),
    .B2(\u_cpu.ALU._0117_ ),
    .C1(\u_cpu.ALU._0118_ ),
    .X(\u_cpu.ALU._0119_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2341_  (.A1(\u_cpu.ALU._0540_ ),
    .A2(\u_cpu.ALU._0058_ ),
    .B1(\u_cpu.ALU._0822_ ),
    .B2(\u_cpu.ALU.Product_Wallace[17] ),
    .C1(\u_cpu.ALU._0119_ ),
    .X(\u_cpu.ALU._0120_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._2342_  (.A1(\u_cpu.ALU._0847_ ),
    .A2(\u_cpu.ALU._0878_ ),
    .B1(\u_cpu.ALU._1124_ ),
    .C1(\u_cpu.ALU._0759_ ),
    .X(\u_cpu.ALU._0121_ ));
 sky130_fd_sc_hd__or4b_2 \u_cpu.ALU._2343_  (.A(\u_cpu.ALU._0113_ ),
    .B(\u_cpu.ALU._0116_ ),
    .C(\u_cpu.ALU._0120_ ),
    .D_N(\u_cpu.ALU._0121_ ),
    .X(\u_cpu.ALU._0122_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2344_  (.A1(\u_cpu.ALU._0108_ ),
    .A2(\u_cpu.ALU._0109_ ),
    .B1(\u_cpu.ALU._0122_ ),
    .Y(\u_cpu.ALU._0123_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._2345_  (.A(\u_cpu.ALU._0123_ ),
    .Y(\u_cpu.ALU.ALUResult[17] ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2346_  (.A1(\u_cpu.ALU._0069_ ),
    .A2(\u_cpu.ALU._0071_ ),
    .B1(\u_cpu.ALU._0102_ ),
    .Y(\u_cpu.ALU._0124_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2347_  (.A(\u_cpu.ALU._0105_ ),
    .B(\u_cpu.ALU._0124_ ),
    .Y(\u_cpu.ALU._0125_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2348_  (.A1(\u_cpu.ALU._0071_ ),
    .A2(\u_cpu.ALU._0069_ ),
    .B1(\u_cpu.ALU._0074_ ),
    .C1(\u_cpu.ALU._0102_ ),
    .D1(\u_cpu.ALU._0105_ ),
    .X(\u_cpu.ALU._0126_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2349_  (.A(\u_cpu.ALU._0087_ ),
    .B(\u_cpu.ALU._0126_ ),
    .Y(\u_cpu.ALU._0127_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2350_  (.A(\u_cpu.ALU._1165_ ),
    .B(\u_cpu.ALU._1297_ ),
    .Y(\u_cpu.ALU._0128_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2351_  (.A(\u_cpu.ALU.SrcB[17] ),
    .B(\u_cpu.ALU.SrcB[16] ),
    .Y(\u_cpu.ALU._0129_ ));
 sky130_fd_sc_hd__a311o_2 \u_cpu.ALU._2352_  (.A1(\u_cpu.ALU._0128_ ),
    .A2(\u_cpu.ALU._0066_ ),
    .A3(\u_cpu.ALU._0129_ ),
    .B1(\u_cpu.ALU._1200_ ),
    .C1(\u_cpu.ALU._0534_ ),
    .X(\u_cpu.ALU._0130_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._2353_  (.A1(\u_cpu.ALU._1200_ ),
    .A2(\u_cpu.ALU._0129_ ),
    .B1(\u_cpu.ALU._0534_ ),
    .C1(\u_cpu.ALU._0068_ ),
    .Y(\u_cpu.ALU._0131_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._2354_  (.A(\u_cpu.ALU._0130_ ),
    .B(\u_cpu.ALU._0131_ ),
    .C(\u_cpu.ALU._0533_ ),
    .Y(\u_cpu.ALU._0132_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2355_  (.A1(\u_cpu.ALU._0130_ ),
    .A2(\u_cpu.ALU._0131_ ),
    .B1(\u_cpu.ALU._0533_ ),
    .X(\u_cpu.ALU._0133_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2356_  (.A(\u_cpu.ALU._0132_ ),
    .B(\u_cpu.ALU._0133_ ),
    .Y(\u_cpu.ALU._0134_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2357_  (.A1(\u_cpu.ALU._0125_ ),
    .A2(\u_cpu.ALU._0127_ ),
    .B1(\u_cpu.ALU._0134_ ),
    .X(\u_cpu.ALU._0135_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._2358_  (.A(\u_cpu.ALU._0544_ ),
    .B(\u_cpu.ALU._0130_ ),
    .C(\u_cpu.ALU._0131_ ),
    .Y(\u_cpu.ALU._0136_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU._2359_  (.A(\u_cpu.ALU._0537_ ),
    .B(\u_cpu.ALU.SrcB[16] ),
    .X(\u_cpu.ALU._0137_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU._2360_  (.A1(\u_cpu.ALU._0711_ ),
    .A2(\u_cpu.ALU._0920_ ),
    .B1(\u_cpu.ALU._0072_ ),
    .B2(\u_cpu.ALU._0137_ ),
    .C1(\u_cpu.ALU._0534_ ),
    .X(\u_cpu.ALU._0138_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._2361_  (.A1(\u_cpu.ALU._0741_ ),
    .A2(\u_cpu.ALU._0811_ ),
    .A3(\u_cpu.ALU._0746_ ),
    .B1(\u_cpu.ALU._0129_ ),
    .X(\u_cpu.ALU._0139_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU._2362_  (.A_N(\u_cpu.ALU._0534_ ),
    .B(\u_cpu.ALU._0068_ ),
    .C(\u_cpu.ALU._0139_ ),
    .Y(\u_cpu.ALU._0140_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU._2363_  (.A_N(\u_cpu.ALU._0138_ ),
    .B(\u_cpu.ALU._0140_ ),
    .C(\u_cpu.ALU._0533_ ),
    .Y(\u_cpu.ALU._0141_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2364_  (.A(\u_cpu.ALU._0136_ ),
    .B(\u_cpu.ALU._0141_ ),
    .Y(\u_cpu.ALU._0142_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2365_  (.A1(\u_cpu.ALU._0105_ ),
    .A2(\u_cpu.ALU._0124_ ),
    .B1(\u_cpu.ALU._0087_ ),
    .B2(\u_cpu.ALU._0126_ ),
    .C1(\u_cpu.ALU._0142_ ),
    .X(\u_cpu.ALU._0143_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2366_  (.A(\u_cpu.ALU._0975_ ),
    .X(\u_cpu.ALU._0144_ ));
 sky130_fd_sc_hd__nor4_2 \u_cpu.ALU._2367_  (.A(\u_cpu.ALU._1331_ ),
    .B(\u_cpu.ALU._1144_ ),
    .C(\u_cpu.ALU._0784_ ),
    .D(\u_cpu.ALU._0942_ ),
    .Y(\u_cpu.ALU._0145_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2368_  (.A1(\u_cpu.ALU._0533_ ),
    .A2(\u_cpu.ALU._0534_ ),
    .B1(\u_cpu.ALU._0061_ ),
    .C1(\u_cpu.ALU._1226_ ),
    .D1(\u_cpu.ALU._0963_ ),
    .X(\u_cpu.ALU._0146_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU._2369_  (.A1(\u_cpu.ALU._0533_ ),
    .A2(\u_cpu.ALU._0534_ ),
    .A3(\u_cpu.ALU._0744_ ),
    .B1(\u_cpu.ALU._0821_ ),
    .B2(\u_cpu.ALU.Product_Wallace[18] ),
    .X(\u_cpu.ALU._0147_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.ALU._2370_  (.A_N(\u_cpu.ALU._0535_ ),
    .B(\u_cpu.ALU._0738_ ),
    .C(\u_cpu.ALU._0890_ ),
    .D(\u_cpu.ALU._1149_ ),
    .X(\u_cpu.ALU._0148_ ));
 sky130_fd_sc_hd__a2111o_2 \u_cpu.ALU._2371_  (.A1(\u_cpu.ALU._0534_ ),
    .A2(\u_cpu.ALU._0060_ ),
    .B1(\u_cpu.ALU._0146_ ),
    .C1(\u_cpu.ALU._0147_ ),
    .D1(\u_cpu.ALU._0148_ ),
    .X(\u_cpu.ALU._0149_ ));
 sky130_fd_sc_hd__or4_2 \u_cpu.ALU._2372_  (.A(\u_cpu.ALU._1149_ ),
    .B(\u_cpu.ALU._0879_ ),
    .C(\u_cpu.ALU._0994_ ),
    .D(\u_cpu.ALU._0784_ ),
    .X(\u_cpu.ALU._0150_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2373_  (.A0(\u_cpu.ALU._0533_ ),
    .A1(\u_cpu.ALU._0536_ ),
    .A2(\u_cpu.ALU._0699_ ),
    .A3(\u_cpu.ALU._0948_ ),
    .S0(\u_cpu.ALU._0794_ ),
    .S1(\u_cpu.ALU._0729_ ),
    .X(\u_cpu.ALU._0151_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2374_  (.A0(\u_cpu.ALU._0023_ ),
    .A1(\u_cpu.ALU._1114_ ),
    .A2(\u_cpu.ALU._0151_ ),
    .A3(\u_cpu.ALU._1258_ ),
    .S0(\u_cpu.ALU._0760_ ),
    .S1(\u_cpu.ALU._0786_ ),
    .X(\u_cpu.ALU._0152_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._2375_  (.A1(\u_cpu.ALU._0962_ ),
    .A2(\u_cpu.ALU._0786_ ),
    .A3(\u_cpu.ALU._1088_ ),
    .B1(\u_cpu.ALU._0879_ ),
    .X(\u_cpu.ALU._0153_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._2376_  (.A1(\u_cpu.ALU._0758_ ),
    .A2(\u_cpu.ALU._0152_ ),
    .B1(\u_cpu.ALU._0153_ ),
    .C1(\u_cpu.ALU._0026_ ),
    .Y(\u_cpu.ALU._0154_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU._2377_  (.A1(\u_cpu.ALU._0759_ ),
    .A2(\u_cpu.ALU._1125_ ),
    .A3(\u_cpu.ALU._0971_ ),
    .B1(\u_cpu.ALU._0150_ ),
    .C1(\u_cpu.ALU._0154_ ),
    .X(\u_cpu.ALU._0155_ ));
 sky130_fd_sc_hd__or3b_2 \u_cpu.ALU._2378_  (.A(\u_cpu.ALU._0145_ ),
    .B(\u_cpu.ALU._0149_ ),
    .C_N(\u_cpu.ALU._0155_ ),
    .X(\u_cpu.ALU._0156_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU._2379_  (.A1(\u_cpu.ALU._0135_ ),
    .A2(\u_cpu.ALU._0143_ ),
    .A3(\u_cpu.ALU._0144_ ),
    .B1(\u_cpu.ALU._0156_ ),
    .Y(\u_cpu.ALU._0157_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._2380_  (.A(\u_cpu.ALU._0157_ ),
    .Y(\u_cpu.ALU.ALUResult[18] ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU._2381_  (.A1(\u_cpu.ALU._0105_ ),
    .A2(\u_cpu.ALU._0124_ ),
    .B1(\u_cpu.ALU._0087_ ),
    .B2(\u_cpu.ALU._0126_ ),
    .Y(\u_cpu.ALU._0158_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2382_  (.A1(\u_cpu.ALU._0134_ ),
    .A2(\u_cpu.ALU._0158_ ),
    .B1(\u_cpu.ALU._0132_ ),
    .Y(\u_cpu.ALU._0159_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2383_  (.A(\u_cpu.ALU._1346_ ),
    .X(\u_cpu.ALU._0160_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU._2384_  (.A1(\u_cpu.ALU._0137_ ),
    .A2(\u_cpu.ALU._0534_ ),
    .A3(\u_cpu.ALU._0072_ ),
    .B1(\u_cpu.ALU._0160_ ),
    .C1(\u_cpu.ALU.SrcB[19] ),
    .X(\u_cpu.ALU._0161_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2385_  (.A(\u_cpu.ALU._0547_ ),
    .B(\u_cpu.ALU._0161_ ),
    .Y(\u_cpu.ALU._0162_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2386_  (.A1(\u_cpu.ALU._0708_ ),
    .A2(\u_cpu.ALU._1018_ ),
    .B1(\u_cpu.ALU.SrcB[18] ),
    .Y(\u_cpu.ALU._0163_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU._2387_  (.A_N(\u_cpu.ALU.SrcB[19] ),
    .B(\u_cpu.ALU._0068_ ),
    .C(\u_cpu.ALU._0139_ ),
    .D(\u_cpu.ALU._0163_ ),
    .Y(\u_cpu.ALU._0164_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.ALU._2388_  (.A1(\u_cpu.ALU._0137_ ),
    .A2(\u_cpu.ALU.SrcB[18] ),
    .A3(\u_cpu.ALU._0072_ ),
    .B1(\u_cpu.ALU._1346_ ),
    .C1(\u_cpu.ALU.SrcB[19] ),
    .Y(\u_cpu.ALU._0165_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU._2389_  (.A1(\u_cpu.ALU._0165_ ),
    .A2(\u_cpu.ALU._0164_ ),
    .B1_N(\u_cpu.ALU._0547_ ),
    .Y(\u_cpu.ALU._0166_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2390_  (.A1(\u_cpu.ALU._0162_ ),
    .A2(\u_cpu.ALU._0164_ ),
    .B1(\u_cpu.ALU._0166_ ),
    .Y(\u_cpu.ALU._0167_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2391_  (.A(\u_cpu.ALU._0159_ ),
    .B(\u_cpu.ALU._0167_ ),
    .Y(\u_cpu.ALU._0168_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2392_  (.A1(\u_cpu.ALU._0162_ ),
    .A2(\u_cpu.ALU._0164_ ),
    .B1(\u_cpu.ALU._0166_ ),
    .X(\u_cpu.ALU._0169_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._2393_  (.A1(\u_cpu.ALU._0134_ ),
    .A2(\u_cpu.ALU._0158_ ),
    .B1(\u_cpu.ALU._0132_ ),
    .C1(\u_cpu.ALU._0169_ ),
    .Y(\u_cpu.ALU._0170_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._2394_  (.A(\u_cpu.ALU._0547_ ),
    .B(\u_cpu.ALU.SrcB[19] ),
    .C(\u_cpu.ALU._0744_ ),
    .X(\u_cpu.ALU._0171_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2395_  (.A1(\u_cpu.ALU._0530_ ),
    .A2(\u_cpu.ALU._0749_ ),
    .B1(\u_cpu.ALU._0822_ ),
    .B2(\u_cpu.ALU.Product_Wallace[19] ),
    .C1(\u_cpu.ALU._0171_ ),
    .X(\u_cpu.ALU._0172_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2396_  (.A1(\u_cpu.ALU.SrcB[19] ),
    .A2(\u_cpu.ALU._0060_ ),
    .B1(\u_cpu.ALU._0813_ ),
    .B2(\u_cpu.ALU._0532_ ),
    .C1(\u_cpu.ALU._0115_ ),
    .X(\u_cpu.ALU._0173_ ));
 sky130_fd_sc_hd__a21bo_2 \u_cpu.ALU._2397_  (.A1(\u_cpu.ALU._1285_ ),
    .A2(\u_cpu.ALU._0761_ ),
    .B1_N(\u_cpu.ALU._1004_ ),
    .X(\u_cpu.ALU._0174_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2398_  (.A1(\u_cpu.ALU._1331_ ),
    .A2(\u_cpu.ALU._1006_ ),
    .B1(\u_cpu.ALU._1158_ ),
    .C1(\u_cpu.ALU._1075_ ),
    .D1(\u_cpu.ALU._0174_ ),
    .X(\u_cpu.ALU._0175_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2399_  (.A0(\u_cpu.ALU._0547_ ),
    .A1(\u_cpu.ALU._0533_ ),
    .A2(\u_cpu.ALU._0536_ ),
    .A3(\u_cpu.ALU._0699_ ),
    .S0(\u_cpu.ALU._0722_ ),
    .S1(\u_cpu.ALU._0790_ ),
    .X(\u_cpu.ALU._0176_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2400_  (.A0(\u_cpu.ALU._1155_ ),
    .A1(\u_cpu.ALU._1276_ ),
    .A2(\u_cpu.ALU._0051_ ),
    .A3(\u_cpu.ALU._0176_ ),
    .S0(\u_cpu.ALU._0786_ ),
    .S1(\u_cpu.ALU._1076_ ),
    .X(\u_cpu.ALU._0177_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._2401_  (.A1(\u_cpu.ALU._1219_ ),
    .A2(\u_cpu.ALU._1279_ ),
    .A3(\u_cpu.ALU._1017_ ),
    .B1(\u_cpu.ALU._0879_ ),
    .X(\u_cpu.ALU._0178_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._2402_  (.A1(\u_cpu.ALU._0759_ ),
    .A2(\u_cpu.ALU._0177_ ),
    .B1(\u_cpu.ALU._0178_ ),
    .C1(\u_cpu.ALU._0026_ ),
    .X(\u_cpu.ALU._0179_ ));
 sky130_fd_sc_hd__or4_2 \u_cpu.ALU._2403_  (.A(\u_cpu.ALU._0172_ ),
    .B(\u_cpu.ALU._0173_ ),
    .C(\u_cpu.ALU._0175_ ),
    .D(\u_cpu.ALU._0179_ ),
    .X(\u_cpu.ALU._0180_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._2404_  (.A1(\u_cpu.ALU._0168_ ),
    .A2(\u_cpu.ALU._0144_ ),
    .A3(\u_cpu.ALU._0170_ ),
    .B1(\u_cpu.ALU._0180_ ),
    .X(\u_cpu.ALU.ALUResult[19] ));
 sky130_fd_sc_hd__a21bo_2 \u_cpu.ALU._2405_  (.A1(\u_cpu.ALU._0165_ ),
    .A2(\u_cpu.ALU._0164_ ),
    .B1_N(\u_cpu.ALU._0547_ ),
    .X(\u_cpu.ALU._0181_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU._2406_  (.A_N(\u_cpu.ALU._0547_ ),
    .B(\u_cpu.ALU._0165_ ),
    .C(\u_cpu.ALU._0164_ ),
    .Y(\u_cpu.ALU._0182_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU._2407_  (.A(\u_cpu.ALU._0126_ ),
    .B(\u_cpu.ALU._0142_ ),
    .C(\u_cpu.ALU._0181_ ),
    .D(\u_cpu.ALU._0182_ ),
    .Y(\u_cpu.ALU._0183_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._2408_  (.A(\u_cpu.ALU._0183_ ),
    .Y(\u_cpu.ALU._0184_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU._2409_  (.A(\u_cpu.ALU._0132_ ),
    .B(\u_cpu.ALU._0133_ ),
    .C(\u_cpu.ALU._0181_ ),
    .D(\u_cpu.ALU._0182_ ),
    .X(\u_cpu.ALU._0185_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU._2410_  (.A1(\u_cpu.ALU._0164_ ),
    .A2(\u_cpu.ALU._0162_ ),
    .B1(\u_cpu.ALU._0181_ ),
    .B2(\u_cpu.ALU._0132_ ),
    .Y(\u_cpu.ALU._0186_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._2411_  (.A1(\u_cpu.ALU._0185_ ),
    .A2(\u_cpu.ALU._0124_ ),
    .A3(\u_cpu.ALU._0105_ ),
    .B1(\u_cpu.ALU._0186_ ),
    .X(\u_cpu.ALU._0187_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2412_  (.A1(\u_cpu.ALU._0087_ ),
    .A2(\u_cpu.ALU._0184_ ),
    .B1(\u_cpu.ALU._0187_ ),
    .Y(\u_cpu.ALU._0188_ ));
 sky130_fd_sc_hd__or4_2 \u_cpu.ALU._2413_  (.A(\u_cpu.ALU.SrcB[19] ),
    .B(\u_cpu.ALU.SrcB[18] ),
    .C(\u_cpu.ALU._0537_ ),
    .D(\u_cpu.ALU.SrcB[16] ),
    .X(\u_cpu.ALU._0189_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._2414_  (.A(\u_cpu.ALU.SrcB[20] ),
    .Y(\u_cpu.ALU._0190_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU._2415_  (.A1(\u_cpu.ALU._0873_ ),
    .A2(\u_cpu.ALU._0920_ ),
    .B1(\u_cpu.ALU._0072_ ),
    .B2(\u_cpu.ALU._0189_ ),
    .C1(\u_cpu.ALU._0190_ ),
    .X(\u_cpu.ALU._0191_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2416_  (.A1(\u_cpu.ALU._0067_ ),
    .A2(\u_cpu.ALU._0189_ ),
    .B1(\u_cpu.ALU._0985_ ),
    .Y(\u_cpu.ALU._0192_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2417_  (.A1(\u_cpu.ALU._0192_ ),
    .A2(\u_cpu.ALU._0557_ ),
    .B1(\u_cpu.ALU._0570_ ),
    .X(\u_cpu.ALU._0193_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2418_  (.A(\u_cpu.ALU._0192_ ),
    .B(\u_cpu.ALU._0557_ ),
    .Y(\u_cpu.ALU._0194_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU._2419_  (.A1(\u_cpu.ALU._0711_ ),
    .A2(\u_cpu.ALU._0920_ ),
    .B1(\u_cpu.ALU._0072_ ),
    .B2(\u_cpu.ALU._0189_ ),
    .C1(\u_cpu.ALU._0190_ ),
    .Y(\u_cpu.ALU._0195_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2420_  (.A1(\u_cpu.ALU._0194_ ),
    .A2(\u_cpu.ALU._0195_ ),
    .B1(\u_cpu.ALU._0837_ ),
    .X(\u_cpu.ALU._0196_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2421_  (.A1(\u_cpu.ALU._0191_ ),
    .A2(\u_cpu.ALU._0193_ ),
    .B1(\u_cpu.ALU._0196_ ),
    .Y(\u_cpu.ALU._0197_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2422_  (.A1(\u_cpu.ALU._0192_ ),
    .A2(\u_cpu.ALU._0557_ ),
    .B1(\u_cpu.ALU._0570_ ),
    .Y(\u_cpu.ALU._0198_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2423_  (.A1(\u_cpu.ALU._0557_ ),
    .A2(\u_cpu.ALU._0192_ ),
    .B1(\u_cpu.ALU._0198_ ),
    .Y(\u_cpu.ALU._0199_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2424_  (.A1(\u_cpu.ALU._0196_ ),
    .A2(\u_cpu.ALU._0199_ ),
    .B1(\u_cpu.ALU._0087_ ),
    .B2(\u_cpu.ALU._0184_ ),
    .C1(\u_cpu.ALU._0187_ ),
    .X(\u_cpu.ALU._0200_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU._2425_  (.A1(\u_cpu.ALU._0188_ ),
    .A2(\u_cpu.ALU._0197_ ),
    .B1(\u_cpu.ALU._0061_ ),
    .C1(\u_cpu.ALU._0890_ ),
    .D1(\u_cpu.ALU._0200_ ),
    .Y(\u_cpu.ALU._0201_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2426_  (.A0(\u_cpu.ALU._0837_ ),
    .A1(\u_cpu.ALU._0547_ ),
    .A2(\u_cpu.ALU._0533_ ),
    .A3(\u_cpu.ALU._0536_ ),
    .S0(\u_cpu.ALU._0722_ ),
    .S1(\u_cpu.ALU._0790_ ),
    .X(\u_cpu.ALU._0202_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2427_  (.A0(\u_cpu.ALU._1194_ ),
    .A1(\u_cpu.ALU._1321_ ),
    .A2(\u_cpu.ALU._0090_ ),
    .A3(\u_cpu.ALU._0202_ ),
    .S0(\u_cpu.ALU._0786_ ),
    .S1(\u_cpu.ALU._1076_ ),
    .X(\u_cpu.ALU._0203_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2428_  (.A1(\u_cpu.ALU._1056_ ),
    .A2(\u_cpu.ALU._1059_ ),
    .B1(\u_cpu.ALU._0784_ ),
    .Y(\u_cpu.ALU._0204_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2429_  (.A1(\u_cpu.ALU._0026_ ),
    .A2(\u_cpu.ALU._0203_ ),
    .B1(\u_cpu.ALU._0204_ ),
    .X(\u_cpu.ALU._0205_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2430_  (.A1(\u_cpu.ALU._1145_ ),
    .A2(\u_cpu.ALU._1045_ ),
    .B1(\u_cpu.ALU._1046_ ),
    .C1(\u_cpu.ALU._1047_ ),
    .D1(\u_cpu.ALU._0759_ ),
    .X(\u_cpu.ALU._0206_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU._2431_  (.A1(\u_cpu.ALU._0837_ ),
    .A2(\u_cpu.ALU._0557_ ),
    .A3(\u_cpu.ALU._0744_ ),
    .B1(\u_cpu.ALU._0821_ ),
    .B2(\u_cpu.ALU.Product_Wallace[20] ),
    .X(\u_cpu.ALU._0207_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._2432_  (.A(\u_cpu.ALU._0812_ ),
    .B(\u_cpu.ALU._0559_ ),
    .C(\u_cpu.ALU._0558_ ),
    .X(\u_cpu.ALU._0208_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU._2433_  (.A1(\u_cpu.ALU._0557_ ),
    .A2(\u_cpu.ALU._0754_ ),
    .B1(\u_cpu.ALU._0748_ ),
    .B2(\u_cpu.ALU._0559_ ),
    .X(\u_cpu.ALU._0209_ ));
 sky130_fd_sc_hd__or4_2 \u_cpu.ALU._2434_  (.A(\u_cpu.ALU._0207_ ),
    .B(\u_cpu.ALU._0208_ ),
    .C(\u_cpu.ALU._0209_ ),
    .D(\u_cpu.ALU._0115_ ),
    .X(\u_cpu.ALU._0210_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._2435_  (.A1(\u_cpu.ALU._1275_ ),
    .A2(\u_cpu.ALU._0205_ ),
    .B1(\u_cpu.ALU._0206_ ),
    .C1(\u_cpu.ALU._0210_ ),
    .X(\u_cpu.ALU._0211_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._2436_  (.A(\u_cpu.ALU._0211_ ),
    .Y(\u_cpu.ALU._0212_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2437_  (.A(\u_cpu.ALU._0201_ ),
    .B(\u_cpu.ALU._0212_ ),
    .Y(\u_cpu.ALU.ALUResult[20] ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.ALU._2438_  (.A1(\u_cpu.ALU._0557_ ),
    .A2(\u_cpu.ALU._0067_ ),
    .A3(\u_cpu.ALU._0189_ ),
    .B1(\u_cpu.ALU._1346_ ),
    .C1(\u_cpu.ALU.SrcB[21] ),
    .Y(\u_cpu.ALU._0213_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._2439_  (.A1(\u_cpu.ALU._1200_ ),
    .A2(\u_cpu.ALU._0190_ ),
    .B1(\u_cpu.ALU._0568_ ),
    .C1(\u_cpu.ALU._0192_ ),
    .Y(\u_cpu.ALU._0214_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2440_  (.A(\u_cpu.ALU._0213_ ),
    .B(\u_cpu.ALU._0214_ ),
    .Y(\u_cpu.ALU._0215_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2441_  (.A(\u_cpu.ALU.SrcA[21] ),
    .X(\u_cpu.ALU._0216_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2442_  (.A(\u_cpu.ALU._0215_ ),
    .B(\u_cpu.ALU._0216_ ),
    .Y(\u_cpu.ALU._0217_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU._2443_  (.A_N(\u_cpu.ALU._0216_ ),
    .B(\u_cpu.ALU._0213_ ),
    .C(\u_cpu.ALU._0214_ ),
    .Y(\u_cpu.ALU._0218_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2444_  (.A1(\u_cpu.ALU._0194_ ),
    .A2(\u_cpu.ALU._0195_ ),
    .B1(\u_cpu.ALU._0837_ ),
    .Y(\u_cpu.ALU._0219_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2445_  (.A1(\u_cpu.ALU._0219_ ),
    .A2(\u_cpu.ALU._0188_ ),
    .B1(\u_cpu.ALU._0199_ ),
    .Y(\u_cpu.ALU._0220_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._2446_  (.A(\u_cpu.ALU._0217_ ),
    .B(\u_cpu.ALU._0218_ ),
    .C(\u_cpu.ALU._0220_ ),
    .Y(\u_cpu.ALU._0221_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2447_  (.A(\u_cpu.ALU._0217_ ),
    .B(\u_cpu.ALU._0218_ ),
    .Y(\u_cpu.ALU._0222_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._2448_  (.A1(\u_cpu.ALU._0197_ ),
    .A2(\u_cpu.ALU._0188_ ),
    .B1(\u_cpu.ALU._0222_ ),
    .C1(\u_cpu.ALU._0199_ ),
    .Y(\u_cpu.ALU._0223_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2449_  (.A(\u_cpu.ALU._0550_ ),
    .B(\u_cpu.ALU._0551_ ),
    .Y(\u_cpu.ALU._0224_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2450_  (.A1(\u_cpu.ALU._0216_ ),
    .A2(\u_cpu.ALU.SrcB[21] ),
    .B1(\u_cpu.ALU._0742_ ),
    .C1(\u_cpu.ALU._1226_ ),
    .D1(\u_cpu.ALU._0963_ ),
    .X(\u_cpu.ALU._0225_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2451_  (.A1(\u_cpu.ALU.SrcB[21] ),
    .A2(\u_cpu.ALU._0060_ ),
    .B1(\u_cpu.ALU._0225_ ),
    .X(\u_cpu.ALU._0226_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2452_  (.A1(\u_cpu.ALU._0550_ ),
    .A2(\u_cpu.ALU._0744_ ),
    .B1(\u_cpu.ALU._0822_ ),
    .B2(\u_cpu.ALU.Product_Wallace[21] ),
    .C1(\u_cpu.ALU._0114_ ),
    .X(\u_cpu.ALU._0227_ ));
 sky130_fd_sc_hd__or4b_2 \u_cpu.ALU._2453_  (.A(\u_cpu.ALU._0890_ ),
    .B(\u_cpu.ALU._0900_ ),
    .C(\u_cpu.ALU._0757_ ),
    .D_N(\u_cpu.ALU._0737_ ),
    .X(\u_cpu.ALU._0228_ ));
 sky130_fd_sc_hd__or3b_2 \u_cpu.ALU._2454_  (.A(\u_cpu.ALU._0806_ ),
    .B(\u_cpu.ALU._1257_ ),
    .C_N(\u_cpu.ALU._1079_ ),
    .X(\u_cpu.ALU._0229_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2455_  (.A0(\u_cpu.ALU._0216_ ),
    .A1(\u_cpu.ALU._0837_ ),
    .A2(\u_cpu.ALU._0547_ ),
    .A3(\u_cpu.ALU._0533_ ),
    .S0(\u_cpu.ALU._0722_ ),
    .S1(\u_cpu.ALU._0790_ ),
    .X(\u_cpu.ALU._0230_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2456_  (.A0(\u_cpu.ALU._1223_ ),
    .A1(\u_cpu.ALU._1329_ ),
    .A2(\u_cpu.ALU._0110_ ),
    .A3(\u_cpu.ALU._0230_ ),
    .S0(\u_cpu.ALU._0769_ ),
    .S1(\u_cpu.ALU._1088_ ),
    .X(\u_cpu.ALU._0231_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU._2457_  (.A1_N(\u_cpu.ALU._0228_ ),
    .A2_N(\u_cpu.ALU._0229_ ),
    .B1(\u_cpu.ALU._0231_ ),
    .B2(\u_cpu.ALU._0759_ ),
    .X(\u_cpu.ALU._0232_ ));
 sky130_fd_sc_hd__a2111o_2 \u_cpu.ALU._2458_  (.A1(\u_cpu.ALU._0224_ ),
    .A2(\u_cpu.ALU._0813_ ),
    .B1(\u_cpu.ALU._0226_ ),
    .C1(\u_cpu.ALU._0227_ ),
    .D1(\u_cpu.ALU._0232_ ),
    .X(\u_cpu.ALU._0233_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2459_  (.A1(\u_cpu.ALU._1275_ ),
    .A2(\u_cpu.ALU._1092_ ),
    .B1(\u_cpu.ALU._0233_ ),
    .X(\u_cpu.ALU._0234_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._2460_  (.A1(\u_cpu.ALU._0221_ ),
    .A2(\u_cpu.ALU._0144_ ),
    .A3(\u_cpu.ALU._0223_ ),
    .B1(\u_cpu.ALU._0234_ ),
    .X(\u_cpu.ALU.ALUResult[21] ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2461_  (.A(\u_cpu.ALU._0216_ ),
    .B(\u_cpu.ALU._0215_ ),
    .Y(\u_cpu.ALU._0235_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU._2462_  (.A1_N(\u_cpu.ALU._0216_ ),
    .A2_N(\u_cpu.ALU._0215_ ),
    .B1(\u_cpu.ALU._0193_ ),
    .B2(\u_cpu.ALU._0191_ ),
    .X(\u_cpu.ALU._0236_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._2463_  (.A1(\u_cpu.ALU._0195_ ),
    .A2(\u_cpu.ALU._0198_ ),
    .B1(\u_cpu.ALU._0219_ ),
    .C1(\u_cpu.ALU._0222_ ),
    .X(\u_cpu.ALU._0237_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU._2464_  (.A1(\u_cpu.ALU._0235_ ),
    .A2(\u_cpu.ALU._0236_ ),
    .B1(\u_cpu.ALU._0237_ ),
    .B2(\u_cpu.ALU._0188_ ),
    .Y(\u_cpu.ALU._0238_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2465_  (.A(\u_cpu.ALU.SrcB[19] ),
    .B(\u_cpu.ALU.SrcB[18] ),
    .Y(\u_cpu.ALU._0239_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU._2466_  (.A(\u_cpu.ALU._0129_ ),
    .B(\u_cpu.ALU._0239_ ),
    .C(\u_cpu.ALU._0568_ ),
    .D(\u_cpu.ALU._0190_ ),
    .Y(\u_cpu.ALU._0240_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._2467_  (.A1(\u_cpu.ALU._0072_ ),
    .A2(\u_cpu.ALU._0240_ ),
    .B1(\u_cpu.ALU.SrcB[22] ),
    .C1(\u_cpu.ALU._0160_ ),
    .Y(\u_cpu.ALU._0241_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2468_  (.A1(\u_cpu.ALU._0072_ ),
    .A2(\u_cpu.ALU._0240_ ),
    .B1(\u_cpu.ALU._1346_ ),
    .X(\u_cpu.ALU._0242_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2469_  (.A1(\u_cpu.ALU.SrcB[22] ),
    .A2(\u_cpu.ALU._0242_ ),
    .B1(\u_cpu.ALU._0562_ ),
    .X(\u_cpu.ALU._0243_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2470_  (.A(\u_cpu.ALU._0067_ ),
    .B(\u_cpu.ALU._0240_ ),
    .Y(\u_cpu.ALU._0244_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2471_  (.A1(\u_cpu.ALU._1200_ ),
    .A2(\u_cpu.ALU._0244_ ),
    .B1(\u_cpu.ALU._0563_ ),
    .Y(\u_cpu.ALU._0245_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2472_  (.A1(\u_cpu.ALU._0245_ ),
    .A2(\u_cpu.ALU._0241_ ),
    .B1(\u_cpu.ALU._0562_ ),
    .Y(\u_cpu.ALU._0246_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2473_  (.A1(\u_cpu.ALU._0241_ ),
    .A2(\u_cpu.ALU._0243_ ),
    .B1(\u_cpu.ALU._0246_ ),
    .Y(\u_cpu.ALU._0247_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2474_  (.A(\u_cpu.ALU._0238_ ),
    .B(\u_cpu.ALU._0247_ ),
    .Y(\u_cpu.ALU._0248_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._2475_  (.A(\u_cpu.ALU._0247_ ),
    .Y(\u_cpu.ALU._0249_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU._2476_  (.A1(\u_cpu.ALU._0235_ ),
    .A2(\u_cpu.ALU._0236_ ),
    .B1(\u_cpu.ALU._0237_ ),
    .B2(\u_cpu.ALU._0188_ ),
    .C1(\u_cpu.ALU._0249_ ),
    .Y(\u_cpu.ALU._0250_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._2477_  (.A1(\u_cpu.ALU._0957_ ),
    .A2(\u_cpu.ALU._0560_ ),
    .B1(\u_cpu.ALU.SrcB[22] ),
    .C1(\u_cpu.ALU._0896_ ),
    .X(\u_cpu.ALU._0251_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2478_  (.A1(\u_cpu.ALU._0562_ ),
    .A2(\u_cpu.ALU._0563_ ),
    .B1(\u_cpu.ALU._0738_ ),
    .C1(\u_cpu.ALU._1149_ ),
    .D1(\u_cpu.ALU._0890_ ),
    .X(\u_cpu.ALU._0252_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.ALU._2479_  (.A1(\u_cpu.ALU._0749_ ),
    .A2(\u_cpu.ALU._0251_ ),
    .A3(\u_cpu.ALU._0252_ ),
    .B1(\u_cpu.ALU.SrcB[22] ),
    .B2(\u_cpu.ALU._0560_ ),
    .X(\u_cpu.ALU._0253_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2480_  (.A0(\u_cpu.ALU._0560_ ),
    .A1(\u_cpu.ALU._0216_ ),
    .A2(\u_cpu.ALU._0837_ ),
    .A3(\u_cpu.ALU._0547_ ),
    .S0(\u_cpu.ALU._0723_ ),
    .S1(\u_cpu.ALU._0899_ ),
    .X(\u_cpu.ALU._0254_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.ALU._2481_  (.A0(\u_cpu.ALU._0151_ ),
    .A1(\u_cpu.ALU._0254_ ),
    .S(\u_cpu.ALU._0786_ ),
    .X(\u_cpu.ALU._0255_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU._2482_  (.A(\u_cpu.ALU._0758_ ),
    .B(\u_cpu.ALU._0761_ ),
    .X(\u_cpu.ALU._0256_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._2483_  (.A1(\u_cpu.ALU._1219_ ),
    .A2(\u_cpu.ALU._1115_ ),
    .A3(\u_cpu.ALU._0026_ ),
    .B1(\u_cpu.ALU._0819_ ),
    .X(\u_cpu.ALU._0257_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU._2484_  (.A1(\u_cpu.ALU._1212_ ),
    .A2(\u_cpu.ALU._0024_ ),
    .B1(\u_cpu.ALU._0255_ ),
    .B2(\u_cpu.ALU._0256_ ),
    .C1(\u_cpu.ALU._0257_ ),
    .Y(\u_cpu.ALU._0258_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2485_  (.A1(\u_cpu.ALU._1144_ ),
    .A2(\u_cpu.ALU._1127_ ),
    .B1(\u_cpu.ALU._0258_ ),
    .Y(\u_cpu.ALU._0259_ ));
 sky130_fd_sc_hd__a2111o_2 \u_cpu.ALU._2486_  (.A1(\u_cpu.ALU.Product_Wallace[22] ),
    .A2(\u_cpu.ALU._1338_ ),
    .B1(\u_cpu.ALU._0115_ ),
    .C1(\u_cpu.ALU._0253_ ),
    .D1(\u_cpu.ALU._0259_ ),
    .X(\u_cpu.ALU._0260_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._2487_  (.A1(\u_cpu.ALU._0248_ ),
    .A2(\u_cpu.ALU._0144_ ),
    .A3(\u_cpu.ALU._0250_ ),
    .B1(\u_cpu.ALU._0260_ ),
    .X(\u_cpu.ALU.ALUResult[22] ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2488_  (.A1(\u_cpu.ALU._0245_ ),
    .A2(\u_cpu.ALU._0241_ ),
    .B1(\u_cpu.ALU._0562_ ),
    .X(\u_cpu.ALU._0261_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU._2489_  (.A(\u_cpu.ALU._0129_ ),
    .B(\u_cpu.ALU._0239_ ),
    .C(\u_cpu.ALU._0568_ ),
    .D(\u_cpu.ALU._0190_ ),
    .X(\u_cpu.ALU._0262_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU._2490_  (.A(\u_cpu.ALU._0128_ ),
    .B(\u_cpu.ALU._0066_ ),
    .C(\u_cpu.ALU._0262_ ),
    .D(\u_cpu.ALU._0563_ ),
    .Y(\u_cpu.ALU._0263_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU._2491_  (.A1(\u_cpu.ALU._0752_ ),
    .A2(\u_cpu.ALU._0873_ ),
    .A3(\u_cpu.ALU._1018_ ),
    .B1(\u_cpu.ALU.SrcB[23] ),
    .C1(\u_cpu.ALU._0263_ ),
    .X(\u_cpu.ALU._0264_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU._2492_  (.A(\u_cpu.ALU._0240_ ),
    .B(\u_cpu.ALU.SrcB[22] ),
    .C(\u_cpu.ALU._0072_ ),
    .Y(\u_cpu.ALU._0265_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2493_  (.A1(\u_cpu.ALU._1200_ ),
    .A2(\u_cpu.ALU._0265_ ),
    .B1(\u_cpu.ALU._0553_ ),
    .Y(\u_cpu.ALU._0266_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2494_  (.A(\u_cpu.ALU._0552_ ),
    .B(\u_cpu.ALU._0266_ ),
    .Y(\u_cpu.ALU._0267_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._2495_  (.A1(\u_cpu.ALU._0873_ ),
    .A2(\u_cpu.ALU._0920_ ),
    .B1(\u_cpu.ALU.SrcB[23] ),
    .C1(\u_cpu.ALU._0263_ ),
    .Y(\u_cpu.ALU._0268_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2496_  (.A1(\u_cpu.ALU._0266_ ),
    .A2(\u_cpu.ALU._0268_ ),
    .B1(\u_cpu.ALU._0552_ ),
    .X(\u_cpu.ALU._0269_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2497_  (.A1(\u_cpu.ALU._0264_ ),
    .A2(\u_cpu.ALU._0267_ ),
    .B1(\u_cpu.ALU._0269_ ),
    .Y(\u_cpu.ALU._0270_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2498_  (.A1(\u_cpu.ALU._0261_ ),
    .A2(\u_cpu.ALU._0248_ ),
    .B1(\u_cpu.ALU._0270_ ),
    .X(\u_cpu.ALU._0271_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2499_  (.A1(\u_cpu.ALU._0873_ ),
    .A2(\u_cpu.ALU._0920_ ),
    .B1(\u_cpu.ALU._0263_ ),
    .Y(\u_cpu.ALU._0272_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2500_  (.A1(\u_cpu.ALU._0553_ ),
    .A2(\u_cpu.ALU._0272_ ),
    .B1(\u_cpu.ALU._0555_ ),
    .Y(\u_cpu.ALU._0273_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2501_  (.A1(\u_cpu.ALU._0266_ ),
    .A2(\u_cpu.ALU._0268_ ),
    .B1(\u_cpu.ALU._0552_ ),
    .Y(\u_cpu.ALU._0274_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2502_  (.A1(\u_cpu.ALU._0273_ ),
    .A2(\u_cpu.ALU._0268_ ),
    .B1(\u_cpu.ALU._0274_ ),
    .Y(\u_cpu.ALU._0275_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._2503_  (.A1(\u_cpu.ALU._0238_ ),
    .A2(\u_cpu.ALU._0247_ ),
    .B1(\u_cpu.ALU._0246_ ),
    .C1(\u_cpu.ALU._0275_ ),
    .X(\u_cpu.ALU._0276_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2504_  (.A0(\u_cpu.ALU._0555_ ),
    .A1(\u_cpu.ALU._0560_ ),
    .A2(\u_cpu.ALU.SrcA[21] ),
    .A3(\u_cpu.ALU._0837_ ),
    .S0(\u_cpu.ALU._0794_ ),
    .S1(\u_cpu.ALU._0826_ ),
    .X(\u_cpu.ALU._0277_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU._2505_  (.A(\u_cpu.ALU._0277_ ),
    .B(\u_cpu.ALU._0769_ ),
    .X(\u_cpu.ALU._0278_ ));
 sky130_fd_sc_hd__a2111oi_2 \u_cpu.ALU._2506_  (.A1(\u_cpu.ALU._1145_ ),
    .A2(\u_cpu.ALU._0176_ ),
    .B1(\u_cpu.ALU._0278_ ),
    .C1(\u_cpu.ALU._0761_ ),
    .D1(\u_cpu.ALU._0758_ ),
    .Y(\u_cpu.ALU._0279_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2507_  (.A(\u_cpu.ALU._1257_ ),
    .B(\u_cpu.ALU._0279_ ),
    .Y(\u_cpu.ALU._0280_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2508_  (.A1(\u_cpu.ALU._1212_ ),
    .A2(\u_cpu.ALU._0052_ ),
    .B1(\u_cpu.ALU._0280_ ),
    .X(\u_cpu.ALU._0281_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2509_  (.A1(\u_cpu.ALU._1151_ ),
    .A2(\u_cpu.ALU._0281_ ),
    .B1(\u_cpu.ALU._1275_ ),
    .X(\u_cpu.ALU._0282_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._2510_  (.A(\u_cpu.ALU._0555_ ),
    .B(\u_cpu.ALU.SrcB[23] ),
    .C(\u_cpu.ALU._0058_ ),
    .X(\u_cpu.ALU._0283_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2511_  (.A1(\u_cpu.ALU.SrcB[23] ),
    .A2(\u_cpu.ALU._0060_ ),
    .B1(\u_cpu.ALU._1338_ ),
    .B2(\u_cpu.ALU.Product_Wallace[23] ),
    .C1(\u_cpu.ALU._0283_ ),
    .X(\u_cpu.ALU._0284_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2512_  (.A1(\u_cpu.ALU._0555_ ),
    .A2(\u_cpu.ALU.SrcB[23] ),
    .B1(\u_cpu.ALU._0061_ ),
    .C1(\u_cpu.ALU._1226_ ),
    .D1(\u_cpu.ALU._1332_ ),
    .X(\u_cpu.ALU._0285_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.ALU._2513_  (.A(\u_cpu.ALU._0554_ ),
    .B(\u_cpu.ALU._0556_ ),
    .C(\u_cpu.ALU._1020_ ),
    .X(\u_cpu.ALU._0286_ ));
 sky130_fd_sc_hd__or3b_2 \u_cpu.ALU._2514_  (.A(\u_cpu.ALU._0115_ ),
    .B(\u_cpu.ALU._0285_ ),
    .C_N(\u_cpu.ALU._0286_ ),
    .X(\u_cpu.ALU._0287_ ));
 sky130_fd_sc_hd__or4b_2 \u_cpu.ALU._2515_  (.A(\u_cpu.ALU._0761_ ),
    .B(\u_cpu.ALU._0279_ ),
    .C(\u_cpu.ALU._1257_ ),
    .D_N(\u_cpu.ALU._1156_ ),
    .X(\u_cpu.ALU._0288_ ));
 sky130_fd_sc_hd__or4b_2 \u_cpu.ALU._2516_  (.A(\u_cpu.ALU._0282_ ),
    .B(\u_cpu.ALU._0284_ ),
    .C(\u_cpu.ALU._0287_ ),
    .D_N(\u_cpu.ALU._0288_ ),
    .X(\u_cpu.ALU._0289_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU._2517_  (.A1(\u_cpu.ALU._0271_ ),
    .A2(\u_cpu.ALU._0144_ ),
    .A3(\u_cpu.ALU._0276_ ),
    .B1(\u_cpu.ALU._0289_ ),
    .Y(\u_cpu.ALU._0290_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._2518_  (.A(\u_cpu.ALU._0290_ ),
    .Y(\u_cpu.ALU.ALUResult[23] ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2519_  (.A(\u_cpu.ALU.SrcB[23] ),
    .B(\u_cpu.ALU.SrcB[22] ),
    .Y(\u_cpu.ALU._0291_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU._2520_  (.A(\u_cpu.ALU._0128_ ),
    .B(\u_cpu.ALU._0066_ ),
    .C(\u_cpu.ALU._0262_ ),
    .D(\u_cpu.ALU._0291_ ),
    .Y(\u_cpu.ALU._0292_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU._2521_  (.A1(\u_cpu.ALU._0160_ ),
    .A2(\u_cpu.ALU._0292_ ),
    .B1_N(\u_cpu.ALU._0444_ ),
    .Y(\u_cpu.ALU._0293_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._2522_  (.A(\u_cpu.ALU._0433_ ),
    .Y(\u_cpu.ALU._0294_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.ALU._2523_  (.A1(\u_cpu.ALU._0746_ ),
    .A2(\u_cpu.ALU._0814_ ),
    .B1(\u_cpu.ALU._0244_ ),
    .B2(\u_cpu.ALU._0291_ ),
    .C1(\u_cpu.ALU._0444_ ),
    .Y(\u_cpu.ALU._0295_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.ALU._2524_  (.A(\u_cpu.ALU._0293_ ),
    .B(\u_cpu.ALU._0294_ ),
    .C(\u_cpu.ALU._0295_ ),
    .X(\u_cpu.ALU._0296_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2525_  (.A(\u_cpu.ALU._0296_ ),
    .X(\u_cpu.ALU._0297_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2526_  (.A1(\u_cpu.ALU._0295_ ),
    .A2(\u_cpu.ALU._0293_ ),
    .B1(\u_cpu.ALU._0294_ ),
    .Y(\u_cpu.ALU._0298_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.ALU._2527_  (.A1(\u_cpu.ALU._0195_ ),
    .A2(\u_cpu.ALU._0198_ ),
    .B1(\u_cpu.ALU._0215_ ),
    .B2(\u_cpu.ALU._0216_ ),
    .C1(\u_cpu.ALU._0219_ ),
    .Y(\u_cpu.ALU._0299_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU._2528_  (.A(\u_cpu.ALU._0299_ ),
    .B(\u_cpu.ALU._0218_ ),
    .C(\u_cpu.ALU._0247_ ),
    .D(\u_cpu.ALU._0275_ ),
    .Y(\u_cpu.ALU._0300_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2529_  (.A(\u_cpu.ALU._0183_ ),
    .B(\u_cpu.ALU._0300_ ),
    .Y(\u_cpu.ALU._0301_ ));
 sky130_fd_sc_hd__a41oi_2 \u_cpu.ALU._2530_  (.A1(\u_cpu.ALU._0167_ ),
    .A2(\u_cpu.ALU._0105_ ),
    .A3(\u_cpu.ALU._0142_ ),
    .A4(\u_cpu.ALU._0124_ ),
    .B1(\u_cpu.ALU._0186_ ),
    .Y(\u_cpu.ALU._0302_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU._2531_  (.A1(\u_cpu.ALU._0837_ ),
    .A2(\u_cpu.ALU._0194_ ),
    .A3(\u_cpu.ALU._0195_ ),
    .B1(\u_cpu.ALU._0215_ ),
    .B2(\u_cpu.ALU._0216_ ),
    .X(\u_cpu.ALU._0303_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU._2532_  (.A1(\u_cpu.ALU._0267_ ),
    .A2(\u_cpu.ALU._0264_ ),
    .B1(\u_cpu.ALU._0246_ ),
    .B2(\u_cpu.ALU._0274_ ),
    .X(\u_cpu.ALU._0304_ ));
 sky130_fd_sc_hd__a41oi_2 \u_cpu.ALU._2533_  (.A1(\u_cpu.ALU._0247_ ),
    .A2(\u_cpu.ALU._0275_ ),
    .A3(\u_cpu.ALU._0303_ ),
    .A4(\u_cpu.ALU._0218_ ),
    .B1(\u_cpu.ALU._0304_ ),
    .Y(\u_cpu.ALU._0305_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2534_  (.A1(\u_cpu.ALU._0302_ ),
    .A2(\u_cpu.ALU._0300_ ),
    .B1(\u_cpu.ALU._0305_ ),
    .Y(\u_cpu.ALU._0306_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2535_  (.A1(\u_cpu.ALU._0297_ ),
    .A2(\u_cpu.ALU._0298_ ),
    .B1(\u_cpu.ALU._0087_ ),
    .B2(\u_cpu.ALU._0301_ ),
    .C1(\u_cpu.ALU._0306_ ),
    .X(\u_cpu.ALU._0307_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2536_  (.A(\u_cpu.ALU._0015_ ),
    .B(\u_cpu.ALU._0084_ ),
    .Y(\u_cpu.ALU._0308_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._2537_  (.A(\u_cpu.ALU._1183_ ),
    .B(\u_cpu.ALU._1307_ ),
    .C(\u_cpu.ALU._0308_ ),
    .Y(\u_cpu.ALU._0309_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2538_  (.A1(\u_cpu.ALU._0193_ ),
    .A2(\u_cpu.ALU._0191_ ),
    .B1(\u_cpu.ALU._0196_ ),
    .C1(\u_cpu.ALU._0217_ ),
    .D1(\u_cpu.ALU._0218_ ),
    .X(\u_cpu.ALU._0310_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._2539_  (.A(\u_cpu.ALU._0562_ ),
    .B(\u_cpu.ALU._0245_ ),
    .C(\u_cpu.ALU._0241_ ),
    .Y(\u_cpu.ALU._0311_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2540_  (.A1(\u_cpu.ALU._0267_ ),
    .A2(\u_cpu.ALU._0264_ ),
    .B1(\u_cpu.ALU._0311_ ),
    .C1(\u_cpu.ALU._0261_ ),
    .D1(\u_cpu.ALU._0269_ ),
    .X(\u_cpu.ALU._0312_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU._2541_  (.A(\u_cpu.ALU._0126_ ),
    .B(\u_cpu.ALU._0185_ ),
    .C(\u_cpu.ALU._0310_ ),
    .D(\u_cpu.ALU._0312_ ),
    .Y(\u_cpu.ALU._0313_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2542_  (.A1(\u_cpu.ALU._0309_ ),
    .A2(\u_cpu.ALU._0086_ ),
    .B1(\u_cpu.ALU._0313_ ),
    .Y(\u_cpu.ALU._0314_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._2543_  (.A1(\u_cpu.ALU._0306_ ),
    .A2(\u_cpu.ALU._0314_ ),
    .B1(\u_cpu.ALU._0298_ ),
    .C1(\u_cpu.ALU._0297_ ),
    .Y(\u_cpu.ALU._0315_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2544_  (.A1(\u_cpu.ALU._1063_ ),
    .A2(\u_cpu.ALU._0056_ ),
    .B1(\u_cpu.ALU._1158_ ),
    .X(\u_cpu.ALU._0316_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU._2545_  (.A1(\u_cpu.ALU._1283_ ),
    .A2(\u_cpu.ALU._0761_ ),
    .A3(\u_cpu.ALU._0766_ ),
    .B1(\u_cpu.ALU._0316_ ),
    .X(\u_cpu.ALU._0317_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU._2546_  (.A1(\u_cpu.ALU._1332_ ),
    .A2(\u_cpu.ALU._1331_ ),
    .A3(\u_cpu.ALU._0061_ ),
    .B1(\u_cpu.ALU._0813_ ),
    .B2(\u_cpu.ALU._0465_ ),
    .X(\u_cpu.ALU._0318_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU._2547_  (.A1(\u_cpu.ALU._0444_ ),
    .A2(\u_cpu.ALU._0754_ ),
    .B1(\u_cpu.ALU._0822_ ),
    .B2(\u_cpu.ALU.Product_Wallace[24] ),
    .X(\u_cpu.ALU._0319_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._2548_  (.A1(\u_cpu.ALU._0433_ ),
    .A2(\u_cpu.ALU._0444_ ),
    .A3(\u_cpu.ALU._0058_ ),
    .B1(\u_cpu.ALU._0319_ ),
    .X(\u_cpu.ALU._0320_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2549_  (.A0(\u_cpu.ALU._0433_ ),
    .A1(\u_cpu.ALU._0555_ ),
    .A2(\u_cpu.ALU._0560_ ),
    .A3(\u_cpu.ALU._0216_ ),
    .S0(\u_cpu.ALU._0722_ ),
    .S1(\u_cpu.ALU._0899_ ),
    .X(\u_cpu.ALU._0321_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2550_  (.A0(\u_cpu.ALU._1321_ ),
    .A1(\u_cpu.ALU._0090_ ),
    .A2(\u_cpu.ALU._0202_ ),
    .A3(\u_cpu.ALU._0321_ ),
    .S0(\u_cpu.ALU._0786_ ),
    .S1(\u_cpu.ALU._1219_ ),
    .X(\u_cpu.ALU._0322_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU._2551_  (.A(\u_cpu.ALU._1196_ ),
    .B(\u_cpu.ALU._0738_ ),
    .C(\u_cpu.ALU._1226_ ),
    .D(\u_cpu.ALU._0963_ ),
    .X(\u_cpu.ALU._0323_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU._2552_  (.A1(\u_cpu.ALU._0322_ ),
    .A2(\u_cpu.ALU._1144_ ),
    .B1(\u_cpu.ALU._0819_ ),
    .B2(\u_cpu.ALU._0323_ ),
    .X(\u_cpu.ALU._0324_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._2553_  (.A1(\u_cpu.ALU._0454_ ),
    .A2(\u_cpu.ALU._0318_ ),
    .B1(\u_cpu.ALU._0320_ ),
    .C1(\u_cpu.ALU._0324_ ),
    .X(\u_cpu.ALU._0325_ ));
 sky130_fd_sc_hd__a311o_2 \u_cpu.ALU._2554_  (.A1(\u_cpu.ALU._0307_ ),
    .A2(\u_cpu.ALU._0975_ ),
    .A3(\u_cpu.ALU._0315_ ),
    .B1(\u_cpu.ALU._0317_ ),
    .C1(\u_cpu.ALU._0325_ ),
    .X(\u_cpu.ALU.ALUResult[24] ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU._2555_  (.A1(\u_cpu.ALU._0750_ ),
    .A2(\u_cpu.ALU._0751_ ),
    .A3(\u_cpu.ALU._0708_ ),
    .B1(\u_cpu.ALU._0444_ ),
    .X(\u_cpu.ALU._0326_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._2556_  (.A1(\u_cpu.ALU._0160_ ),
    .A2(\u_cpu.ALU._0292_ ),
    .B1(\u_cpu.ALU._0326_ ),
    .C1(\u_cpu.ALU.SrcB[25] ),
    .X(\u_cpu.ALU._0327_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU._2557_  (.A1(\u_cpu.ALU._0873_ ),
    .A2(\u_cpu.ALU._0920_ ),
    .B1(\u_cpu.ALU._0444_ ),
    .B2(\u_cpu.ALU._0292_ ),
    .C1(\u_cpu.ALU.SrcB[25] ),
    .Y(\u_cpu.ALU._0328_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU._2558_  (.A1(\u_cpu.ALU._0327_ ),
    .A2(\u_cpu.ALU._0328_ ),
    .B1_N(\u_cpu.ALU._0475_ ),
    .Y(\u_cpu.ALU._0329_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU._2559_  (.A_N(\u_cpu.ALU._0475_ ),
    .B(\u_cpu.ALU._0327_ ),
    .C(\u_cpu.ALU._0328_ ),
    .Y(\u_cpu.ALU._0330_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.ALU._2560_  (.A(\u_cpu.ALU._0329_ ),
    .B_N(\u_cpu.ALU._0330_ ),
    .X(\u_cpu.ALU._0331_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2561_  (.A1(\u_cpu.ALU._0297_ ),
    .A2(\u_cpu.ALU._0315_ ),
    .B1(\u_cpu.ALU._0331_ ),
    .Y(\u_cpu.ALU._0332_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._2562_  (.A1(\u_cpu.ALU._0297_ ),
    .A2(\u_cpu.ALU._0315_ ),
    .A3(\u_cpu.ALU._0331_ ),
    .B1(\u_cpu.ALU._0921_ ),
    .X(\u_cpu.ALU._0333_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2563_  (.A1(\u_cpu.ALU._0475_ ),
    .A2(\u_cpu.ALU.SrcB[25] ),
    .B1(\u_cpu.ALU._0061_ ),
    .C1(\u_cpu.ALU._1331_ ),
    .D1(\u_cpu.ALU._1332_ ),
    .X(\u_cpu.ALU._0334_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.ALU._2564_  (.A1(\u_cpu.ALU.SrcB[25] ),
    .A2(\u_cpu.ALU._0060_ ),
    .B1(\u_cpu.ALU._0813_ ),
    .B2(\u_cpu.ALU._0507_ ),
    .C1(\u_cpu.ALU._0334_ ),
    .Y(\u_cpu.ALU._0335_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.ALU._2565_  (.A1(\u_cpu.ALU._0496_ ),
    .A2(\u_cpu.ALU._0058_ ),
    .B1(\u_cpu.ALU._1338_ ),
    .B2(\u_cpu.ALU.Product_Wallace[25] ),
    .C1(\u_cpu.ALU._0115_ ),
    .Y(\u_cpu.ALU._0336_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2566_  (.A0(\u_cpu.ALU._0475_ ),
    .A1(\u_cpu.ALU._0433_ ),
    .A2(\u_cpu.ALU._0555_ ),
    .A3(\u_cpu.ALU._0560_ ),
    .S0(\u_cpu.ALU._0723_ ),
    .S1(\u_cpu.ALU._0899_ ),
    .X(\u_cpu.ALU._0337_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2567_  (.A0(\u_cpu.ALU._1329_ ),
    .A1(\u_cpu.ALU._0110_ ),
    .A2(\u_cpu.ALU._0230_ ),
    .A3(\u_cpu.ALU._0337_ ),
    .S0(\u_cpu.ALU._1279_ ),
    .S1(\u_cpu.ALU._1212_ ),
    .X(\u_cpu.ALU._0339_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU._2568_  (.A1(\u_cpu.ALU._0819_ ),
    .A2(\u_cpu.ALU._1227_ ),
    .B1(\u_cpu.ALU._0339_ ),
    .B2(\u_cpu.ALU._1283_ ),
    .Y(\u_cpu.ALU._0340_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2569_  (.A1(\u_cpu.ALU._1283_ ),
    .A2(\u_cpu.ALU._1214_ ),
    .B1(\u_cpu.ALU._0335_ ),
    .C1(\u_cpu.ALU._0336_ ),
    .D1(\u_cpu.ALU._0340_ ),
    .X(\u_cpu.ALU._0341_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2570_  (.A1(\u_cpu.ALU._0332_ ),
    .A2(\u_cpu.ALU._0333_ ),
    .B1(\u_cpu.ALU._0341_ ),
    .Y(\u_cpu.ALU.ALUResult[25] ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2571_  (.A1(\u_cpu.ALU.SrcA[26] ),
    .A2(\u_cpu.ALU.SrcB[26] ),
    .B1(\u_cpu.ALU._0061_ ),
    .C1(\u_cpu.ALU._1226_ ),
    .D1(\u_cpu.ALU._1332_ ),
    .X(\u_cpu.ALU._0342_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2572_  (.A1(\u_cpu.ALU.SrcB[26] ),
    .A2(\u_cpu.ALU._0060_ ),
    .B1(\u_cpu.ALU._0813_ ),
    .B2(\u_cpu.ALU._0423_ ),
    .C1(\u_cpu.ALU._0342_ ),
    .X(\u_cpu.ALU._0343_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2573_  (.A1(\u_cpu.ALU._0412_ ),
    .A2(\u_cpu.ALU._0058_ ),
    .B1(\u_cpu.ALU._1338_ ),
    .B2(\u_cpu.ALU.Product_Wallace[26] ),
    .C1(\u_cpu.ALU._0115_ ),
    .X(\u_cpu.ALU._0344_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU._2574_  (.A1(\u_cpu.ALU._1275_ ),
    .A2(\u_cpu.ALU._1249_ ),
    .B1(\u_cpu.ALU._0343_ ),
    .C1(\u_cpu.ALU._0344_ ),
    .X(\u_cpu.ALU._0345_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2575_  (.A0(\u_cpu.ALU.SrcA[26] ),
    .A1(\u_cpu.ALU._0475_ ),
    .A2(\u_cpu.ALU._0433_ ),
    .A3(\u_cpu.ALU._0555_ ),
    .S0(\u_cpu.ALU._0723_ ),
    .S1(\u_cpu.ALU._0899_ ),
    .X(\u_cpu.ALU._0346_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2576_  (.A0(\u_cpu.ALU._0023_ ),
    .A1(\u_cpu.ALU._0151_ ),
    .A2(\u_cpu.ALU._0254_ ),
    .A3(\u_cpu.ALU._0346_ ),
    .S0(\u_cpu.ALU._1279_ ),
    .S1(\u_cpu.ALU._1212_ ),
    .X(\u_cpu.ALU._0347_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU._2577_  (.A1_N(\u_cpu.ALU._0228_ ),
    .A2_N(\u_cpu.ALU._1262_ ),
    .B1(\u_cpu.ALU._0347_ ),
    .B2(\u_cpu.ALU._1283_ ),
    .X(\u_cpu.ALU._0349_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._2578_  (.A(\u_cpu.ALU._0330_ ),
    .Y(\u_cpu.ALU._0350_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU._2579_  (.A(\u_cpu.ALU._0293_ ),
    .B(\u_cpu.ALU._0294_ ),
    .C(\u_cpu.ALU._0295_ ),
    .Y(\u_cpu.ALU._0351_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2580_  (.A(\u_cpu.ALU._0351_ ),
    .B(\u_cpu.ALU._0329_ ),
    .Y(\u_cpu.ALU._0352_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU._2581_  (.A_N(\u_cpu.ALU._0331_ ),
    .B(\u_cpu.ALU._0298_ ),
    .C(\u_cpu.ALU._0297_ ),
    .Y(\u_cpu.ALU._0353_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2582_  (.A1(\u_cpu.ALU._0087_ ),
    .A2(\u_cpu.ALU._0301_ ),
    .B1(\u_cpu.ALU._0306_ ),
    .Y(\u_cpu.ALU._0354_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU._2583_  (.A1(\u_cpu.ALU._0350_ ),
    .A2(\u_cpu.ALU._0352_ ),
    .B1(\u_cpu.ALU._0353_ ),
    .B2(\u_cpu.ALU._0354_ ),
    .Y(\u_cpu.ALU._0355_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2584_  (.A(\u_cpu.ALU.SrcB[25] ),
    .B(\u_cpu.ALU._0444_ ),
    .Y(\u_cpu.ALU._0356_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU._2585_  (.A_N(\u_cpu.ALU._0067_ ),
    .B(\u_cpu.ALU._0262_ ),
    .C(\u_cpu.ALU._0291_ ),
    .D(\u_cpu.ALU._0356_ ),
    .Y(\u_cpu.ALU._0357_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU._2586_  (.A1(\u_cpu.ALU._0963_ ),
    .A2(\u_cpu.ALU._0900_ ),
    .A3(\u_cpu.ALU._1018_ ),
    .B1(\u_cpu.ALU.SrcB[26] ),
    .C1(\u_cpu.ALU._0357_ ),
    .X(\u_cpu.ALU._0358_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2587_  (.A1(\u_cpu.ALU._0160_ ),
    .A2(\u_cpu.ALU._0357_ ),
    .B1(\u_cpu.ALU.SrcB[26] ),
    .X(\u_cpu.ALU._0360_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2588_  (.A(\u_cpu.ALU._0588_ ),
    .B(\u_cpu.ALU._0360_ ),
    .Y(\u_cpu.ALU._0361_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._2589_  (.A1(\u_cpu.ALU._0873_ ),
    .A2(\u_cpu.ALU._0920_ ),
    .B1(\u_cpu.ALU.SrcB[26] ),
    .C1(\u_cpu.ALU._0357_ ),
    .Y(\u_cpu.ALU._0362_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2590_  (.A1(\u_cpu.ALU._0360_ ),
    .A2(\u_cpu.ALU._0362_ ),
    .B1(\u_cpu.ALU._0588_ ),
    .X(\u_cpu.ALU._0363_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2591_  (.A1(\u_cpu.ALU._0358_ ),
    .A2(\u_cpu.ALU._0361_ ),
    .B1(\u_cpu.ALU._0363_ ),
    .X(\u_cpu.ALU._0364_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2592_  (.A(\u_cpu.ALU._0355_ ),
    .B(\u_cpu.ALU._0364_ ),
    .Y(\u_cpu.ALU._0365_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2593_  (.A1(\u_cpu.ALU._0360_ ),
    .A2(\u_cpu.ALU._0362_ ),
    .B1(\u_cpu.ALU._0588_ ),
    .Y(\u_cpu.ALU._0366_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._2594_  (.A(\u_cpu.ALU._0588_ ),
    .B(\u_cpu.ALU._0360_ ),
    .C(\u_cpu.ALU._0362_ ),
    .X(\u_cpu.ALU._0367_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2595_  (.A1(\u_cpu.ALU._0351_ ),
    .A2(\u_cpu.ALU._0329_ ),
    .B1(\u_cpu.ALU._0330_ ),
    .Y(\u_cpu.ALU._0368_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU._2596_  (.A1(\u_cpu.ALU._0366_ ),
    .A2(\u_cpu.ALU._0367_ ),
    .B1(\u_cpu.ALU._0353_ ),
    .B2(\u_cpu.ALU._0354_ ),
    .C1(\u_cpu.ALU._0368_ ),
    .Y(\u_cpu.ALU._0369_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU._2597_  (.A(\u_cpu.ALU._0890_ ),
    .B(\u_cpu.ALU._0365_ ),
    .C(\u_cpu.ALU._0369_ ),
    .D(\u_cpu.ALU._0061_ ),
    .Y(\u_cpu.ALU._0371_ ));
 sky130_fd_sc_hd__or3b_2 \u_cpu.ALU._2598_  (.A(\u_cpu.ALU._0345_ ),
    .B(\u_cpu.ALU._0349_ ),
    .C_N(\u_cpu.ALU._0371_ ),
    .X(\u_cpu.ALU._0372_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU._2599_  (.A(\u_cpu.ALU._0372_ ),
    .X(\u_cpu.ALU.ALUResult[26] ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2600_  (.A1(\u_cpu.ALU._0358_ ),
    .A2(\u_cpu.ALU._0361_ ),
    .B1(\u_cpu.ALU._0355_ ),
    .Y(\u_cpu.ALU._0373_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU._2601_  (.A(\u_cpu.ALU.SrcB[26] ),
    .B(\u_cpu.ALU.SrcB[25] ),
    .C(\u_cpu.ALU._0444_ ),
    .Y(\u_cpu.ALU._0374_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU._2602_  (.A_N(\u_cpu.ALU._0067_ ),
    .B(\u_cpu.ALU._0262_ ),
    .C(\u_cpu.ALU._0291_ ),
    .D(\u_cpu.ALU._0374_ ),
    .Y(\u_cpu.ALU._0375_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2603_  (.A1(\u_cpu.ALU._0160_ ),
    .A2(\u_cpu.ALU._0375_ ),
    .B1(\u_cpu.ALU.SrcB[27] ),
    .X(\u_cpu.ALU._0376_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU._2604_  (.A1(\u_cpu.ALU._0711_ ),
    .A2(\u_cpu.ALU._0920_ ),
    .B1(\u_cpu.ALU.SrcB[26] ),
    .B2(\u_cpu.ALU._0357_ ),
    .C1(\u_cpu.ALU.SrcB[27] ),
    .Y(\u_cpu.ALU._0377_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2605_  (.A1(\u_cpu.ALU._0376_ ),
    .A2(\u_cpu.ALU._0377_ ),
    .B1(\u_cpu.ALU._0338_ ),
    .Y(\u_cpu.ALU._0378_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._2606_  (.A(\u_cpu.ALU._0376_ ),
    .B(\u_cpu.ALU._0377_ ),
    .C(\u_cpu.ALU._0338_ ),
    .X(\u_cpu.ALU._0379_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU._2607_  (.A1_N(\u_cpu.ALU._0363_ ),
    .A2_N(\u_cpu.ALU._0373_ ),
    .B1(\u_cpu.ALU._0378_ ),
    .B2(\u_cpu.ALU._0379_ ),
    .Y(\u_cpu.ALU._0381_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._2608_  (.A(\u_cpu.ALU._0359_ ),
    .B(\u_cpu.ALU._0376_ ),
    .C(\u_cpu.ALU._0377_ ),
    .Y(\u_cpu.ALU._0382_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2609_  (.A1(\u_cpu.ALU._0376_ ),
    .A2(\u_cpu.ALU._0377_ ),
    .B1(\u_cpu.ALU._0359_ ),
    .X(\u_cpu.ALU._0383_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU._2610_  (.A1(\u_cpu.ALU._0382_ ),
    .A2(\u_cpu.ALU._0383_ ),
    .B1(\u_cpu.ALU._0355_ ),
    .B2(\u_cpu.ALU._0364_ ),
    .Y(\u_cpu.ALU._0384_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2611_  (.A(\u_cpu.ALU._0384_ ),
    .B(\u_cpu.ALU._0363_ ),
    .Y(\u_cpu.ALU._0385_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2612_  (.A1(\u_cpu.ALU._0338_ ),
    .A2(\u_cpu.ALU.SrcB[27] ),
    .B1(\u_cpu.ALU._0061_ ),
    .C1(\u_cpu.ALU._1331_ ),
    .D1(\u_cpu.ALU._1332_ ),
    .X(\u_cpu.ALU._0386_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2613_  (.A1(\u_cpu.ALU._0380_ ),
    .A2(\u_cpu.ALU._0058_ ),
    .B1(\u_cpu.ALU._1338_ ),
    .B2(\u_cpu.ALU.Product_Wallace[27] ),
    .C1(\u_cpu.ALU._0386_ ),
    .X(\u_cpu.ALU._0387_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2614_  (.A1(\u_cpu.ALU.SrcB[27] ),
    .A2(\u_cpu.ALU._0060_ ),
    .B1(\u_cpu.ALU._0813_ ),
    .B2(\u_cpu.ALU._0391_ ),
    .C1(\u_cpu.ALU._0115_ ),
    .X(\u_cpu.ALU._0388_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.ALU._2615_  (.A_N(\u_cpu.ALU._1278_ ),
    .B(\u_cpu.ALU._0738_ ),
    .C(\u_cpu.ALU._1331_ ),
    .D(\u_cpu.ALU._1332_ ),
    .X(\u_cpu.ALU._0389_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2616_  (.A0(\u_cpu.ALU._0338_ ),
    .A1(\u_cpu.ALU.SrcA[26] ),
    .A2(\u_cpu.ALU._0475_ ),
    .A3(\u_cpu.ALU._0433_ ),
    .S0(\u_cpu.ALU._0722_ ),
    .S1(\u_cpu.ALU._0790_ ),
    .X(\u_cpu.ALU._0390_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2617_  (.A0(\u_cpu.ALU._0051_ ),
    .A1(\u_cpu.ALU._0176_ ),
    .A2(\u_cpu.ALU._0277_ ),
    .A3(\u_cpu.ALU._0390_ ),
    .S0(\u_cpu.ALU._0786_ ),
    .S1(\u_cpu.ALU._1076_ ),
    .X(\u_cpu.ALU._0392_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2618_  (.A1(\u_cpu.ALU._0759_ ),
    .A2(\u_cpu.ALU._0392_ ),
    .B1(\u_cpu.ALU._0738_ ),
    .C1(\u_cpu.ALU._1332_ ),
    .D1(\u_cpu.ALU._1331_ ),
    .X(\u_cpu.ALU._0393_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU._2619_  (.A1(\u_cpu.ALU._1275_ ),
    .A2(\u_cpu.ALU._0389_ ),
    .B1(\u_cpu.ALU._1287_ ),
    .B2(\u_cpu.ALU._0393_ ),
    .X(\u_cpu.ALU._0394_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.ALU._2620_  (.A(\u_cpu.ALU._0387_ ),
    .B(\u_cpu.ALU._0388_ ),
    .C(\u_cpu.ALU._0394_ ),
    .X(\u_cpu.ALU._0395_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU._2621_  (.A1(\u_cpu.ALU._0381_ ),
    .A2(\u_cpu.ALU._0385_ ),
    .A3(\u_cpu.ALU._0144_ ),
    .B1(\u_cpu.ALU._0395_ ),
    .Y(\u_cpu.ALU._0396_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._2622_  (.A(\u_cpu.ALU._0396_ ),
    .Y(\u_cpu.ALU.ALUResult[27] ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU._2623_  (.A1(\u_cpu.ALU._0358_ ),
    .A2(\u_cpu.ALU._0361_ ),
    .B1(\u_cpu.ALU._0378_ ),
    .B2(\u_cpu.ALU._0379_ ),
    .C1(\u_cpu.ALU._0363_ ),
    .X(\u_cpu.ALU._0397_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU._2624_  (.A_N(\u_cpu.ALU._0331_ ),
    .B(\u_cpu.ALU._0397_ ),
    .C(\u_cpu.ALU._0297_ ),
    .D(\u_cpu.ALU._0298_ ),
    .Y(\u_cpu.ALU._0398_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU._2625_  (.A1(\u_cpu.ALU._0306_ ),
    .A2(\u_cpu.ALU._0314_ ),
    .B1_N(\u_cpu.ALU._0398_ ),
    .Y(\u_cpu.ALU._0399_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2626_  (.A1(\u_cpu.ALU._0378_ ),
    .A2(\u_cpu.ALU._0379_ ),
    .B1(\u_cpu.ALU._0364_ ),
    .Y(\u_cpu.ALU._0400_ ));
 sky130_fd_sc_hd__a32oi_2 \u_cpu.ALU._2627_  (.A1(\u_cpu.ALU._0359_ ),
    .A2(\u_cpu.ALU._0376_ ),
    .A3(\u_cpu.ALU._0377_ ),
    .B1(\u_cpu.ALU._0383_ ),
    .B2(\u_cpu.ALU._0363_ ),
    .Y(\u_cpu.ALU._0402_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.ALU._2628_  (.A1(\u_cpu.ALU._0368_ ),
    .A2(\u_cpu.ALU._0400_ ),
    .B1_N(\u_cpu.ALU._0402_ ),
    .X(\u_cpu.ALU._0403_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU._2629_  (.A1(\u_cpu.ALU._0900_ ),
    .A2(\u_cpu.ALU._0921_ ),
    .B1(\u_cpu.ALU.SrcB[27] ),
    .B2(\u_cpu.ALU._0375_ ),
    .C1(\u_cpu.ALU._0582_ ),
    .X(\u_cpu.ALU._0404_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU._2630_  (.A(\u_cpu.ALU._0244_ ),
    .B(\u_cpu.ALU._0291_ ),
    .C(\u_cpu.ALU._0374_ ),
    .D(\u_cpu.ALU._0370_ ),
    .Y(\u_cpu.ALU._0405_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2631_  (.A1(\u_cpu.ALU._0160_ ),
    .A2(\u_cpu.ALU._0405_ ),
    .B1(\u_cpu.ALU._0582_ ),
    .Y(\u_cpu.ALU._0406_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU._2632_  (.A(\u_cpu.ALU._0581_ ),
    .B(\u_cpu.ALU._0406_ ),
    .X(\u_cpu.ALU._0407_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2633_  (.A1(\u_cpu.ALU._0406_ ),
    .A2(\u_cpu.ALU._0404_ ),
    .B1(\u_cpu.ALU._0581_ ),
    .Y(\u_cpu.ALU._0408_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2634_  (.A1(\u_cpu.ALU._0404_ ),
    .A2(\u_cpu.ALU._0407_ ),
    .B1(\u_cpu.ALU._0408_ ),
    .Y(\u_cpu.ALU._0409_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2635_  (.A1(\u_cpu.ALU._0399_ ),
    .A2(\u_cpu.ALU._0403_ ),
    .B1(\u_cpu.ALU._0409_ ),
    .X(\u_cpu.ALU._0410_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._2636_  (.A1(\u_cpu.ALU._0398_ ),
    .A2(\u_cpu.ALU._0354_ ),
    .B1(\u_cpu.ALU._0409_ ),
    .C1(\u_cpu.ALU._0403_ ),
    .Y(\u_cpu.ALU._0411_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU._2637_  (.A(\u_cpu.ALU._0410_ ),
    .B(\u_cpu.ALU._0144_ ),
    .C(\u_cpu.ALU._0411_ ),
    .Y(\u_cpu.ALU._0413_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2638_  (.A0(\u_cpu.ALU._0581_ ),
    .A1(\u_cpu.ALU._0338_ ),
    .A2(\u_cpu.ALU.SrcA[26] ),
    .A3(\u_cpu.ALU._0475_ ),
    .S0(\u_cpu.ALU._0723_ ),
    .S1(\u_cpu.ALU._0899_ ),
    .X(\u_cpu.ALU._0414_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2639_  (.A0(\u_cpu.ALU._0090_ ),
    .A1(\u_cpu.ALU._0202_ ),
    .A2(\u_cpu.ALU._0321_ ),
    .A3(\u_cpu.ALU._0414_ ),
    .S0(\u_cpu.ALU._1279_ ),
    .S1(\u_cpu.ALU._1212_ ),
    .X(\u_cpu.ALU._0415_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.ALU._2640_  (.A0(\u_cpu.ALU._0415_ ),
    .A1(\u_cpu.ALU._1322_ ),
    .S(\u_cpu.ALU._1144_ ),
    .X(\u_cpu.ALU._0416_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU._2641_  (.A(\u_cpu.ALU._1158_ ),
    .B(\u_cpu.ALU._1075_ ),
    .C(\u_cpu.ALU._1149_ ),
    .X(\u_cpu.ALU._0417_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2642_  (.A1(\u_cpu.ALU._1316_ ),
    .A2(\u_cpu.ALU._1317_ ),
    .B1(\u_cpu.ALU._0879_ ),
    .X(\u_cpu.ALU._0418_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2643_  (.A1(\u_cpu.ALU._1144_ ),
    .A2(\u_cpu.ALU._0577_ ),
    .B1(\u_cpu.ALU._0418_ ),
    .X(\u_cpu.ALU._0419_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU._2644_  (.A(\u_cpu.ALU._0737_ ),
    .B(\u_cpu.ALU._0520_ ),
    .C(\u_cpu.ALU._0900_ ),
    .D(\u_cpu.ALU._0890_ ),
    .X(\u_cpu.ALU._0420_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU._2645_  (.A1(\u_cpu.ALU._0581_ ),
    .A2(\u_cpu.ALU._0582_ ),
    .B1(\u_cpu.ALU._0748_ ),
    .B2(\u_cpu.ALU._0420_ ),
    .X(\u_cpu.ALU._0421_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2646_  (.A1(\u_cpu.ALU._0582_ ),
    .A2(\u_cpu.ALU._0754_ ),
    .B1(\u_cpu.ALU._0822_ ),
    .B2(\u_cpu.ALU.Product_Wallace[28] ),
    .C1(\u_cpu.ALU._0421_ ),
    .X(\u_cpu.ALU._0422_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU._2647_  (.A1(\u_cpu.ALU._0581_ ),
    .A2(\u_cpu.ALU._0582_ ),
    .A3(\u_cpu.ALU._0058_ ),
    .B1(\u_cpu.ALU._0422_ ),
    .X(\u_cpu.ALU._0424_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2648_  (.A1(\u_cpu.ALU._1316_ ),
    .A2(\u_cpu.ALU._0417_ ),
    .B1(\u_cpu.ALU._0419_ ),
    .B2(\u_cpu.ALU._0874_ ),
    .C1(\u_cpu.ALU._0424_ ),
    .X(\u_cpu.ALU._0425_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2649_  (.A1(\u_cpu.ALU._0026_ ),
    .A2(\u_cpu.ALU._0416_ ),
    .B1(\u_cpu.ALU._0425_ ),
    .Y(\u_cpu.ALU._0426_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2650_  (.A(\u_cpu.ALU._0413_ ),
    .B(\u_cpu.ALU._0426_ ),
    .Y(\u_cpu.ALU.ALUResult[28] ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2651_  (.A1(\u_cpu.ALU._0406_ ),
    .A2(\u_cpu.ALU._0404_ ),
    .B1(\u_cpu.ALU._0581_ ),
    .X(\u_cpu.ALU._0427_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2652_  (.A1(\u_cpu.ALU._0399_ ),
    .A2(\u_cpu.ALU._0403_ ),
    .B1(\u_cpu.ALU._0409_ ),
    .Y(\u_cpu.ALU._0428_ ));
 sky130_fd_sc_hd__or4bb_2 \u_cpu.ALU._2653_  (.A(\u_cpu.ALU._0582_ ),
    .B(\u_cpu.ALU._0292_ ),
    .C_N(\u_cpu.ALU._0374_ ),
    .D_N(\u_cpu.ALU._0370_ ),
    .X(\u_cpu.ALU._0429_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2654_  (.A1(\u_cpu.ALU._0160_ ),
    .A2(\u_cpu.ALU._0429_ ),
    .B1(\u_cpu.ALU.SrcB[29] ),
    .Y(\u_cpu.ALU._0430_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU._2655_  (.A1(\u_cpu.ALU._0582_ ),
    .A2(\u_cpu.ALU.SrcB[27] ),
    .A3(\u_cpu.ALU._0375_ ),
    .B1(\u_cpu.ALU._0160_ ),
    .C1(\u_cpu.ALU.SrcB[29] ),
    .X(\u_cpu.ALU._0431_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2656_  (.A1(\u_cpu.ALU._0430_ ),
    .A2(\u_cpu.ALU._0431_ ),
    .B1(\u_cpu.ALU._0579_ ),
    .X(\u_cpu.ALU._0432_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU._2657_  (.A(\u_cpu.ALU._0579_ ),
    .B(\u_cpu.ALU._0430_ ),
    .C(\u_cpu.ALU._0431_ ),
    .Y(\u_cpu.ALU._0434_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU._2658_  (.A(\u_cpu.ALU._0432_ ),
    .B(\u_cpu.ALU._0434_ ),
    .X(\u_cpu.ALU._0435_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU._2659_  (.A1(\u_cpu.ALU._0427_ ),
    .A2(\u_cpu.ALU._0428_ ),
    .B1_N(\u_cpu.ALU._0435_ ),
    .Y(\u_cpu.ALU._0436_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2660_  (.A1(\u_cpu.ALU._0398_ ),
    .A2(\u_cpu.ALU._0354_ ),
    .B1(\u_cpu.ALU._0403_ ),
    .X(\u_cpu.ALU._0437_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU._2661_  (.A1(\u_cpu.ALU._0432_ ),
    .A2(\u_cpu.ALU._0434_ ),
    .B1(\u_cpu.ALU._0409_ ),
    .B2(\u_cpu.ALU._0437_ ),
    .C1(\u_cpu.ALU._0408_ ),
    .Y(\u_cpu.ALU._0438_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2662_  (.A0(\u_cpu.ALU._0579_ ),
    .A1(\u_cpu.ALU._0581_ ),
    .A2(\u_cpu.ALU._0338_ ),
    .A3(\u_cpu.ALU.SrcA[26] ),
    .S0(\u_cpu.ALU._0723_ ),
    .S1(\u_cpu.ALU._0899_ ),
    .X(\u_cpu.ALU._0439_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2663_  (.A0(\u_cpu.ALU._0110_ ),
    .A1(\u_cpu.ALU._0230_ ),
    .A2(\u_cpu.ALU._0337_ ),
    .A3(\u_cpu.ALU._0439_ ),
    .S0(\u_cpu.ALU._1279_ ),
    .S1(\u_cpu.ALU._1212_ ),
    .X(\u_cpu.ALU._0440_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU._2664_  (.A1(\u_cpu.ALU._0819_ ),
    .A2(\u_cpu.ALU._1333_ ),
    .B1(\u_cpu.ALU._0440_ ),
    .B2(\u_cpu.ALU._1283_ ),
    .Y(\u_cpu.ALU._0441_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2665_  (.A(\u_cpu.ALU._0521_ ),
    .B(\u_cpu.ALU._0522_ ),
    .Y(\u_cpu.ALU._0442_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2666_  (.A1(\u_cpu.ALU._0579_ ),
    .A2(\u_cpu.ALU.SrcB[29] ),
    .B1(\u_cpu.ALU._0061_ ),
    .C1(\u_cpu.ALU._1331_ ),
    .D1(\u_cpu.ALU._1332_ ),
    .X(\u_cpu.ALU._0443_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2667_  (.A1(\u_cpu.ALU._0522_ ),
    .A2(\u_cpu.ALU._0058_ ),
    .B1(\u_cpu.ALU._0813_ ),
    .B2(\u_cpu.ALU._0442_ ),
    .C1(\u_cpu.ALU._0443_ ),
    .X(\u_cpu.ALU._0445_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2668_  (.A1(\u_cpu.ALU.SrcB[29] ),
    .A2(\u_cpu.ALU._0060_ ),
    .B1(\u_cpu.ALU._1338_ ),
    .B2(\u_cpu.ALU.Product_Wallace[29] ),
    .C1(\u_cpu.ALU._0115_ ),
    .X(\u_cpu.ALU._0446_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2669_  (.A(\u_cpu.ALU._0445_ ),
    .B(\u_cpu.ALU._0446_ ),
    .Y(\u_cpu.ALU._0447_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU._2670_  (.A1(\u_cpu.ALU._1283_ ),
    .A2(\u_cpu.ALU._1337_ ),
    .B1(\u_cpu.ALU._0441_ ),
    .C1(\u_cpu.ALU._0447_ ),
    .Y(\u_cpu.ALU._0448_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU._2671_  (.A1(\u_cpu.ALU._0436_ ),
    .A2(\u_cpu.ALU._0438_ ),
    .A3(\u_cpu.ALU._0144_ ),
    .B1(\u_cpu.ALU._0448_ ),
    .Y(\u_cpu.ALU._0449_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._2672_  (.A(\u_cpu.ALU._0449_ ),
    .Y(\u_cpu.ALU.ALUResult[29] ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.ALU._2673_  (.A1(\u_cpu.ALU._0579_ ),
    .A2(\u_cpu.ALU._0430_ ),
    .A3(\u_cpu.ALU._0431_ ),
    .B1(\u_cpu.ALU._0432_ ),
    .B2(\u_cpu.ALU._0427_ ),
    .X(\u_cpu.ALU._0450_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.ALU._2674_  (.A(\u_cpu.ALU._0432_ ),
    .B(\u_cpu.ALU._0434_ ),
    .C(\u_cpu.ALU._0409_ ),
    .X(\u_cpu.ALU._0451_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2675_  (.A1(\u_cpu.ALU._0399_ ),
    .A2(\u_cpu.ALU._0403_ ),
    .B1(\u_cpu.ALU._0451_ ),
    .Y(\u_cpu.ALU._0452_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.ALU._2676_  (.A1(\u_cpu.ALU.SrcB[29] ),
    .A2(\u_cpu.ALU._0582_ ),
    .A3(\u_cpu.ALU._0405_ ),
    .B1(\u_cpu.ALU._0921_ ),
    .B2(\u_cpu.ALU._1149_ ),
    .X(\u_cpu.ALU._0453_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu.ALU._2677_  (.A(\u_cpu.ALU.SrcB[30] ),
    .B(\u_cpu.ALU._0453_ ),
    .Y(\u_cpu.ALU._0455_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu.ALU._2678_  (.A(\u_cpu.ALU._0516_ ),
    .B(\u_cpu.ALU._0455_ ),
    .Y(\u_cpu.ALU._0456_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU._2679_  (.A1(\u_cpu.ALU._0450_ ),
    .A2(\u_cpu.ALU._0452_ ),
    .B1_N(\u_cpu.ALU._0456_ ),
    .Y(\u_cpu.ALU._0457_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2680_  (.A(\u_cpu.ALU._0427_ ),
    .B(\u_cpu.ALU._0432_ ),
    .Y(\u_cpu.ALU._0458_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU._2681_  (.A1(\u_cpu.ALU._0434_ ),
    .A2(\u_cpu.ALU._0458_ ),
    .B1(\u_cpu.ALU._0451_ ),
    .B2(\u_cpu.ALU._0437_ ),
    .C1(\u_cpu.ALU._0456_ ),
    .Y(\u_cpu.ALU._0459_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2682_  (.A0(\u_cpu.ALU._0516_ ),
    .A1(\u_cpu.ALU._0579_ ),
    .A2(\u_cpu.ALU._0581_ ),
    .A3(\u_cpu.ALU._0338_ ),
    .S0(\u_cpu.ALU._0723_ ),
    .S1(\u_cpu.ALU._0899_ ),
    .X(\u_cpu.ALU._0460_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2683_  (.A0(\u_cpu.ALU._0151_ ),
    .A1(\u_cpu.ALU._0254_ ),
    .A2(\u_cpu.ALU._0346_ ),
    .A3(\u_cpu.ALU._0460_ ),
    .S0(\u_cpu.ALU._1279_ ),
    .S1(\u_cpu.ALU._1212_ ),
    .X(\u_cpu.ALU._0461_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.ALU._2684_  (.A0(\u_cpu.ALU._0025_ ),
    .A1(\u_cpu.ALU._0461_ ),
    .S(\u_cpu.ALU._1275_ ),
    .X(\u_cpu.ALU._0462_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2685_  (.A1(\u_cpu.ALU._0516_ ),
    .A2(\u_cpu.ALU.SrcB[30] ),
    .B1(\u_cpu.ALU._1020_ ),
    .Y(\u_cpu.ALU._0463_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU._2686_  (.A1(\u_cpu.ALU._0516_ ),
    .A2(\u_cpu.ALU.SrcB[30] ),
    .B1(\u_cpu.ALU._0749_ ),
    .B2(\u_cpu.ALU._0463_ ),
    .X(\u_cpu.ALU._0464_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU._2687_  (.A1(\u_cpu.ALU._0957_ ),
    .A2(\u_cpu.ALU._0516_ ),
    .B1(\u_cpu.ALU.SrcB[30] ),
    .C1(\u_cpu.ALU._0896_ ),
    .X(\u_cpu.ALU._0466_ ));
 sky130_fd_sc_hd__a2111oi_2 \u_cpu.ALU._2688_  (.A1(\u_cpu.ALU.Product_Wallace[30] ),
    .A2(\u_cpu.ALU._1338_ ),
    .B1(\u_cpu.ALU._0115_ ),
    .C1(\u_cpu.ALU._0464_ ),
    .D1(\u_cpu.ALU._0466_ ),
    .Y(\u_cpu.ALU._0467_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU._2689_  (.A1(\u_cpu.ALU._1283_ ),
    .A2(\u_cpu.ALU._0034_ ),
    .B1(\u_cpu.ALU._0467_ ),
    .Y(\u_cpu.ALU._0468_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU._2690_  (.A1(\u_cpu.ALU._0462_ ),
    .A2(\u_cpu.ALU._0026_ ),
    .B1(\u_cpu.ALU._0468_ ),
    .X(\u_cpu.ALU._0469_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU._2691_  (.A1(\u_cpu.ALU._0457_ ),
    .A2(\u_cpu.ALU._0459_ ),
    .A3(\u_cpu.ALU._0144_ ),
    .B1(\u_cpu.ALU._0469_ ),
    .Y(\u_cpu.ALU._0470_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._2692_  (.A(\u_cpu.ALU._0470_ ),
    .Y(\u_cpu.ALU.ALUResult[30] ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2693_  (.A(\u_cpu.ALU._0455_ ),
    .B(\u_cpu.ALU._0516_ ),
    .Y(\u_cpu.ALU._0471_ ));
 sky130_fd_sc_hd__nor4_2 \u_cpu.ALU._2694_  (.A(\u_cpu.ALU.SrcB[30] ),
    .B(\u_cpu.ALU.SrcB[29] ),
    .C(\u_cpu.ALU._0582_ ),
    .D(\u_cpu.ALU._0405_ ),
    .Y(\u_cpu.ALU._0472_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU._2695_  (.A1(\u_cpu.ALU._1200_ ),
    .A2(\u_cpu.ALU._0472_ ),
    .B1(\u_cpu.ALU._0526_ ),
    .X(\u_cpu.ALU._0473_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU._2696_  (.A1(\u_cpu.ALU.SrcB[30] ),
    .A2(\u_cpu.ALU.SrcB[29] ),
    .A3(\u_cpu.ALU._0429_ ),
    .B1(\u_cpu.ALU._0160_ ),
    .C1(\u_cpu.ALU._0527_ ),
    .X(\u_cpu.ALU._0474_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU._2697_  (.A(\u_cpu.ALU._0473_ ),
    .B(\u_cpu.ALU._0474_ ),
    .X(\u_cpu.ALU._0476_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU._2698_  (.A1(\u_cpu.ALU._0471_ ),
    .A2(\u_cpu.ALU._0457_ ),
    .B1(\u_cpu.ALU._0476_ ),
    .Y(\u_cpu.ALU._0477_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU._2699_  (.A(\u_cpu.ALU._0434_ ),
    .Y(\u_cpu.ALU._0478_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU._2700_  (.A(\u_cpu.ALU._0427_ ),
    .B(\u_cpu.ALU._0432_ ),
    .X(\u_cpu.ALU._0479_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU._2701_  (.A1(\u_cpu.ALU._0368_ ),
    .A2(\u_cpu.ALU._0400_ ),
    .B1_N(\u_cpu.ALU._0402_ ),
    .Y(\u_cpu.ALU._0480_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU._2702_  (.A1(\u_cpu.ALU._0398_ ),
    .A2(\u_cpu.ALU._0354_ ),
    .B1_N(\u_cpu.ALU._0480_ ),
    .Y(\u_cpu.ALU._0481_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU._2703_  (.A(\u_cpu.ALU._0409_ ),
    .B(\u_cpu.ALU._0435_ ),
    .Y(\u_cpu.ALU._0482_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU._2704_  (.A1(\u_cpu.ALU._0478_ ),
    .A2(\u_cpu.ALU._0479_ ),
    .B1(\u_cpu.ALU._0481_ ),
    .B2(\u_cpu.ALU._0482_ ),
    .Y(\u_cpu.ALU._0483_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU._2705_  (.A1(\u_cpu.ALU._0473_ ),
    .A2(\u_cpu.ALU._0474_ ),
    .B1(\u_cpu.ALU._0456_ ),
    .B2(\u_cpu.ALU._0483_ ),
    .C1(\u_cpu.ALU._0471_ ),
    .Y(\u_cpu.ALU._0484_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU._2706_  (.A(\u_cpu.ALU._0484_ ),
    .B(\u_cpu.ALU._0144_ ),
    .Y(\u_cpu.ALU._0485_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU._2707_  (.A1(\u_cpu.ALU._0524_ ),
    .A2(\u_cpu.ALU._0058_ ),
    .B1(\u_cpu.ALU._0060_ ),
    .B2(\u_cpu.ALU.SrcB[31] ),
    .X(\u_cpu.ALU._0487_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU._2708_  (.A1(\u_cpu.ALU.Product_Wallace[31] ),
    .A2(\u_cpu.ALU._1338_ ),
    .B1(\u_cpu.ALU._0874_ ),
    .B2(\u_cpu.ALU._0577_ ),
    .C1(\u_cpu.ALU._0487_ ),
    .X(\u_cpu.ALU._0488_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2709_  (.A0(\u_cpu.ALU.SrcA[31] ),
    .A1(\u_cpu.ALU._0516_ ),
    .A2(\u_cpu.ALU._0579_ ),
    .A3(\u_cpu.ALU._0581_ ),
    .S0(\u_cpu.ALU._0723_ ),
    .S1(\u_cpu.ALU._0899_ ),
    .X(\u_cpu.ALU._0489_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.ALU._2710_  (.A0(\u_cpu.ALU._0176_ ),
    .A1(\u_cpu.ALU._0277_ ),
    .A2(\u_cpu.ALU._0390_ ),
    .A3(\u_cpu.ALU._0489_ ),
    .S0(\u_cpu.ALU._0786_ ),
    .S1(\u_cpu.ALU._1219_ ),
    .X(\u_cpu.ALU._0490_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.ALU._2711_  (.A0(\u_cpu.ALU._0053_ ),
    .A1(\u_cpu.ALU._0490_ ),
    .S(\u_cpu.ALU._1075_ ),
    .X(\u_cpu.ALU._0491_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU._2712_  (.A1(\u_cpu.ALU._0994_ ),
    .A2(\u_cpu.ALU._0576_ ),
    .B1(\u_cpu.ALU._0738_ ),
    .C1(\u_cpu.ALU._1149_ ),
    .D1(\u_cpu.ALU._0890_ ),
    .X(\u_cpu.ALU._0492_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU._2713_  (.A1(\u_cpu.ALU._0577_ ),
    .A2(\u_cpu.ALU.SrcB[31] ),
    .B1(\u_cpu.ALU._0749_ ),
    .B2(\u_cpu.ALU._0492_ ),
    .X(\u_cpu.ALU._0493_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU._2714_  (.A1(\u_cpu.ALU._0491_ ),
    .A2(\u_cpu.ALU._0738_ ),
    .A3(\u_cpu.ALU._1331_ ),
    .A4(\u_cpu.ALU._1332_ ),
    .B1(\u_cpu.ALU._0493_ ),
    .X(\u_cpu.ALU._0494_ ));
 sky130_fd_sc_hd__a311o_2 \u_cpu.ALU._2715_  (.A1(\u_cpu.ALU._0577_ ),
    .A2(\u_cpu.ALU._0801_ ),
    .A3(\u_cpu.ALU._0417_ ),
    .B1(\u_cpu.ALU._0488_ ),
    .C1(\u_cpu.ALU._0494_ ),
    .X(\u_cpu.ALU._0495_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU._2716_  (.A1(\u_cpu.ALU._0477_ ),
    .A2(\u_cpu.ALU._0485_ ),
    .B1_N(\u_cpu.ALU._0495_ ),
    .Y(\u_cpu.ALU.ALUResult[31] ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._4935_  (.A(\u_cpu.ALU.SrcB[0] ),
    .Y(\u_cpu.ALU.u_wallace._4912_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4936_  (.A(\u_cpu.ALU.u_wallace._4912_ ),
    .X(\u_cpu.ALU.u_wallace._4923_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4937_  (.A(\u_cpu.ALU.u_wallace._4923_ ),
    .X(\u_cpu.ALU.u_wallace._4934_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4938_  (.A(\u_cpu.ALU.SrcA[0] ),
    .X(\u_cpu.ALU.u_wallace._0010_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4939_  (.A(\u_cpu.ALU.u_wallace._0010_ ),
    .X(\u_cpu.ALU.u_wallace._0021_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._4940_  (.A(\u_cpu.ALU.u_wallace._0021_ ),
    .Y(\u_cpu.ALU.u_wallace._0032_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4941_  (.A(\u_cpu.ALU.u_wallace._0032_ ),
    .X(\u_cpu.ALU.u_wallace._0043_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._4942_  (.A(\u_cpu.ALU.u_wallace._4934_ ),
    .B(\u_cpu.ALU.u_wallace._0043_ ),
    .Y(\u_cpu.ALU.Product_Wallace[0] ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4943_  (.A(\u_cpu.ALU.SrcB[0] ),
    .X(\u_cpu.ALU.u_wallace._0064_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4944_  (.A(\u_cpu.ALU.u_wallace._0064_ ),
    .X(\u_cpu.ALU.u_wallace._0075_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4945_  (.A(\u_cpu.ALU.u_wallace._0075_ ),
    .X(\u_cpu.ALU.u_wallace._0086_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4946_  (.A(\u_cpu.ALU.u_wallace._0086_ ),
    .X(\u_cpu.ALU.u_wallace._0097_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4947_  (.A(\u_cpu.ALU.u_wallace._0021_ ),
    .X(\u_cpu.ALU.u_wallace._0108_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4948_  (.A(\u_cpu.ALU.u_wallace._0108_ ),
    .X(\u_cpu.ALU.u_wallace._0118_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4949_  (.A(\u_cpu.ALU.u_wallace._0118_ ),
    .X(\u_cpu.ALU.u_wallace._0129_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4950_  (.A(\u_cpu.ALU.SrcA[1] ),
    .X(\u_cpu.ALU.u_wallace._0140_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4951_  (.A(\u_cpu.ALU.u_wallace._0140_ ),
    .X(\u_cpu.ALU.u_wallace._0151_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4952_  (.A(\u_cpu.ALU.u_wallace._0151_ ),
    .X(\u_cpu.ALU.u_wallace._0162_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4953_  (.A(\u_cpu.ALU.u_wallace._0162_ ),
    .X(\u_cpu.ALU.u_wallace._0173_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4954_  (.A(\u_cpu.ALU.u_wallace._0173_ ),
    .X(\u_cpu.ALU.u_wallace._0184_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4955_  (.A(\u_cpu.ALU.SrcB[1] ),
    .X(\u_cpu.ALU.u_wallace._0195_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4956_  (.A(\u_cpu.ALU.u_wallace._0195_ ),
    .X(\u_cpu.ALU.u_wallace._0206_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4957_  (.A(\u_cpu.ALU.u_wallace._0206_ ),
    .X(\u_cpu.ALU.u_wallace._0217_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4958_  (.A(\u_cpu.ALU.u_wallace._0217_ ),
    .X(\u_cpu.ALU.u_wallace._0228_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._4959_  (.A(\u_cpu.ALU.u_wallace._0097_ ),
    .B(\u_cpu.ALU.u_wallace._0129_ ),
    .C(\u_cpu.ALU.u_wallace._0184_ ),
    .D(\u_cpu.ALU.u_wallace._0228_ ),
    .Y(\u_cpu.ALU.u_wallace._0239_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4960_  (.A(\u_cpu.ALU.SrcA[1] ),
    .X(\u_cpu.ALU.u_wallace._0250_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4961_  (.A(\u_cpu.ALU.u_wallace._0250_ ),
    .X(\u_cpu.ALU.u_wallace._0261_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4962_  (.A(\u_cpu.ALU.u_wallace._0261_ ),
    .X(\u_cpu.ALU.u_wallace._0272_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4963_  (.A(\u_cpu.ALU.SrcB[2] ),
    .X(\u_cpu.ALU.u_wallace._0282_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4964_  (.A(\u_cpu.ALU.u_wallace._0282_ ),
    .X(\u_cpu.ALU.u_wallace._0293_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4965_  (.A(\u_cpu.ALU.u_wallace._0293_ ),
    .X(\u_cpu.ALU.u_wallace._0304_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4966_  (.A(\u_cpu.ALU.u_wallace._0304_ ),
    .X(\u_cpu.ALU.u_wallace._0315_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._4967_  (.A(\u_cpu.ALU.u_wallace._0118_ ),
    .B(\u_cpu.ALU.u_wallace._0272_ ),
    .C(\u_cpu.ALU.u_wallace._0228_ ),
    .D(\u_cpu.ALU.u_wallace._0315_ ),
    .X(\u_cpu.ALU.u_wallace._0326_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._4968_  (.A1(\u_cpu.ALU.u_wallace._0173_ ),
    .A2(\u_cpu.ALU.u_wallace._0228_ ),
    .B1(\u_cpu.ALU.u_wallace._0315_ ),
    .B2(\u_cpu.ALU.u_wallace._0118_ ),
    .X(\u_cpu.ALU.u_wallace._0337_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4969_  (.A(\u_cpu.ALU.SrcA[2] ),
    .X(\u_cpu.ALU.u_wallace._0348_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4970_  (.A(\u_cpu.ALU.u_wallace._0348_ ),
    .X(\u_cpu.ALU.u_wallace._0359_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4971_  (.A(\u_cpu.ALU.u_wallace._0359_ ),
    .X(\u_cpu.ALU.u_wallace._0370_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.ALU.u_wallace._4972_  (.A_N(\u_cpu.ALU.u_wallace._0326_ ),
    .B(\u_cpu.ALU.u_wallace._0337_ ),
    .C(\u_cpu.ALU.u_wallace._0097_ ),
    .D(\u_cpu.ALU.u_wallace._0370_ ),
    .X(\u_cpu.ALU.u_wallace._0381_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4973_  (.A(\u_cpu.ALU.SrcA[2] ),
    .X(\u_cpu.ALU.u_wallace._0392_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._4974_  (.A(\u_cpu.ALU.u_wallace._0392_ ),
    .Y(\u_cpu.ALU.u_wallace._0403_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4975_  (.A(\u_cpu.ALU.u_wallace._0403_ ),
    .X(\u_cpu.ALU.u_wallace._0414_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._4976_  (.A1(\u_cpu.ALU.u_wallace._0184_ ),
    .A2(\u_cpu.ALU.u_wallace._0228_ ),
    .B1(\u_cpu.ALU.u_wallace._0315_ ),
    .B2(\u_cpu.ALU.u_wallace._0129_ ),
    .Y(\u_cpu.ALU.u_wallace._0425_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._4977_  (.A1(\u_cpu.ALU.u_wallace._4934_ ),
    .A2(\u_cpu.ALU.u_wallace._0414_ ),
    .B1(\u_cpu.ALU.u_wallace._0326_ ),
    .B2(\u_cpu.ALU.u_wallace._0425_ ),
    .X(\u_cpu.ALU.u_wallace._0435_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4978_  (.A(\u_cpu.ALU.u_wallace._0010_ ),
    .X(\u_cpu.ALU.u_wallace._0446_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4979_  (.A(\u_cpu.ALU.SrcB[3] ),
    .X(\u_cpu.ALU.u_wallace._0457_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4980_  (.A(\u_cpu.ALU.u_wallace._0457_ ),
    .X(\u_cpu.ALU.u_wallace._0468_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4981_  (.A(\u_cpu.ALU.u_wallace._0195_ ),
    .X(\u_cpu.ALU.u_wallace._0479_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4982_  (.A(\u_cpu.ALU.u_wallace._0282_ ),
    .X(\u_cpu.ALU.u_wallace._0490_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._4983_  (.A1(\u_cpu.ALU.u_wallace._0348_ ),
    .A2(\u_cpu.ALU.u_wallace._0479_ ),
    .B1(\u_cpu.ALU.u_wallace._0490_ ),
    .B2(\u_cpu.ALU.u_wallace._0140_ ),
    .X(\u_cpu.ALU.u_wallace._0501_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4984_  (.A(\u_cpu.ALU.SrcA[2] ),
    .X(\u_cpu.ALU.u_wallace._0512_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4985_  (.A(\u_cpu.ALU.u_wallace._0195_ ),
    .X(\u_cpu.ALU.u_wallace._0523_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4986_  (.A(\u_cpu.ALU.u_wallace._0282_ ),
    .X(\u_cpu.ALU.u_wallace._0534_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4987_  (.A(\u_cpu.ALU.u_wallace._0534_ ),
    .X(\u_cpu.ALU.u_wallace._0545_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._4988_  (.A(\u_cpu.ALU.u_wallace._0512_ ),
    .B(\u_cpu.ALU.u_wallace._0250_ ),
    .C(\u_cpu.ALU.u_wallace._0523_ ),
    .D(\u_cpu.ALU.u_wallace._0545_ ),
    .Y(\u_cpu.ALU.u_wallace._0556_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._4989_  (.A1(\u_cpu.ALU.u_wallace._0446_ ),
    .A2(\u_cpu.ALU.u_wallace._0468_ ),
    .B1(\u_cpu.ALU.u_wallace._0501_ ),
    .B2(\u_cpu.ALU.u_wallace._0556_ ),
    .X(\u_cpu.ALU.u_wallace._0567_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4990_  (.A(\u_cpu.ALU.u_wallace._0457_ ),
    .X(\u_cpu.ALU.u_wallace._0578_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._4991_  (.A(\u_cpu.ALU.u_wallace._0501_ ),
    .B(\u_cpu.ALU.u_wallace._0556_ ),
    .C(\u_cpu.ALU.u_wallace._0446_ ),
    .D(\u_cpu.ALU.u_wallace._0578_ ),
    .Y(\u_cpu.ALU.u_wallace._0589_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4992_  (.A(\u_cpu.ALU.SrcA[3] ),
    .X(\u_cpu.ALU.u_wallace._0600_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._4993_  (.A(\u_cpu.ALU.u_wallace._0600_ ),
    .Y(\u_cpu.ALU.u_wallace._0610_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._4994_  (.A(\u_cpu.ALU.u_wallace._0610_ ),
    .X(\u_cpu.ALU.u_wallace._0621_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._4995_  (.A(\u_cpu.ALU.u_wallace._4934_ ),
    .B(\u_cpu.ALU.u_wallace._0621_ ),
    .Y(\u_cpu.ALU.u_wallace._0632_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._4996_  (.A(\u_cpu.ALU.u_wallace._0567_ ),
    .B(\u_cpu.ALU.u_wallace._0589_ ),
    .C(\u_cpu.ALU.u_wallace._0632_ ),
    .X(\u_cpu.ALU.u_wallace._0643_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU.u_wallace._4997_  (.A1_N(\u_cpu.ALU.u_wallace._0567_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0589_ ),
    .B1(\u_cpu.ALU.u_wallace._4934_ ),
    .B2(\u_cpu.ALU.u_wallace._0621_ ),
    .X(\u_cpu.ALU.u_wallace._0654_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._4998_  (.A(\u_cpu.ALU.u_wallace._0643_ ),
    .B(\u_cpu.ALU.u_wallace._0654_ ),
    .Y(\u_cpu.ALU.u_wallace._0665_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._4999_  (.A1(\u_cpu.ALU.u_wallace._0326_ ),
    .A2(\u_cpu.ALU.u_wallace._0381_ ),
    .B1(\u_cpu.ALU.u_wallace._0665_ ),
    .Y(\u_cpu.ALU.u_wallace._0676_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._5000_  (.A1(\u_cpu.ALU.u_wallace._0337_ ),
    .A2(\u_cpu.ALU.u_wallace._0370_ ),
    .A3(\u_cpu.ALU.u_wallace._0097_ ),
    .B1(\u_cpu.ALU.u_wallace._0326_ ),
    .X(\u_cpu.ALU.u_wallace._0687_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._5001_  (.A1(\u_cpu.ALU.u_wallace._0643_ ),
    .A2(\u_cpu.ALU.u_wallace._0654_ ),
    .B1_N(\u_cpu.ALU.u_wallace._0687_ ),
    .Y(\u_cpu.ALU.u_wallace._0698_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._5002_  (.A(\u_cpu.ALU.u_wallace._0676_ ),
    .B(\u_cpu.ALU.u_wallace._0698_ ),
    .X(\u_cpu.ALU.u_wallace._0709_ ));
 sky130_fd_sc_hd__or4b_2 \u_cpu.ALU.u_wallace._5003_  (.A(\u_cpu.ALU.u_wallace._0239_ ),
    .B(\u_cpu.ALU.u_wallace._0381_ ),
    .C(\u_cpu.ALU.u_wallace._0435_ ),
    .D_N(\u_cpu.ALU.u_wallace._0709_ ),
    .X(\u_cpu.ALU.u_wallace._0720_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5004_  (.A(\u_cpu.ALU.u_wallace._0140_ ),
    .X(\u_cpu.ALU.u_wallace._0731_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5005_  (.A(\u_cpu.ALU.SrcB[3] ),
    .X(\u_cpu.ALU.u_wallace._0742_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5006_  (.A(\u_cpu.ALU.u_wallace._0742_ ),
    .X(\u_cpu.ALU.u_wallace._0753_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5007_  (.A(\u_cpu.ALU.SrcA[3] ),
    .X(\u_cpu.ALU.u_wallace._0764_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5008_  (.A(\u_cpu.ALU.SrcB[1] ),
    .X(\u_cpu.ALU.u_wallace._0775_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5009_  (.A1(\u_cpu.ALU.SrcA[2] ),
    .A2(\u_cpu.ALU.u_wallace._0534_ ),
    .B1(\u_cpu.ALU.u_wallace._0764_ ),
    .B2(\u_cpu.ALU.u_wallace._0775_ ),
    .X(\u_cpu.ALU.u_wallace._0786_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5010_  (.A(\u_cpu.ALU.u_wallace._0195_ ),
    .X(\u_cpu.ALU.u_wallace._0797_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5011_  (.A(\u_cpu.ALU.u_wallace._0282_ ),
    .X(\u_cpu.ALU.u_wallace._0807_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5012_  (.A(\u_cpu.ALU.SrcA[2] ),
    .B(\u_cpu.ALU.u_wallace._0797_ ),
    .C(\u_cpu.ALU.u_wallace._0807_ ),
    .D(\u_cpu.ALU.u_wallace._0764_ ),
    .Y(\u_cpu.ALU.u_wallace._0818_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5013_  (.A1(\u_cpu.ALU.u_wallace._0731_ ),
    .A2(\u_cpu.ALU.u_wallace._0753_ ),
    .B1(\u_cpu.ALU.u_wallace._0786_ ),
    .B2(\u_cpu.ALU.u_wallace._0818_ ),
    .X(\u_cpu.ALU.u_wallace._0829_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5014_  (.A(\u_cpu.ALU.u_wallace._0742_ ),
    .X(\u_cpu.ALU.u_wallace._0840_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5015_  (.A(\u_cpu.ALU.u_wallace._0786_ ),
    .B(\u_cpu.ALU.u_wallace._0818_ ),
    .C(\u_cpu.ALU.u_wallace._0151_ ),
    .D(\u_cpu.ALU.u_wallace._0840_ ),
    .Y(\u_cpu.ALU.u_wallace._0851_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5016_  (.A(\u_cpu.ALU.u_wallace._0064_ ),
    .X(\u_cpu.ALU.u_wallace._0862_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5017_  (.A(\u_cpu.ALU.u_wallace._0862_ ),
    .X(\u_cpu.ALU.u_wallace._0873_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5018_  (.A(\u_cpu.ALU.u_wallace._0873_ ),
    .X(\u_cpu.ALU.u_wallace._0884_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5019_  (.A(\u_cpu.ALU.SrcA[4] ),
    .X(\u_cpu.ALU.u_wallace._0895_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5020_  (.A(\u_cpu.ALU.u_wallace._0895_ ),
    .X(\u_cpu.ALU.u_wallace._0906_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5021_  (.A(\u_cpu.ALU.u_wallace._0906_ ),
    .X(\u_cpu.ALU.u_wallace._0917_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5022_  (.A(\u_cpu.ALU.u_wallace._0829_ ),
    .B(\u_cpu.ALU.u_wallace._0851_ ),
    .C(\u_cpu.ALU.u_wallace._0884_ ),
    .D(\u_cpu.ALU.u_wallace._0917_ ),
    .Y(\u_cpu.ALU.u_wallace._0928_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._5023_  (.A(\u_cpu.ALU.u_wallace._0895_ ),
    .Y(\u_cpu.ALU.u_wallace._0939_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5024_  (.A1_N(\u_cpu.ALU.u_wallace._0829_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0851_ ),
    .B1(\u_cpu.ALU.u_wallace._4934_ ),
    .B2(\u_cpu.ALU.u_wallace._0939_ ),
    .Y(\u_cpu.ALU.u_wallace._0950_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._5025_  (.A1(\u_cpu.ALU.u_wallace._0632_ ),
    .A2(\u_cpu.ALU.u_wallace._0567_ ),
    .A3(\u_cpu.ALU.u_wallace._0589_ ),
    .B1(\u_cpu.ALU.u_wallace._0928_ ),
    .B2(\u_cpu.ALU.u_wallace._0950_ ),
    .X(\u_cpu.ALU.u_wallace._0961_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5026_  (.A(\u_cpu.ALU.u_wallace._0643_ ),
    .B(\u_cpu.ALU.u_wallace._0928_ ),
    .C(\u_cpu.ALU.u_wallace._0950_ ),
    .Y(\u_cpu.ALU.u_wallace._0972_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5027_  (.A(\u_cpu.ALU.u_wallace._0753_ ),
    .X(\u_cpu.ALU.u_wallace._0983_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5028_  (.A(\u_cpu.ALU.u_wallace._0010_ ),
    .X(\u_cpu.ALU.u_wallace._0994_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5029_  (.A(\u_cpu.ALU.u_wallace._0512_ ),
    .B(\u_cpu.ALU.u_wallace._0250_ ),
    .C(\u_cpu.ALU.u_wallace._0523_ ),
    .D(\u_cpu.ALU.u_wallace._0545_ ),
    .X(\u_cpu.ALU.u_wallace._1005_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._5030_  (.A1(\u_cpu.ALU.u_wallace._0501_ ),
    .A2(\u_cpu.ALU.u_wallace._0983_ ),
    .A3(\u_cpu.ALU.u_wallace._0994_ ),
    .B1(\u_cpu.ALU.u_wallace._1005_ ),
    .X(\u_cpu.ALU.u_wallace._1016_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5031_  (.A(\u_cpu.ALU.SrcB[4] ),
    .X(\u_cpu.ALU.u_wallace._1026_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._5032_  (.A(\u_cpu.ALU.u_wallace._1026_ ),
    .Y(\u_cpu.ALU.u_wallace._1037_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5033_  (.A(\u_cpu.ALU.u_wallace._0032_ ),
    .B(\u_cpu.ALU.u_wallace._1037_ ),
    .Y(\u_cpu.ALU.u_wallace._1048_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5034_  (.A(\u_cpu.ALU.u_wallace._1016_ ),
    .B(\u_cpu.ALU.u_wallace._1048_ ),
    .Y(\u_cpu.ALU.u_wallace._1059_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5035_  (.A(\u_cpu.ALU.u_wallace._0446_ ),
    .X(\u_cpu.ALU.u_wallace._1070_ ));
 sky130_fd_sc_hd__a311o_2 \u_cpu.ALU.u_wallace._5036_  (.A1(\u_cpu.ALU.u_wallace._1070_ ),
    .A2(\u_cpu.ALU.u_wallace._0983_ ),
    .A3(\u_cpu.ALU.u_wallace._0501_ ),
    .B1(\u_cpu.ALU.u_wallace._1005_ ),
    .C1(\u_cpu.ALU.u_wallace._1048_ ),
    .X(\u_cpu.ALU.u_wallace._1081_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5037_  (.A(\u_cpu.ALU.u_wallace._0961_ ),
    .B(\u_cpu.ALU.u_wallace._0972_ ),
    .C(\u_cpu.ALU.u_wallace._1059_ ),
    .D(\u_cpu.ALU.u_wallace._1081_ ),
    .Y(\u_cpu.ALU.u_wallace._1092_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5038_  (.A1(\u_cpu.ALU.u_wallace._0961_ ),
    .A2(\u_cpu.ALU.u_wallace._0972_ ),
    .B1(\u_cpu.ALU.u_wallace._1059_ ),
    .B2(\u_cpu.ALU.u_wallace._1081_ ),
    .X(\u_cpu.ALU.u_wallace._1103_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5039_  (.A(\u_cpu.ALU.SrcA[5] ),
    .X(\u_cpu.ALU.u_wallace._1114_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5040_  (.A(\u_cpu.ALU.u_wallace._1114_ ),
    .X(\u_cpu.ALU.u_wallace._1125_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5041_  (.A(\u_cpu.ALU.u_wallace._1125_ ),
    .X(\u_cpu.ALU.u_wallace._1136_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5042_  (.A1(\u_cpu.ALU.u_wallace._0775_ ),
    .A2(\u_cpu.ALU.SrcA[4] ),
    .B1(\u_cpu.ALU.u_wallace._0764_ ),
    .B2(\u_cpu.ALU.u_wallace._0293_ ),
    .Y(\u_cpu.ALU.u_wallace._1147_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5043_  (.A(\u_cpu.ALU.u_wallace._0775_ ),
    .X(\u_cpu.ALU.u_wallace._1158_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5044_  (.A(\u_cpu.ALU.u_wallace._0534_ ),
    .X(\u_cpu.ALU.u_wallace._1169_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5045_  (.A(\u_cpu.ALU.SrcA[4] ),
    .X(\u_cpu.ALU.u_wallace._1180_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5046_  (.A(\u_cpu.ALU.u_wallace._0764_ ),
    .X(\u_cpu.ALU.u_wallace._1191_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5047_  (.A(\u_cpu.ALU.u_wallace._1158_ ),
    .B(\u_cpu.ALU.u_wallace._1169_ ),
    .C(\u_cpu.ALU.u_wallace._1180_ ),
    .D(\u_cpu.ALU.u_wallace._1191_ ),
    .Y(\u_cpu.ALU.u_wallace._1202_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._5048_  (.A_N(\u_cpu.ALU.u_wallace._1147_ ),
    .B(\u_cpu.ALU.u_wallace._1202_ ),
    .C(\u_cpu.ALU.u_wallace._0359_ ),
    .D(\u_cpu.ALU.u_wallace._0578_ ),
    .Y(\u_cpu.ALU.u_wallace._1213_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._5049_  (.A(\u_cpu.ALU.SrcB[3] ),
    .Y(\u_cpu.ALU.u_wallace._1224_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5050_  (.A(\u_cpu.ALU.u_wallace._0797_ ),
    .B(\u_cpu.ALU.u_wallace._0293_ ),
    .C(\u_cpu.ALU.u_wallace._0895_ ),
    .D(\u_cpu.ALU.u_wallace._0764_ ),
    .X(\u_cpu.ALU.u_wallace._1235_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5051_  (.A1(\u_cpu.ALU.u_wallace._0403_ ),
    .A2(\u_cpu.ALU.u_wallace._1224_ ),
    .B1(\u_cpu.ALU.u_wallace._1147_ ),
    .B2(\u_cpu.ALU.u_wallace._1235_ ),
    .Y(\u_cpu.ALU.u_wallace._1246_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5052_  (.A1(\u_cpu.ALU.u_wallace._0884_ ),
    .A2(\u_cpu.ALU.u_wallace._1136_ ),
    .B1(\u_cpu.ALU.u_wallace._1213_ ),
    .B2(\u_cpu.ALU.u_wallace._1246_ ),
    .X(\u_cpu.ALU.u_wallace._1256_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5053_  (.A(\u_cpu.ALU.SrcA[4] ),
    .X(\u_cpu.ALU.u_wallace._1267_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5054_  (.A(\u_cpu.ALU.SrcA[3] ),
    .X(\u_cpu.ALU.u_wallace._1278_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5055_  (.A(\u_cpu.ALU.u_wallace._0392_ ),
    .B(\u_cpu.ALU.u_wallace._0742_ ),
    .Y(\u_cpu.ALU.u_wallace._1289_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._5056_  (.A1(\u_cpu.ALU.u_wallace._0523_ ),
    .A2(\u_cpu.ALU.u_wallace._0545_ ),
    .A3(\u_cpu.ALU.u_wallace._1267_ ),
    .A4(\u_cpu.ALU.u_wallace._1278_ ),
    .B1(\u_cpu.ALU.u_wallace._1289_ ),
    .X(\u_cpu.ALU.u_wallace._1300_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5057_  (.A(\u_cpu.ALU.SrcA[5] ),
    .X(\u_cpu.ALU.u_wallace._1311_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5058_  (.A(\u_cpu.ALU.u_wallace._1311_ ),
    .X(\u_cpu.ALU.u_wallace._1322_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5059_  (.A(\u_cpu.ALU.u_wallace._1322_ ),
    .X(\u_cpu.ALU.u_wallace._1333_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._5060_  (.A1(\u_cpu.ALU.u_wallace._1147_ ),
    .A2(\u_cpu.ALU.u_wallace._1300_ ),
    .B1(\u_cpu.ALU.u_wallace._0884_ ),
    .C1(\u_cpu.ALU.u_wallace._1333_ ),
    .D1(\u_cpu.ALU.u_wallace._1246_ ),
    .Y(\u_cpu.ALU.u_wallace._1344_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._5061_  (.A_N(\u_cpu.ALU.u_wallace._0928_ ),
    .B(\u_cpu.ALU.u_wallace._1256_ ),
    .C(\u_cpu.ALU.u_wallace._1344_ ),
    .Y(\u_cpu.ALU.u_wallace._1355_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5062_  (.A1(\u_cpu.ALU.u_wallace._0884_ ),
    .A2(\u_cpu.ALU.u_wallace._1136_ ),
    .B1(\u_cpu.ALU.u_wallace._1213_ ),
    .B2(\u_cpu.ALU.u_wallace._1246_ ),
    .Y(\u_cpu.ALU.u_wallace._1366_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._5063_  (.A1(\u_cpu.ALU.u_wallace._1147_ ),
    .A2(\u_cpu.ALU.u_wallace._1300_ ),
    .B1(\u_cpu.ALU.u_wallace._0086_ ),
    .C1(\u_cpu.ALU.u_wallace._1136_ ),
    .D1(\u_cpu.ALU.u_wallace._1246_ ),
    .X(\u_cpu.ALU.u_wallace._1377_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5064_  (.A1(\u_cpu.ALU.u_wallace._1366_ ),
    .A2(\u_cpu.ALU.u_wallace._1377_ ),
    .B1(\u_cpu.ALU.u_wallace._0928_ ),
    .Y(\u_cpu.ALU.u_wallace._1388_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5065_  (.A(\u_cpu.ALU.u_wallace._0151_ ),
    .B(\u_cpu.ALU.u_wallace._0840_ ),
    .Y(\u_cpu.ALU.u_wallace._1399_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5066_  (.A(\u_cpu.ALU.SrcA[2] ),
    .X(\u_cpu.ALU.u_wallace._1410_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5067_  (.A(\u_cpu.ALU.u_wallace._0764_ ),
    .X(\u_cpu.ALU.u_wallace._1421_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5068_  (.A1(\u_cpu.ALU.u_wallace._1410_ ),
    .A2(\u_cpu.ALU.u_wallace._1169_ ),
    .B1(\u_cpu.ALU.u_wallace._1421_ ),
    .B2(\u_cpu.ALU.u_wallace._1158_ ),
    .Y(\u_cpu.ALU.u_wallace._1432_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5069_  (.A1(\u_cpu.ALU.u_wallace._1399_ ),
    .A2(\u_cpu.ALU.u_wallace._1432_ ),
    .B1(\u_cpu.ALU.u_wallace._0818_ ),
    .Y(\u_cpu.ALU.u_wallace._1443_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5070_  (.A(\u_cpu.ALU.u_wallace._0140_ ),
    .X(\u_cpu.ALU.u_wallace._1454_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5071_  (.A(\u_cpu.ALU.SrcB[4] ),
    .X(\u_cpu.ALU.u_wallace._1465_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5072_  (.A(\u_cpu.ALU.u_wallace._1465_ ),
    .X(\u_cpu.ALU.u_wallace._1476_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5073_  (.A(\u_cpu.ALU.SrcB[5] ),
    .X(\u_cpu.ALU.u_wallace._1486_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5074_  (.A(\u_cpu.ALU.u_wallace._1486_ ),
    .X(\u_cpu.ALU.u_wallace._1497_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5075_  (.A(\u_cpu.ALU.u_wallace._1497_ ),
    .X(\u_cpu.ALU.u_wallace._1508_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5076_  (.A(\u_cpu.ALU.u_wallace._0021_ ),
    .B(\u_cpu.ALU.u_wallace._1454_ ),
    .C(\u_cpu.ALU.u_wallace._1476_ ),
    .D(\u_cpu.ALU.u_wallace._1508_ ),
    .Y(\u_cpu.ALU.u_wallace._1519_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5077_  (.A(\u_cpu.ALU.u_wallace._1026_ ),
    .X(\u_cpu.ALU.u_wallace._1530_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5078_  (.A(\u_cpu.ALU.SrcB[5] ),
    .X(\u_cpu.ALU.u_wallace._1541_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5079_  (.A(\u_cpu.ALU.u_wallace._1541_ ),
    .X(\u_cpu.ALU.u_wallace._1552_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5080_  (.A1(\u_cpu.ALU.u_wallace._0731_ ),
    .A2(\u_cpu.ALU.u_wallace._1530_ ),
    .B1(\u_cpu.ALU.u_wallace._1552_ ),
    .B2(\u_cpu.ALU.u_wallace._0021_ ),
    .X(\u_cpu.ALU.u_wallace._1563_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5081_  (.A(\u_cpu.ALU.u_wallace._1443_ ),
    .B(\u_cpu.ALU.u_wallace._1519_ ),
    .C(\u_cpu.ALU.u_wallace._1563_ ),
    .X(\u_cpu.ALU.u_wallace._1574_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5082_  (.A(\u_cpu.ALU.u_wallace._1519_ ),
    .B(\u_cpu.ALU.u_wallace._1563_ ),
    .Y(\u_cpu.ALU.u_wallace._1585_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5083_  (.A1(\u_cpu.ALU.u_wallace._1399_ ),
    .A2(\u_cpu.ALU.u_wallace._1432_ ),
    .B1(\u_cpu.ALU.u_wallace._0818_ ),
    .C1(\u_cpu.ALU.u_wallace._1585_ ),
    .X(\u_cpu.ALU.u_wallace._1596_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5084_  (.A1_N(\u_cpu.ALU.u_wallace._1355_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1388_ ),
    .B1(\u_cpu.ALU.u_wallace._1574_ ),
    .B2(\u_cpu.ALU.u_wallace._1596_ ),
    .Y(\u_cpu.ALU.u_wallace._1607_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5085_  (.A(\u_cpu.ALU.u_wallace._1574_ ),
    .B(\u_cpu.ALU.u_wallace._1596_ ),
    .Y(\u_cpu.ALU.u_wallace._1618_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5086_  (.A(\u_cpu.ALU.u_wallace._1355_ ),
    .B(\u_cpu.ALU.u_wallace._1388_ ),
    .C(\u_cpu.ALU.u_wallace._1618_ ),
    .Y(\u_cpu.ALU.u_wallace._1629_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5087_  (.A(\u_cpu.ALU.u_wallace._1059_ ),
    .B(\u_cpu.ALU.u_wallace._1081_ ),
    .Y(\u_cpu.ALU.u_wallace._1640_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5088_  (.A1(\u_cpu.ALU.u_wallace._0928_ ),
    .A2(\u_cpu.ALU.u_wallace._0950_ ),
    .B1(\u_cpu.ALU.u_wallace._0643_ ),
    .Y(\u_cpu.ALU.u_wallace._1651_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5089_  (.A1(\u_cpu.ALU.u_wallace._1640_ ),
    .A2(\u_cpu.ALU.u_wallace._1651_ ),
    .B1(\u_cpu.ALU.u_wallace._0972_ ),
    .Y(\u_cpu.ALU.u_wallace._1662_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5090_  (.A1(\u_cpu.ALU.u_wallace._1607_ ),
    .A2(\u_cpu.ALU.u_wallace._1629_ ),
    .B1(\u_cpu.ALU.u_wallace._1662_ ),
    .X(\u_cpu.ALU.u_wallace._1673_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5091_  (.A(\u_cpu.ALU.u_wallace._1662_ ),
    .B(\u_cpu.ALU.u_wallace._1607_ ),
    .C(\u_cpu.ALU.u_wallace._1629_ ),
    .Y(\u_cpu.ALU.u_wallace._1684_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5092_  (.A1(\u_cpu.ALU.u_wallace._1016_ ),
    .A2(\u_cpu.ALU.u_wallace._1048_ ),
    .B1(\u_cpu.ALU.u_wallace._1673_ ),
    .B2(\u_cpu.ALU.u_wallace._1684_ ),
    .X(\u_cpu.ALU.u_wallace._1694_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5093_  (.A(\u_cpu.ALU.u_wallace._1016_ ),
    .B(\u_cpu.ALU.u_wallace._1684_ ),
    .C(\u_cpu.ALU.u_wallace._1673_ ),
    .D(\u_cpu.ALU.u_wallace._1048_ ),
    .Y(\u_cpu.ALU.u_wallace._1705_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5094_  (.A(\u_cpu.ALU.u_wallace._1092_ ),
    .B(\u_cpu.ALU.u_wallace._1103_ ),
    .C(\u_cpu.ALU.u_wallace._1694_ ),
    .D(\u_cpu.ALU.u_wallace._1705_ ),
    .Y(\u_cpu.ALU.u_wallace._1716_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5095_  (.A(\u_cpu.ALU.u_wallace._0687_ ),
    .B(\u_cpu.ALU.u_wallace._1103_ ),
    .C(\u_cpu.ALU.u_wallace._0665_ ),
    .D(\u_cpu.ALU.u_wallace._1092_ ),
    .X(\u_cpu.ALU.u_wallace._1727_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5096_  (.A(\u_cpu.ALU.u_wallace._1694_ ),
    .B(\u_cpu.ALU.u_wallace._1705_ ),
    .C(\u_cpu.ALU.u_wallace._1727_ ),
    .Y(\u_cpu.ALU.u_wallace._1738_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5097_  (.A(\u_cpu.ALU.u_wallace._0064_ ),
    .X(\u_cpu.ALU.u_wallace._1749_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5098_  (.A(\u_cpu.ALU.SrcB[6] ),
    .X(\u_cpu.ALU.u_wallace._1760_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5099_  (.A(\u_cpu.ALU.u_wallace._1760_ ),
    .X(\u_cpu.ALU.u_wallace._1771_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5100_  (.A(\u_cpu.ALU.SrcA[6] ),
    .X(\u_cpu.ALU.u_wallace._1782_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5101_  (.A(\u_cpu.ALU.u_wallace._1782_ ),
    .X(\u_cpu.ALU.u_wallace._1793_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5102_  (.A(\u_cpu.ALU.u_wallace._1749_ ),
    .B(\u_cpu.ALU.u_wallace._0010_ ),
    .C(\u_cpu.ALU.u_wallace._1771_ ),
    .D(\u_cpu.ALU.u_wallace._1793_ ),
    .X(\u_cpu.ALU.u_wallace._1804_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5103_  (.A(\u_cpu.ALU.SrcB[6] ),
    .X(\u_cpu.ALU.u_wallace._1815_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5104_  (.A(\u_cpu.ALU.u_wallace._1815_ ),
    .X(\u_cpu.ALU.u_wallace._1826_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5105_  (.A(\u_cpu.ALU.SrcA[6] ),
    .X(\u_cpu.ALU.u_wallace._1837_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5106_  (.A(\u_cpu.ALU.u_wallace._1837_ ),
    .X(\u_cpu.ALU.u_wallace._1848_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5107_  (.A(\u_cpu.ALU.u_wallace._0064_ ),
    .X(\u_cpu.ALU.u_wallace._1859_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5108_  (.A1(\u_cpu.ALU.u_wallace._0021_ ),
    .A2(\u_cpu.ALU.u_wallace._1826_ ),
    .B1(\u_cpu.ALU.u_wallace._1848_ ),
    .B2(\u_cpu.ALU.u_wallace._1859_ ),
    .Y(\u_cpu.ALU.u_wallace._1870_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5109_  (.A(\u_cpu.ALU.u_wallace._1804_ ),
    .B(\u_cpu.ALU.u_wallace._1870_ ),
    .Y(\u_cpu.ALU.u_wallace._1881_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5110_  (.A(\u_cpu.ALU.u_wallace._1224_ ),
    .X(\u_cpu.ALU.u_wallace._1892_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5111_  (.A(\u_cpu.ALU.u_wallace._0195_ ),
    .X(\u_cpu.ALU.u_wallace._1903_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5112_  (.A(\u_cpu.ALU.u_wallace._0282_ ),
    .X(\u_cpu.ALU.u_wallace._1914_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5113_  (.A1(\u_cpu.ALU.u_wallace._1903_ ),
    .A2(\u_cpu.ALU.u_wallace._1311_ ),
    .B1(\u_cpu.ALU.u_wallace._0895_ ),
    .B2(\u_cpu.ALU.u_wallace._1914_ ),
    .Y(\u_cpu.ALU.u_wallace._1924_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5114_  (.A(\u_cpu.ALU.u_wallace._0479_ ),
    .B(\u_cpu.ALU.u_wallace._0807_ ),
    .C(\u_cpu.ALU.u_wallace._1311_ ),
    .D(\u_cpu.ALU.u_wallace._0895_ ),
    .X(\u_cpu.ALU.u_wallace._1935_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5115_  (.A1(\u_cpu.ALU.u_wallace._1892_ ),
    .A2(\u_cpu.ALU.u_wallace._0610_ ),
    .B1(\u_cpu.ALU.u_wallace._1924_ ),
    .B2(\u_cpu.ALU.u_wallace._1935_ ),
    .Y(\u_cpu.ALU.u_wallace._1946_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5116_  (.A(\u_cpu.ALU.u_wallace._0195_ ),
    .X(\u_cpu.ALU.u_wallace._1957_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5117_  (.A(\u_cpu.ALU.u_wallace._0282_ ),
    .X(\u_cpu.ALU.u_wallace._1968_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5118_  (.A(\u_cpu.ALU.u_wallace._1114_ ),
    .X(\u_cpu.ALU.u_wallace._1979_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5119_  (.A(\u_cpu.ALU.u_wallace._1957_ ),
    .B(\u_cpu.ALU.u_wallace._1968_ ),
    .C(\u_cpu.ALU.u_wallace._1979_ ),
    .D(\u_cpu.ALU.u_wallace._1267_ ),
    .Y(\u_cpu.ALU.u_wallace._1990_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._5120_  (.A_N(\u_cpu.ALU.u_wallace._1924_ ),
    .B(\u_cpu.ALU.u_wallace._1990_ ),
    .C(\u_cpu.ALU.u_wallace._0468_ ),
    .D(\u_cpu.ALU.u_wallace._1421_ ),
    .Y(\u_cpu.ALU.u_wallace._2001_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5121_  (.A(\u_cpu.ALU.u_wallace._1881_ ),
    .B(\u_cpu.ALU.u_wallace._1946_ ),
    .C(\u_cpu.ALU.u_wallace._2001_ ),
    .X(\u_cpu.ALU.u_wallace._2012_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5122_  (.A1_N(\u_cpu.ALU.u_wallace._2001_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1946_ ),
    .B1(\u_cpu.ALU.u_wallace._1804_ ),
    .B2(\u_cpu.ALU.u_wallace._1870_ ),
    .Y(\u_cpu.ALU.u_wallace._2023_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5123_  (.A(\u_cpu.ALU.u_wallace._1377_ ),
    .B(\u_cpu.ALU.u_wallace._2023_ ),
    .Y(\u_cpu.ALU.u_wallace._2034_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5124_  (.A(\u_cpu.ALU.SrcB[4] ),
    .X(\u_cpu.ALU.u_wallace._2045_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5125_  (.A(\u_cpu.ALU.u_wallace._1486_ ),
    .X(\u_cpu.ALU.u_wallace._2056_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5126_  (.A(\u_cpu.ALU.u_wallace._0512_ ),
    .B(\u_cpu.ALU.u_wallace._0250_ ),
    .C(\u_cpu.ALU.u_wallace._2045_ ),
    .D(\u_cpu.ALU.u_wallace._2056_ ),
    .Y(\u_cpu.ALU.u_wallace._2067_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5127_  (.A(\u_cpu.ALU.u_wallace._1486_ ),
    .X(\u_cpu.ALU.u_wallace._2078_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5128_  (.A1(\u_cpu.ALU.u_wallace._0348_ ),
    .A2(\u_cpu.ALU.u_wallace._1465_ ),
    .B1(\u_cpu.ALU.u_wallace._2078_ ),
    .B2(\u_cpu.ALU.u_wallace._0250_ ),
    .X(\u_cpu.ALU.u_wallace._2089_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5129_  (.A(\u_cpu.ALU.u_wallace._2067_ ),
    .B(\u_cpu.ALU.u_wallace._2089_ ),
    .Y(\u_cpu.ALU.u_wallace._2100_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5130_  (.A1(\u_cpu.ALU.u_wallace._1289_ ),
    .A2(\u_cpu.ALU.u_wallace._1147_ ),
    .B1(\u_cpu.ALU.u_wallace._1202_ ),
    .C1(\u_cpu.ALU.u_wallace._2100_ ),
    .Y(\u_cpu.ALU.u_wallace._2111_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5131_  (.A1(\u_cpu.ALU.u_wallace._1289_ ),
    .A2(\u_cpu.ALU.u_wallace._1147_ ),
    .B1(\u_cpu.ALU.u_wallace._1202_ ),
    .Y(\u_cpu.ALU.u_wallace._2122_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5132_  (.A(\u_cpu.ALU.u_wallace._2122_ ),
    .B(\u_cpu.ALU.u_wallace._2067_ ),
    .C(\u_cpu.ALU.u_wallace._2089_ ),
    .Y(\u_cpu.ALU.u_wallace._2133_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5133_  (.A(\u_cpu.ALU.SrcB[4] ),
    .X(\u_cpu.ALU.u_wallace._2144_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5134_  (.A(\u_cpu.ALU.u_wallace._2144_ ),
    .X(\u_cpu.ALU.u_wallace._2155_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5135_  (.A(\u_cpu.ALU.u_wallace._2155_ ),
    .X(\u_cpu.ALU.u_wallace._2166_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5136_  (.A(\u_cpu.ALU.u_wallace._0162_ ),
    .B(\u_cpu.ALU.u_wallace._2166_ ),
    .Y(\u_cpu.ALU.u_wallace._2176_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5137_  (.A(\u_cpu.ALU.u_wallace._1541_ ),
    .X(\u_cpu.ALU.u_wallace._2187_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5138_  (.A(\u_cpu.ALU.u_wallace._2187_ ),
    .X(\u_cpu.ALU.u_wallace._2198_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5139_  (.A(\u_cpu.ALU.u_wallace._0108_ ),
    .B(\u_cpu.ALU.u_wallace._2198_ ),
    .Y(\u_cpu.ALU.u_wallace._2209_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5140_  (.A1_N(\u_cpu.ALU.u_wallace._2111_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2133_ ),
    .B1(\u_cpu.ALU.u_wallace._2176_ ),
    .B2(\u_cpu.ALU.u_wallace._2209_ ),
    .Y(\u_cpu.ALU.u_wallace._2220_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5141_  (.A(\u_cpu.ALU.u_wallace._0446_ ),
    .B(\u_cpu.ALU.u_wallace._0261_ ),
    .C(\u_cpu.ALU.u_wallace._1476_ ),
    .D(\u_cpu.ALU.u_wallace._1508_ ),
    .X(\u_cpu.ALU.u_wallace._2231_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5142_  (.A(\u_cpu.ALU.u_wallace._2133_ ),
    .B(\u_cpu.ALU.u_wallace._2231_ ),
    .C(\u_cpu.ALU.u_wallace._2111_ ),
    .Y(\u_cpu.ALU.u_wallace._2242_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5143_  (.A1(\u_cpu.ALU.u_wallace._2012_ ),
    .A2(\u_cpu.ALU.u_wallace._2034_ ),
    .B1(\u_cpu.ALU.u_wallace._2220_ ),
    .C1(\u_cpu.ALU.u_wallace._2242_ ),
    .Y(\u_cpu.ALU.u_wallace._2253_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5144_  (.A(\u_cpu.ALU.u_wallace._1881_ ),
    .B(\u_cpu.ALU.u_wallace._1946_ ),
    .C(\u_cpu.ALU.u_wallace._2001_ ),
    .Y(\u_cpu.ALU.u_wallace._2264_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5145_  (.A1(\u_cpu.ALU.u_wallace._2023_ ),
    .A2(\u_cpu.ALU.u_wallace._2264_ ),
    .B1(\u_cpu.ALU.u_wallace._1377_ ),
    .Y(\u_cpu.ALU.u_wallace._2275_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._5146_  (.A(\u_cpu.ALU.u_wallace._0928_ ),
    .B(\u_cpu.ALU.u_wallace._1366_ ),
    .C(\u_cpu.ALU.u_wallace._1377_ ),
    .Y(\u_cpu.ALU.u_wallace._2286_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5147_  (.A1(\u_cpu.ALU.u_wallace._1388_ ),
    .A2(\u_cpu.ALU.u_wallace._1618_ ),
    .B1(\u_cpu.ALU.u_wallace._2286_ ),
    .X(\u_cpu.ALU.u_wallace._2297_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5148_  (.A(\u_cpu.ALU.u_wallace._1377_ ),
    .B(\u_cpu.ALU.u_wallace._2023_ ),
    .C(\u_cpu.ALU.u_wallace._2264_ ),
    .X(\u_cpu.ALU.u_wallace._2308_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5149_  (.A(\u_cpu.ALU.u_wallace._2220_ ),
    .B(\u_cpu.ALU.u_wallace._2242_ ),
    .Y(\u_cpu.ALU.u_wallace._2319_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5150_  (.A1(\u_cpu.ALU.u_wallace._2308_ ),
    .A2(\u_cpu.ALU.u_wallace._2275_ ),
    .B1(\u_cpu.ALU.u_wallace._2319_ ),
    .Y(\u_cpu.ALU.u_wallace._2330_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5151_  (.A1(\u_cpu.ALU.u_wallace._2253_ ),
    .A2(\u_cpu.ALU.u_wallace._2275_ ),
    .B1(\u_cpu.ALU.u_wallace._2297_ ),
    .C1(\u_cpu.ALU.u_wallace._2330_ ),
    .Y(\u_cpu.ALU.u_wallace._2341_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5152_  (.A1(\u_cpu.ALU.u_wallace._2012_ ),
    .A2(\u_cpu.ALU.u_wallace._2034_ ),
    .B1(\u_cpu.ALU.u_wallace._2275_ ),
    .B2(\u_cpu.ALU.u_wallace._2319_ ),
    .Y(\u_cpu.ALU.u_wallace._2352_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5153_  (.A1(\u_cpu.ALU.u_wallace._1388_ ),
    .A2(\u_cpu.ALU.u_wallace._1618_ ),
    .B1(\u_cpu.ALU.u_wallace._2286_ ),
    .Y(\u_cpu.ALU.u_wallace._2363_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5154_  (.A1(\u_cpu.ALU.u_wallace._2308_ ),
    .A2(\u_cpu.ALU.u_wallace._2275_ ),
    .B1(\u_cpu.ALU.u_wallace._2220_ ),
    .C1(\u_cpu.ALU.u_wallace._2242_ ),
    .Y(\u_cpu.ALU.u_wallace._2374_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5155_  (.A1(\u_cpu.ALU.u_wallace._2275_ ),
    .A2(\u_cpu.ALU.u_wallace._2352_ ),
    .B1(\u_cpu.ALU.u_wallace._2363_ ),
    .C1(\u_cpu.ALU.u_wallace._2374_ ),
    .Y(\u_cpu.ALU.u_wallace._2385_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5156_  (.A(\u_cpu.ALU.u_wallace._2341_ ),
    .B(\u_cpu.ALU.u_wallace._2385_ ),
    .C(\u_cpu.ALU.u_wallace._1574_ ),
    .Y(\u_cpu.ALU.u_wallace._2396_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._5157_  (.A(\u_cpu.ALU.u_wallace._1443_ ),
    .Y(\u_cpu.ALU.u_wallace._2407_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5158_  (.A1_N(\u_cpu.ALU.u_wallace._2341_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2385_ ),
    .B1(\u_cpu.ALU.u_wallace._2407_ ),
    .B2(\u_cpu.ALU.u_wallace._1585_ ),
    .Y(\u_cpu.ALU.u_wallace._2418_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5159_  (.A1(\u_cpu.ALU.u_wallace._1607_ ),
    .A2(\u_cpu.ALU.u_wallace._1629_ ),
    .B1(\u_cpu.ALU.u_wallace._1662_ ),
    .Y(\u_cpu.ALU.u_wallace._2429_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5160_  (.A1(\u_cpu.ALU.u_wallace._1059_ ),
    .A2(\u_cpu.ALU.u_wallace._2429_ ),
    .B1(\u_cpu.ALU.u_wallace._1684_ ),
    .Y(\u_cpu.ALU.u_wallace._2440_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5161_  (.A1(\u_cpu.ALU.u_wallace._2396_ ),
    .A2(\u_cpu.ALU.u_wallace._2418_ ),
    .B1(\u_cpu.ALU.u_wallace._2440_ ),
    .Y(\u_cpu.ALU.u_wallace._2451_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5162_  (.A(\u_cpu.ALU.u_wallace._1738_ ),
    .B(\u_cpu.ALU.u_wallace._2451_ ),
    .Y(\u_cpu.ALU.u_wallace._2462_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5163_  (.A(\u_cpu.ALU.u_wallace._2440_ ),
    .B(\u_cpu.ALU.u_wallace._2396_ ),
    .C(\u_cpu.ALU.u_wallace._2418_ ),
    .X(\u_cpu.ALU.u_wallace._2472_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5164_  (.A1(\u_cpu.ALU.u_wallace._2451_ ),
    .A2(\u_cpu.ALU.u_wallace._2472_ ),
    .B1(\u_cpu.ALU.u_wallace._1738_ ),
    .Y(\u_cpu.ALU.u_wallace._2483_ ));
 sky130_fd_sc_hd__nor4b_2 \u_cpu.ALU.u_wallace._5165_  (.A(\u_cpu.ALU.u_wallace._0720_ ),
    .B(\u_cpu.ALU.u_wallace._1716_ ),
    .C(\u_cpu.ALU.u_wallace._2462_ ),
    .D_N(\u_cpu.ALU.u_wallace._2483_ ),
    .Y(\u_cpu.ALU.u_wallace._2494_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5166_  (.A(\u_cpu.ALU.u_wallace._2341_ ),
    .B(\u_cpu.ALU.u_wallace._2396_ ),
    .Y(\u_cpu.ALU.u_wallace._2505_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5167_  (.A(\u_cpu.ALU.u_wallace._0468_ ),
    .B(\u_cpu.ALU.u_wallace._1421_ ),
    .Y(\u_cpu.ALU.u_wallace._2516_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5168_  (.A(\u_cpu.ALU.u_wallace._2516_ ),
    .B(\u_cpu.ALU.u_wallace._1924_ ),
    .Y(\u_cpu.ALU.u_wallace._2527_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5169_  (.A(\u_cpu.ALU.SrcB[5] ),
    .X(\u_cpu.ALU.u_wallace._2538_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5170_  (.A(\u_cpu.ALU.SrcA[3] ),
    .X(\u_cpu.ALU.u_wallace._2549_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5171_  (.A1(\u_cpu.ALU.u_wallace._0392_ ),
    .A2(\u_cpu.ALU.u_wallace._2538_ ),
    .B1(\u_cpu.ALU.u_wallace._2549_ ),
    .B2(\u_cpu.ALU.u_wallace._1465_ ),
    .X(\u_cpu.ALU.u_wallace._2560_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5172_  (.A(\u_cpu.ALU.SrcB[4] ),
    .X(\u_cpu.ALU.u_wallace._2571_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5173_  (.A(\u_cpu.ALU.u_wallace._1486_ ),
    .X(\u_cpu.ALU.u_wallace._2582_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5174_  (.A(\u_cpu.ALU.u_wallace._0348_ ),
    .B(\u_cpu.ALU.u_wallace._2571_ ),
    .C(\u_cpu.ALU.u_wallace._2582_ ),
    .D(\u_cpu.ALU.u_wallace._1278_ ),
    .Y(\u_cpu.ALU.u_wallace._2593_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5175_  (.A(\u_cpu.ALU.SrcB[7] ),
    .X(\u_cpu.ALU.u_wallace._2604_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5176_  (.A(\u_cpu.ALU.u_wallace._2560_ ),
    .B(\u_cpu.ALU.u_wallace._2593_ ),
    .C(\u_cpu.ALU.u_wallace._0446_ ),
    .D(\u_cpu.ALU.u_wallace._2604_ ),
    .Y(\u_cpu.ALU.u_wallace._2615_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5177_  (.A(\u_cpu.ALU.SrcB[7] ),
    .X(\u_cpu.ALU.u_wallace._2626_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5178_  (.A1(\u_cpu.ALU.u_wallace._0021_ ),
    .A2(\u_cpu.ALU.u_wallace._2626_ ),
    .B1(\u_cpu.ALU.u_wallace._2560_ ),
    .B2(\u_cpu.ALU.u_wallace._2593_ ),
    .X(\u_cpu.ALU.u_wallace._2637_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5179_  (.A1(\u_cpu.ALU.u_wallace._1935_ ),
    .A2(\u_cpu.ALU.u_wallace._2527_ ),
    .B1(\u_cpu.ALU.u_wallace._2615_ ),
    .C1(\u_cpu.ALU.u_wallace._2637_ ),
    .X(\u_cpu.ALU.u_wallace._2648_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5180_  (.A1(\u_cpu.ALU.u_wallace._2516_ ),
    .A2(\u_cpu.ALU.u_wallace._1924_ ),
    .B1(\u_cpu.ALU.u_wallace._1990_ ),
    .Y(\u_cpu.ALU.u_wallace._2659_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5181_  (.A1(\u_cpu.ALU.u_wallace._2615_ ),
    .A2(\u_cpu.ALU.u_wallace._2637_ ),
    .B1(\u_cpu.ALU.u_wallace._2659_ ),
    .Y(\u_cpu.ALU.u_wallace._2670_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5182_  (.A1(\u_cpu.ALU.u_wallace._2648_ ),
    .A2(\u_cpu.ALU.u_wallace._2670_ ),
    .B1(\u_cpu.ALU.u_wallace._2067_ ),
    .Y(\u_cpu.ALU.u_wallace._2681_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5183_  (.A(\u_cpu.ALU.u_wallace._0370_ ),
    .B(\u_cpu.ALU.u_wallace._0272_ ),
    .C(\u_cpu.ALU.u_wallace._2166_ ),
    .D(\u_cpu.ALU.u_wallace._2198_ ),
    .X(\u_cpu.ALU.u_wallace._2692_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5184_  (.A1(\u_cpu.ALU.u_wallace._1935_ ),
    .A2(\u_cpu.ALU.u_wallace._2527_ ),
    .B1(\u_cpu.ALU.u_wallace._2615_ ),
    .C1(\u_cpu.ALU.u_wallace._2637_ ),
    .Y(\u_cpu.ALU.u_wallace._2703_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._5185_  (.A_N(\u_cpu.ALU.u_wallace._2670_ ),
    .B(\u_cpu.ALU.u_wallace._2692_ ),
    .C(\u_cpu.ALU.u_wallace._2703_ ),
    .Y(\u_cpu.ALU.u_wallace._2714_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5186_  (.A(\u_cpu.ALU.SrcA[7] ),
    .X(\u_cpu.ALU.u_wallace._2725_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5187_  (.A1(\u_cpu.ALU.u_wallace._1859_ ),
    .A2(\u_cpu.ALU.u_wallace._2725_ ),
    .B1(\u_cpu.ALU.u_wallace._0731_ ),
    .B2(\u_cpu.ALU.u_wallace._1826_ ),
    .X(\u_cpu.ALU.u_wallace._2736_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5188_  (.A(\u_cpu.ALU.u_wallace._0064_ ),
    .X(\u_cpu.ALU.u_wallace._2747_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5189_  (.A(\u_cpu.ALU.u_wallace._2747_ ),
    .X(\u_cpu.ALU.u_wallace._2757_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5190_  (.A(\u_cpu.ALU.SrcB[6] ),
    .X(\u_cpu.ALU.u_wallace._2768_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5191_  (.A(\u_cpu.ALU.u_wallace._2768_ ),
    .X(\u_cpu.ALU.u_wallace._2779_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5192_  (.A(\u_cpu.ALU.SrcA[7] ),
    .X(\u_cpu.ALU.u_wallace._2790_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5193_  (.A(\u_cpu.ALU.u_wallace._2790_ ),
    .X(\u_cpu.ALU.u_wallace._2801_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5194_  (.A(\u_cpu.ALU.u_wallace._2757_ ),
    .B(\u_cpu.ALU.u_wallace._2779_ ),
    .C(\u_cpu.ALU.u_wallace._2801_ ),
    .D(\u_cpu.ALU.u_wallace._0151_ ),
    .Y(\u_cpu.ALU.u_wallace._2812_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5195_  (.A(\u_cpu.ALU.u_wallace._1804_ ),
    .B(\u_cpu.ALU.u_wallace._2736_ ),
    .C(\u_cpu.ALU.u_wallace._2812_ ),
    .Y(\u_cpu.ALU.u_wallace._2823_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5196_  (.A(\u_cpu.ALU.u_wallace._1782_ ),
    .X(\u_cpu.ALU.u_wallace._2834_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5197_  (.A(\u_cpu.ALU.u_wallace._2747_ ),
    .B(\u_cpu.ALU.u_wallace._2834_ ),
    .Y(\u_cpu.ALU.u_wallace._2845_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5198_  (.A(\u_cpu.ALU.u_wallace._1760_ ),
    .X(\u_cpu.ALU.u_wallace._2856_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5199_  (.A(\u_cpu.ALU.u_wallace._0010_ ),
    .B(\u_cpu.ALU.u_wallace._2856_ ),
    .Y(\u_cpu.ALU.u_wallace._2867_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5200_  (.A(\u_cpu.ALU.SrcA[7] ),
    .X(\u_cpu.ALU.u_wallace._2878_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5201_  (.A1(\u_cpu.ALU.u_wallace._0862_ ),
    .A2(\u_cpu.ALU.u_wallace._2878_ ),
    .B1(\u_cpu.ALU.u_wallace._0140_ ),
    .B2(\u_cpu.ALU.u_wallace._2768_ ),
    .Y(\u_cpu.ALU.u_wallace._2889_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5202_  (.A(\u_cpu.ALU.u_wallace._0064_ ),
    .B(\u_cpu.ALU.u_wallace._1760_ ),
    .C(\u_cpu.ALU.SrcA[7] ),
    .D(\u_cpu.ALU.SrcA[1] ),
    .X(\u_cpu.ALU.u_wallace._2900_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5203_  (.A1(\u_cpu.ALU.u_wallace._2845_ ),
    .A2(\u_cpu.ALU.u_wallace._2867_ ),
    .B1(\u_cpu.ALU.u_wallace._2889_ ),
    .B2(\u_cpu.ALU.u_wallace._2900_ ),
    .Y(\u_cpu.ALU.u_wallace._2911_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5204_  (.A(\u_cpu.ALU.SrcA[4] ),
    .X(\u_cpu.ALU.u_wallace._2922_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5205_  (.A(\u_cpu.ALU.u_wallace._2922_ ),
    .X(\u_cpu.ALU.u_wallace._2933_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5206_  (.A1(\u_cpu.ALU.u_wallace._0479_ ),
    .A2(\u_cpu.ALU.u_wallace._1837_ ),
    .B1(\u_cpu.ALU.u_wallace._1311_ ),
    .B2(\u_cpu.ALU.u_wallace._0490_ ),
    .X(\u_cpu.ALU.u_wallace._2944_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5207_  (.A(\u_cpu.ALU.u_wallace._1114_ ),
    .X(\u_cpu.ALU.u_wallace._2955_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5208_  (.A(\u_cpu.ALU.u_wallace._0206_ ),
    .B(\u_cpu.ALU.u_wallace._0490_ ),
    .C(\u_cpu.ALU.u_wallace._2834_ ),
    .D(\u_cpu.ALU.u_wallace._2955_ ),
    .Y(\u_cpu.ALU.u_wallace._2966_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5209_  (.A1(\u_cpu.ALU.u_wallace._0983_ ),
    .A2(\u_cpu.ALU.u_wallace._2933_ ),
    .B1(\u_cpu.ALU.u_wallace._2944_ ),
    .B2(\u_cpu.ALU.u_wallace._2966_ ),
    .Y(\u_cpu.ALU.u_wallace._2977_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5210_  (.A(\u_cpu.ALU.u_wallace._2944_ ),
    .B(\u_cpu.ALU.u_wallace._2966_ ),
    .C(\u_cpu.ALU.u_wallace._0840_ ),
    .D(\u_cpu.ALU.u_wallace._0906_ ),
    .X(\u_cpu.ALU.u_wallace._2988_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5211_  (.A1_N(\u_cpu.ALU.u_wallace._2823_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2911_ ),
    .B1(\u_cpu.ALU.u_wallace._2977_ ),
    .B2(\u_cpu.ALU.u_wallace._2988_ ),
    .Y(\u_cpu.ALU.u_wallace._2999_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5212_  (.A1(\u_cpu.ALU.u_wallace._0775_ ),
    .A2(\u_cpu.ALU.u_wallace._1782_ ),
    .B1(\u_cpu.ALU.u_wallace._1114_ ),
    .B2(\u_cpu.ALU.u_wallace._0534_ ),
    .Y(\u_cpu.ALU.u_wallace._3010_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5213_  (.A(\u_cpu.ALU.u_wallace._0195_ ),
    .B(\u_cpu.ALU.u_wallace._0282_ ),
    .C(\u_cpu.ALU.u_wallace._1782_ ),
    .D(\u_cpu.ALU.u_wallace._1114_ ),
    .X(\u_cpu.ALU.u_wallace._3021_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5214_  (.A1(\u_cpu.ALU.u_wallace._1224_ ),
    .A2(\u_cpu.ALU.u_wallace._0939_ ),
    .B1(\u_cpu.ALU.u_wallace._3010_ ),
    .B2(\u_cpu.ALU.u_wallace._3021_ ),
    .Y(\u_cpu.ALU.u_wallace._3032_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5215_  (.A(\u_cpu.ALU.u_wallace._2944_ ),
    .B(\u_cpu.ALU.u_wallace._2966_ ),
    .C(\u_cpu.ALU.u_wallace._0983_ ),
    .D(\u_cpu.ALU.u_wallace._0917_ ),
    .Y(\u_cpu.ALU.u_wallace._3042_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5216_  (.A(\u_cpu.ALU.u_wallace._2823_ ),
    .B(\u_cpu.ALU.u_wallace._2911_ ),
    .C(\u_cpu.ALU.u_wallace._3032_ ),
    .D(\u_cpu.ALU.u_wallace._3042_ ),
    .Y(\u_cpu.ALU.u_wallace._3053_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5217_  (.A1(\u_cpu.ALU.u_wallace._2999_ ),
    .A2(\u_cpu.ALU.u_wallace._3053_ ),
    .B1(\u_cpu.ALU.u_wallace._2012_ ),
    .Y(\u_cpu.ALU.u_wallace._3064_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5218_  (.A(\u_cpu.ALU.u_wallace._2012_ ),
    .B(\u_cpu.ALU.u_wallace._2999_ ),
    .C(\u_cpu.ALU.u_wallace._3053_ ),
    .X(\u_cpu.ALU.u_wallace._3075_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5219_  (.A1_N(\u_cpu.ALU.u_wallace._2681_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2714_ ),
    .B1(\u_cpu.ALU.u_wallace._3064_ ),
    .B2(\u_cpu.ALU.u_wallace._3075_ ),
    .Y(\u_cpu.ALU.u_wallace._3086_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5220_  (.A1(\u_cpu.ALU.u_wallace._2999_ ),
    .A2(\u_cpu.ALU.u_wallace._3053_ ),
    .B1(\u_cpu.ALU.u_wallace._2012_ ),
    .X(\u_cpu.ALU.u_wallace._3097_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5221_  (.A(\u_cpu.ALU.u_wallace._1804_ ),
    .B(\u_cpu.ALU.u_wallace._2736_ ),
    .C(\u_cpu.ALU.u_wallace._2812_ ),
    .X(\u_cpu.ALU.u_wallace._3108_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5222_  (.A(\u_cpu.ALU.u_wallace._0742_ ),
    .B(\u_cpu.ALU.u_wallace._0895_ ),
    .Y(\u_cpu.ALU.u_wallace._3119_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._5223_  (.A1(\u_cpu.ALU.u_wallace._1957_ ),
    .A2(\u_cpu.ALU.u_wallace._1968_ ),
    .A3(\u_cpu.ALU.u_wallace._1793_ ),
    .A4(\u_cpu.ALU.u_wallace._1979_ ),
    .B1(\u_cpu.ALU.u_wallace._3119_ ),
    .X(\u_cpu.ALU.u_wallace._3130_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5224_  (.A1(\u_cpu.ALU.u_wallace._3010_ ),
    .A2(\u_cpu.ALU.u_wallace._3130_ ),
    .B1(\u_cpu.ALU.u_wallace._3032_ ),
    .C1(\u_cpu.ALU.u_wallace._2911_ ),
    .Y(\u_cpu.ALU.u_wallace._3141_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5225_  (.A1(\u_cpu.ALU.u_wallace._3108_ ),
    .A2(\u_cpu.ALU.u_wallace._3141_ ),
    .B1(\u_cpu.ALU.u_wallace._2999_ ),
    .C1(\u_cpu.ALU.u_wallace._2012_ ),
    .Y(\u_cpu.ALU.u_wallace._3152_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5226_  (.A(\u_cpu.ALU.u_wallace._2681_ ),
    .B(\u_cpu.ALU.u_wallace._2714_ ),
    .C(\u_cpu.ALU.u_wallace._3097_ ),
    .D(\u_cpu.ALU.u_wallace._3152_ ),
    .Y(\u_cpu.ALU.u_wallace._3163_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5227_  (.A1(\u_cpu.ALU.u_wallace._3086_ ),
    .A2(\u_cpu.ALU.u_wallace._3163_ ),
    .B1(\u_cpu.ALU.u_wallace._2352_ ),
    .Y(\u_cpu.ALU.u_wallace._3174_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5228_  (.A(\u_cpu.ALU.u_wallace._2681_ ),
    .B(\u_cpu.ALU.u_wallace._2714_ ),
    .C(\u_cpu.ALU.u_wallace._3152_ ),
    .Y(\u_cpu.ALU.u_wallace._3185_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5229_  (.A1(\u_cpu.ALU.u_wallace._3064_ ),
    .A2(\u_cpu.ALU.u_wallace._3185_ ),
    .B1(\u_cpu.ALU.u_wallace._3086_ ),
    .C1(\u_cpu.ALU.u_wallace._2352_ ),
    .Y(\u_cpu.ALU.u_wallace._3196_ ));
 sky130_fd_sc_hd__a21bo_2 \u_cpu.ALU.u_wallace._5230_  (.A1(\u_cpu.ALU.u_wallace._2231_ ),
    .A2(\u_cpu.ALU.u_wallace._2111_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2133_ ),
    .X(\u_cpu.ALU.u_wallace._3207_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._5231_  (.A_N(\u_cpu.ALU.u_wallace._3174_ ),
    .B(\u_cpu.ALU.u_wallace._3196_ ),
    .C(\u_cpu.ALU.u_wallace._3207_ ),
    .Y(\u_cpu.ALU.u_wallace._3218_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5232_  (.A1(\u_cpu.ALU.u_wallace._3064_ ),
    .A2(\u_cpu.ALU.u_wallace._3185_ ),
    .B1(\u_cpu.ALU.u_wallace._3086_ ),
    .C1(\u_cpu.ALU.u_wallace._2352_ ),
    .X(\u_cpu.ALU.u_wallace._3229_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._5233_  (.A1(\u_cpu.ALU.u_wallace._3174_ ),
    .A2(\u_cpu.ALU.u_wallace._3229_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3207_ ),
    .Y(\u_cpu.ALU.u_wallace._3240_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5234_  (.A(\u_cpu.ALU.u_wallace._2505_ ),
    .B(\u_cpu.ALU.u_wallace._3218_ ),
    .C(\u_cpu.ALU.u_wallace._3240_ ),
    .X(\u_cpu.ALU.u_wallace._3251_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5235_  (.A(\u_cpu.ALU.u_wallace._2440_ ),
    .B(\u_cpu.ALU.u_wallace._2396_ ),
    .C(\u_cpu.ALU.u_wallace._2418_ ),
    .Y(\u_cpu.ALU.u_wallace._3262_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5236_  (.A1(\u_cpu.ALU.u_wallace._3218_ ),
    .A2(\u_cpu.ALU.u_wallace._3240_ ),
    .B1(\u_cpu.ALU.u_wallace._2505_ ),
    .X(\u_cpu.ALU.u_wallace._3273_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5237_  (.A1(\u_cpu.ALU.u_wallace._1738_ ),
    .A2(\u_cpu.ALU.u_wallace._2451_ ),
    .B1(\u_cpu.ALU.u_wallace._3262_ ),
    .C1(\u_cpu.ALU.u_wallace._3273_ ),
    .Y(\u_cpu.ALU.u_wallace._3284_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5238_  (.A1(\u_cpu.ALU.u_wallace._3218_ ),
    .A2(\u_cpu.ALU.u_wallace._3240_ ),
    .B1(\u_cpu.ALU.u_wallace._2505_ ),
    .Y(\u_cpu.ALU.u_wallace._3295_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5239_  (.A1(\u_cpu.ALU.u_wallace._2472_ ),
    .A2(\u_cpu.ALU.u_wallace._2462_ ),
    .B1(\u_cpu.ALU.u_wallace._3251_ ),
    .B2(\u_cpu.ALU.u_wallace._3295_ ),
    .Y(\u_cpu.ALU.u_wallace._3306_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5240_  (.A1(\u_cpu.ALU.u_wallace._3251_ ),
    .A2(\u_cpu.ALU.u_wallace._3284_ ),
    .B1(\u_cpu.ALU.u_wallace._3306_ ),
    .Y(\u_cpu.ALU.u_wallace._3317_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5241_  (.A(\u_cpu.ALU.u_wallace._2505_ ),
    .B(\u_cpu.ALU.u_wallace._3218_ ),
    .C(\u_cpu.ALU.u_wallace._3240_ ),
    .Y(\u_cpu.ALU.u_wallace._3328_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._5242_  (.A1(\u_cpu.ALU.u_wallace._2681_ ),
    .A2(\u_cpu.ALU.u_wallace._2714_ ),
    .A3(\u_cpu.ALU.u_wallace._3097_ ),
    .B1(\u_cpu.ALU.u_wallace._3075_ ),
    .X(\u_cpu.ALU.u_wallace._3338_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5243_  (.A1(\u_cpu.ALU.u_wallace._2922_ ),
    .A2(\u_cpu.ALU.u_wallace._1465_ ),
    .B1(\u_cpu.ALU.u_wallace._2582_ ),
    .B2(\u_cpu.ALU.u_wallace._0600_ ),
    .Y(\u_cpu.ALU.u_wallace._3349_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5244_  (.A(\u_cpu.ALU.u_wallace._0895_ ),
    .B(\u_cpu.ALU.u_wallace._1026_ ),
    .C(\u_cpu.ALU.u_wallace._1541_ ),
    .D(\u_cpu.ALU.u_wallace._0764_ ),
    .X(\u_cpu.ALU.u_wallace._3360_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._5245_  (.A(\u_cpu.ALU.u_wallace._0140_ ),
    .B(\u_cpu.ALU.SrcB[7] ),
    .X(\u_cpu.ALU.u_wallace._3371_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._5246_  (.A1(\u_cpu.ALU.u_wallace._3349_ ),
    .A2(\u_cpu.ALU.u_wallace._3360_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3371_ ),
    .Y(\u_cpu.ALU.u_wallace._3382_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5247_  (.A(\u_cpu.ALU.u_wallace._2922_ ),
    .B(\u_cpu.ALU.u_wallace._2078_ ),
    .C(\u_cpu.ALU.u_wallace._0600_ ),
    .Y(\u_cpu.ALU.u_wallace._3393_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5248_  (.A(\u_cpu.ALU.SrcB[7] ),
    .X(\u_cpu.ALU.u_wallace._3404_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5249_  (.A1(\u_cpu.ALU.u_wallace._0895_ ),
    .A2(\u_cpu.ALU.u_wallace._2144_ ),
    .B1(\u_cpu.ALU.u_wallace._2538_ ),
    .B2(\u_cpu.ALU.u_wallace._2549_ ),
    .X(\u_cpu.ALU.u_wallace._3415_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._5250_  (.A1(\u_cpu.ALU.u_wallace._1037_ ),
    .A2(\u_cpu.ALU.u_wallace._3393_ ),
    .B1(\u_cpu.ALU.u_wallace._3404_ ),
    .C1(\u_cpu.ALU.u_wallace._1454_ ),
    .D1(\u_cpu.ALU.u_wallace._3415_ ),
    .Y(\u_cpu.ALU.u_wallace._3426_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5251_  (.A1(\u_cpu.ALU.u_wallace._3119_ ),
    .A2(\u_cpu.ALU.u_wallace._3010_ ),
    .B1(\u_cpu.ALU.u_wallace._2966_ ),
    .Y(\u_cpu.ALU.u_wallace._3437_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5252_  (.A1(\u_cpu.ALU.u_wallace._3382_ ),
    .A2(\u_cpu.ALU.u_wallace._3426_ ),
    .B1(\u_cpu.ALU.u_wallace._3437_ ),
    .Y(\u_cpu.ALU.u_wallace._3448_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5253_  (.A(\u_cpu.ALU.u_wallace._3119_ ),
    .B(\u_cpu.ALU.u_wallace._3010_ ),
    .Y(\u_cpu.ALU.u_wallace._3459_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5254_  (.A1(\u_cpu.ALU.u_wallace._3021_ ),
    .A2(\u_cpu.ALU.u_wallace._3459_ ),
    .B1(\u_cpu.ALU.u_wallace._3382_ ),
    .C1(\u_cpu.ALU.u_wallace._3426_ ),
    .X(\u_cpu.ALU.u_wallace._3470_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5255_  (.A(\u_cpu.ALU.u_wallace._3404_ ),
    .X(\u_cpu.ALU.u_wallace._3481_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5256_  (.A(\u_cpu.ALU.u_wallace._0512_ ),
    .B(\u_cpu.ALU.u_wallace._2045_ ),
    .C(\u_cpu.ALU.u_wallace._1552_ ),
    .D(\u_cpu.ALU.u_wallace._1191_ ),
    .X(\u_cpu.ALU.u_wallace._3492_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._5257_  (.A1(\u_cpu.ALU.u_wallace._2560_ ),
    .A2(\u_cpu.ALU.u_wallace._3481_ ),
    .A3(\u_cpu.ALU.u_wallace._0994_ ),
    .B1(\u_cpu.ALU.u_wallace._3492_ ),
    .X(\u_cpu.ALU.u_wallace._3503_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._5258_  (.A1(\u_cpu.ALU.u_wallace._3448_ ),
    .A2(\u_cpu.ALU.u_wallace._3470_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3503_ ),
    .Y(\u_cpu.ALU.u_wallace._3514_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5259_  (.A(\u_cpu.ALU.u_wallace._0906_ ),
    .B(\u_cpu.ALU.u_wallace._1530_ ),
    .C(\u_cpu.ALU.u_wallace._1552_ ),
    .D(\u_cpu.ALU.u_wallace._1191_ ),
    .Y(\u_cpu.ALU.u_wallace._3525_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5260_  (.A1(\u_cpu.ALU.u_wallace._0261_ ),
    .A2(\u_cpu.ALU.u_wallace._2626_ ),
    .B1(\u_cpu.ALU.u_wallace._3415_ ),
    .B2(\u_cpu.ALU.u_wallace._3525_ ),
    .Y(\u_cpu.ALU.u_wallace._3536_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5261_  (.A1(\u_cpu.ALU.u_wallace._1037_ ),
    .A2(\u_cpu.ALU.u_wallace._3393_ ),
    .B1(\u_cpu.ALU.u_wallace._3371_ ),
    .C1(\u_cpu.ALU.u_wallace._3415_ ),
    .X(\u_cpu.ALU.u_wallace._3547_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._5262_  (.A1(\u_cpu.ALU.u_wallace._3536_ ),
    .A2(\u_cpu.ALU.u_wallace._3547_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3437_ ),
    .Y(\u_cpu.ALU.u_wallace._3558_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5263_  (.A1(\u_cpu.ALU.u_wallace._3021_ ),
    .A2(\u_cpu.ALU.u_wallace._3459_ ),
    .B1(\u_cpu.ALU.u_wallace._3382_ ),
    .C1(\u_cpu.ALU.u_wallace._3426_ ),
    .Y(\u_cpu.ALU.u_wallace._3569_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5264_  (.A(\u_cpu.ALU.u_wallace._3558_ ),
    .B(\u_cpu.ALU.u_wallace._3569_ ),
    .C(\u_cpu.ALU.u_wallace._3503_ ),
    .Y(\u_cpu.ALU.u_wallace._3580_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5265_  (.A1(\u_cpu.ALU.u_wallace._3010_ ),
    .A2(\u_cpu.ALU.u_wallace._3130_ ),
    .B1(\u_cpu.ALU.u_wallace._3032_ ),
    .C1(\u_cpu.ALU.u_wallace._2911_ ),
    .X(\u_cpu.ALU.u_wallace._3591_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5266_  (.A(\u_cpu.ALU.u_wallace._1859_ ),
    .B(\u_cpu.ALU.u_wallace._2725_ ),
    .Y(\u_cpu.ALU.u_wallace._3602_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5267_  (.A(\u_cpu.ALU.u_wallace._1826_ ),
    .B(\u_cpu.ALU.u_wallace._0250_ ),
    .Y(\u_cpu.ALU.u_wallace._3613_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5268_  (.A(\u_cpu.ALU.SrcA[8] ),
    .X(\u_cpu.ALU.u_wallace._3623_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5269_  (.A1(\u_cpu.ALU.u_wallace._1771_ ),
    .A2(\u_cpu.ALU.u_wallace._0348_ ),
    .B1(\u_cpu.ALU.u_wallace._3623_ ),
    .B2(\u_cpu.ALU.u_wallace._1749_ ),
    .Y(\u_cpu.ALU.u_wallace._3634_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5270_  (.A(\u_cpu.ALU.SrcA[8] ),
    .X(\u_cpu.ALU.u_wallace._3645_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5271_  (.A(\u_cpu.ALU.u_wallace._0862_ ),
    .B(\u_cpu.ALU.u_wallace._2768_ ),
    .C(\u_cpu.ALU.SrcA[2] ),
    .D(\u_cpu.ALU.u_wallace._3645_ ),
    .X(\u_cpu.ALU.u_wallace._3656_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5272_  (.A1(\u_cpu.ALU.u_wallace._3602_ ),
    .A2(\u_cpu.ALU.u_wallace._3613_ ),
    .B1(\u_cpu.ALU.u_wallace._3634_ ),
    .B2(\u_cpu.ALU.u_wallace._3656_ ),
    .Y(\u_cpu.ALU.u_wallace._3667_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5273_  (.A(\u_cpu.ALU.SrcB[6] ),
    .X(\u_cpu.ALU.u_wallace._3678_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5274_  (.A(\u_cpu.ALU.SrcA[8] ),
    .X(\u_cpu.ALU.u_wallace._3689_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5275_  (.A1(\u_cpu.ALU.u_wallace._3678_ ),
    .A2(\u_cpu.ALU.u_wallace._0392_ ),
    .B1(\u_cpu.ALU.u_wallace._3689_ ),
    .B2(\u_cpu.ALU.u_wallace._0862_ ),
    .X(\u_cpu.ALU.u_wallace._3700_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5276_  (.A(\u_cpu.ALU.u_wallace._2747_ ),
    .B(\u_cpu.ALU.u_wallace._2856_ ),
    .C(\u_cpu.ALU.u_wallace._0392_ ),
    .D(\u_cpu.ALU.u_wallace._3689_ ),
    .Y(\u_cpu.ALU.u_wallace._3711_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5277_  (.A(\u_cpu.ALU.u_wallace._2900_ ),
    .B(\u_cpu.ALU.u_wallace._3700_ ),
    .C(\u_cpu.ALU.u_wallace._3711_ ),
    .Y(\u_cpu.ALU.u_wallace._3722_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5278_  (.A1(\u_cpu.ALU.u_wallace._2790_ ),
    .A2(\u_cpu.ALU.u_wallace._0797_ ),
    .B1(\u_cpu.ALU.u_wallace._1914_ ),
    .B2(\u_cpu.ALU.u_wallace._1837_ ),
    .Y(\u_cpu.ALU.u_wallace._3733_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5279_  (.A(\u_cpu.ALU.u_wallace._2790_ ),
    .B(\u_cpu.ALU.u_wallace._1903_ ),
    .C(\u_cpu.ALU.u_wallace._0807_ ),
    .D(\u_cpu.ALU.u_wallace._1837_ ),
    .X(\u_cpu.ALU.u_wallace._3744_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5280_  (.A(\u_cpu.ALU.u_wallace._0457_ ),
    .B(\u_cpu.ALU.u_wallace._2955_ ),
    .Y(\u_cpu.ALU.u_wallace._3755_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5281_  (.A1(\u_cpu.ALU.u_wallace._3733_ ),
    .A2(\u_cpu.ALU.u_wallace._3744_ ),
    .B1(\u_cpu.ALU.u_wallace._3755_ ),
    .Y(\u_cpu.ALU.u_wallace._3766_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5282_  (.A(\u_cpu.ALU.u_wallace._1782_ ),
    .X(\u_cpu.ALU.u_wallace._3777_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5283_  (.A(\u_cpu.ALU.u_wallace._2725_ ),
    .B(\u_cpu.ALU.u_wallace._1957_ ),
    .C(\u_cpu.ALU.u_wallace._1968_ ),
    .D(\u_cpu.ALU.u_wallace._3777_ ),
    .Y(\u_cpu.ALU.u_wallace._3788_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._5284_  (.A_N(\u_cpu.ALU.u_wallace._3733_ ),
    .B(\u_cpu.ALU.u_wallace._3788_ ),
    .C(\u_cpu.ALU.u_wallace._0468_ ),
    .D(\u_cpu.ALU.u_wallace._1322_ ),
    .Y(\u_cpu.ALU.u_wallace._3799_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5285_  (.A1(\u_cpu.ALU.u_wallace._3667_ ),
    .A2(\u_cpu.ALU.u_wallace._3722_ ),
    .B1(\u_cpu.ALU.u_wallace._3766_ ),
    .B2(\u_cpu.ALU.u_wallace._3799_ ),
    .X(\u_cpu.ALU.u_wallace._3810_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5286_  (.A(\u_cpu.ALU.u_wallace._2878_ ),
    .X(\u_cpu.ALU.u_wallace._3821_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5287_  (.A(\u_cpu.ALU.u_wallace._1782_ ),
    .X(\u_cpu.ALU.u_wallace._3832_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._5288_  (.A1(\u_cpu.ALU.u_wallace._3821_ ),
    .A2(\u_cpu.ALU.u_wallace._1158_ ),
    .A3(\u_cpu.ALU.u_wallace._0304_ ),
    .A4(\u_cpu.ALU.u_wallace._3832_ ),
    .B1(\u_cpu.ALU.u_wallace._3755_ ),
    .X(\u_cpu.ALU.u_wallace._3843_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._5289_  (.A1(\u_cpu.ALU.u_wallace._3843_ ),
    .A2(\u_cpu.ALU.u_wallace._3733_ ),
    .B1(\u_cpu.ALU.u_wallace._3722_ ),
    .C1(\u_cpu.ALU.u_wallace._3667_ ),
    .D1(\u_cpu.ALU.u_wallace._3766_ ),
    .Y(\u_cpu.ALU.u_wallace._3854_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5290_  (.A1(\u_cpu.ALU.u_wallace._3108_ ),
    .A2(\u_cpu.ALU.u_wallace._3591_ ),
    .B1(\u_cpu.ALU.u_wallace._3810_ ),
    .C1(\u_cpu.ALU.u_wallace._3854_ ),
    .Y(\u_cpu.ALU.u_wallace._3865_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5291_  (.A1(\u_cpu.ALU.u_wallace._3667_ ),
    .A2(\u_cpu.ALU.u_wallace._3722_ ),
    .B1(\u_cpu.ALU.u_wallace._3766_ ),
    .B2(\u_cpu.ALU.u_wallace._3799_ ),
    .Y(\u_cpu.ALU.u_wallace._3876_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._5292_  (.A1(\u_cpu.ALU.u_wallace._3843_ ),
    .A2(\u_cpu.ALU.u_wallace._3733_ ),
    .B1(\u_cpu.ALU.u_wallace._3722_ ),
    .C1(\u_cpu.ALU.u_wallace._3667_ ),
    .D1(\u_cpu.ALU.u_wallace._3766_ ),
    .X(\u_cpu.ALU.u_wallace._3887_ ));
 sky130_fd_sc_hd__o41a_2 \u_cpu.ALU.u_wallace._5293_  (.A1(\u_cpu.ALU.u_wallace._2845_ ),
    .A2(\u_cpu.ALU.u_wallace._2867_ ),
    .A3(\u_cpu.ALU.u_wallace._2889_ ),
    .A4(\u_cpu.ALU.u_wallace._2900_ ),
    .B1(\u_cpu.ALU.u_wallace._3141_ ),
    .X(\u_cpu.ALU.u_wallace._3898_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5294_  (.A1(\u_cpu.ALU.u_wallace._3876_ ),
    .A2(\u_cpu.ALU.u_wallace._3887_ ),
    .B1(\u_cpu.ALU.u_wallace._3898_ ),
    .Y(\u_cpu.ALU.u_wallace._3908_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5295_  (.A1(\u_cpu.ALU.u_wallace._3514_ ),
    .A2(\u_cpu.ALU.u_wallace._3580_ ),
    .B1(\u_cpu.ALU.u_wallace._3865_ ),
    .B2(\u_cpu.ALU.u_wallace._3908_ ),
    .X(\u_cpu.ALU.u_wallace._3919_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5296_  (.A(\u_cpu.ALU.u_wallace._3558_ ),
    .B(\u_cpu.ALU.u_wallace._3503_ ),
    .Y(\u_cpu.ALU.u_wallace._3930_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._5297_  (.A1(\u_cpu.ALU.u_wallace._3470_ ),
    .A2(\u_cpu.ALU.u_wallace._3930_ ),
    .B1(\u_cpu.ALU.u_wallace._3865_ ),
    .C1(\u_cpu.ALU.u_wallace._3908_ ),
    .D1(\u_cpu.ALU.u_wallace._3514_ ),
    .Y(\u_cpu.ALU.u_wallace._3941_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5298_  (.A(\u_cpu.ALU.u_wallace._3338_ ),
    .B(\u_cpu.ALU.u_wallace._3919_ ),
    .C(\u_cpu.ALU.u_wallace._3941_ ),
    .Y(\u_cpu.ALU.u_wallace._3952_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5299_  (.A1(\u_cpu.ALU.u_wallace._3514_ ),
    .A2(\u_cpu.ALU.u_wallace._3580_ ),
    .B1(\u_cpu.ALU.u_wallace._3865_ ),
    .B2(\u_cpu.ALU.u_wallace._3908_ ),
    .Y(\u_cpu.ALU.u_wallace._3963_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._5300_  (.A1(\u_cpu.ALU.u_wallace._3930_ ),
    .A2(\u_cpu.ALU.u_wallace._3470_ ),
    .B1(\u_cpu.ALU.u_wallace._3514_ ),
    .C1(\u_cpu.ALU.u_wallace._3865_ ),
    .D1(\u_cpu.ALU.u_wallace._3908_ ),
    .X(\u_cpu.ALU.u_wallace._3974_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._5301_  (.A1(\u_cpu.ALU.u_wallace._3064_ ),
    .A2(\u_cpu.ALU.u_wallace._3185_ ),
    .B1(\u_cpu.ALU.u_wallace._3963_ ),
    .B2(\u_cpu.ALU.u_wallace._3974_ ),
    .C1(\u_cpu.ALU.u_wallace._3152_ ),
    .Y(\u_cpu.ALU.u_wallace._3985_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5302_  (.A(\u_cpu.ALU.u_wallace._1070_ ),
    .X(\u_cpu.ALU.u_wallace._3996_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5303_  (.A(\u_cpu.ALU.SrcB[8] ),
    .X(\u_cpu.ALU.u_wallace._4007_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5304_  (.A(\u_cpu.ALU.u_wallace._4007_ ),
    .X(\u_cpu.ALU.u_wallace._4018_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5305_  (.A(\u_cpu.ALU.u_wallace._4018_ ),
    .X(\u_cpu.ALU.u_wallace._4029_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5306_  (.A(\u_cpu.ALU.u_wallace._3996_ ),
    .B(\u_cpu.ALU.u_wallace._4029_ ),
    .Y(\u_cpu.ALU.u_wallace._4040_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5307_  (.A1(\u_cpu.ALU.u_wallace._2703_ ),
    .A2(\u_cpu.ALU.u_wallace._2714_ ),
    .B1(\u_cpu.ALU.u_wallace._4040_ ),
    .Y(\u_cpu.ALU.u_wallace._4051_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5308_  (.A(\u_cpu.ALU.u_wallace._0370_ ),
    .B(\u_cpu.ALU.u_wallace._2166_ ),
    .Y(\u_cpu.ALU.u_wallace._4062_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5309_  (.A(\u_cpu.ALU.u_wallace._0173_ ),
    .B(\u_cpu.ALU.u_wallace._2198_ ),
    .Y(\u_cpu.ALU.u_wallace._4073_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU.u_wallace._5310_  (.A1(\u_cpu.ALU.u_wallace._4062_ ),
    .A2(\u_cpu.ALU.u_wallace._4073_ ),
    .A3(\u_cpu.ALU.u_wallace._2670_ ),
    .B1(\u_cpu.ALU.u_wallace._4040_ ),
    .C1(\u_cpu.ALU.u_wallace._2703_ ),
    .X(\u_cpu.ALU.u_wallace._4084_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5311_  (.A(\u_cpu.ALU.u_wallace._4051_ ),
    .B(\u_cpu.ALU.u_wallace._4084_ ),
    .Y(\u_cpu.ALU.u_wallace._4095_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5312_  (.A1(\u_cpu.ALU.u_wallace._3952_ ),
    .A2(\u_cpu.ALU.u_wallace._3985_ ),
    .B1(\u_cpu.ALU.u_wallace._4095_ ),
    .Y(\u_cpu.ALU.u_wallace._4106_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5313_  (.A(\u_cpu.ALU.u_wallace._3985_ ),
    .B(\u_cpu.ALU.u_wallace._4095_ ),
    .C(\u_cpu.ALU.u_wallace._3952_ ),
    .X(\u_cpu.ALU.u_wallace._4117_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._5314_  (.A1(\u_cpu.ALU.u_wallace._3196_ ),
    .A2(\u_cpu.ALU.u_wallace._3218_ ),
    .B1(\u_cpu.ALU.u_wallace._4106_ ),
    .C1(\u_cpu.ALU.u_wallace._4117_ ),
    .X(\u_cpu.ALU.u_wallace._4128_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5315_  (.A1(\u_cpu.ALU.u_wallace._4106_ ),
    .A2(\u_cpu.ALU.u_wallace._4117_ ),
    .B1(\u_cpu.ALU.u_wallace._3196_ ),
    .C1(\u_cpu.ALU.u_wallace._3218_ ),
    .Y(\u_cpu.ALU.u_wallace._4139_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._5316_  (.A1(\u_cpu.ALU.u_wallace._3295_ ),
    .A2(\u_cpu.ALU.u_wallace._3262_ ),
    .B1(\u_cpu.ALU.u_wallace._3328_ ),
    .C1(\u_cpu.ALU.u_wallace._4128_ ),
    .D1(\u_cpu.ALU.u_wallace._4139_ ),
    .Y(\u_cpu.ALU.u_wallace._4150_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU.u_wallace._5317_  (.A1(\u_cpu.ALU.u_wallace._3196_ ),
    .A2(\u_cpu.ALU.u_wallace._3218_ ),
    .B1(\u_cpu.ALU.u_wallace._4106_ ),
    .C1(\u_cpu.ALU.u_wallace._4117_ ),
    .Y(\u_cpu.ALU.u_wallace._4161_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5318_  (.A1(\u_cpu.ALU.u_wallace._4106_ ),
    .A2(\u_cpu.ALU.u_wallace._4117_ ),
    .B1(\u_cpu.ALU.u_wallace._3196_ ),
    .C1(\u_cpu.ALU.u_wallace._3218_ ),
    .X(\u_cpu.ALU.u_wallace._4172_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5319_  (.A1(\u_cpu.ALU.u_wallace._3262_ ),
    .A2(\u_cpu.ALU.u_wallace._3295_ ),
    .B1(\u_cpu.ALU.u_wallace._3328_ ),
    .Y(\u_cpu.ALU.u_wallace._4183_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5320_  (.A1(\u_cpu.ALU.u_wallace._4161_ ),
    .A2(\u_cpu.ALU.u_wallace._4172_ ),
    .B1(\u_cpu.ALU.u_wallace._4183_ ),
    .Y(\u_cpu.ALU.u_wallace._4194_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5321_  (.A(\u_cpu.ALU.u_wallace._2462_ ),
    .B(\u_cpu.ALU.u_wallace._3273_ ),
    .Y(\u_cpu.ALU.u_wallace._4205_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5322_  (.A(\u_cpu.ALU.u_wallace._4150_ ),
    .B(\u_cpu.ALU.u_wallace._4194_ ),
    .C(\u_cpu.ALU.u_wallace._4205_ ),
    .Y(\u_cpu.ALU.u_wallace._4215_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5323_  (.A1(\u_cpu.ALU.u_wallace._4150_ ),
    .A2(\u_cpu.ALU.u_wallace._4194_ ),
    .B1(\u_cpu.ALU.u_wallace._4205_ ),
    .X(\u_cpu.ALU.u_wallace._4226_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5324_  (.A1(\u_cpu.ALU.u_wallace._2494_ ),
    .A2(\u_cpu.ALU.u_wallace._3317_ ),
    .B1(\u_cpu.ALU.u_wallace._4226_ ),
    .B2(\u_cpu.ALU.u_wallace._4215_ ),
    .Y(\u_cpu.ALU.u_wallace._4237_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._5325_  (.A1(\u_cpu.ALU.u_wallace._2494_ ),
    .A2(\u_cpu.ALU.u_wallace._3317_ ),
    .A3(\u_cpu.ALU.u_wallace._4215_ ),
    .B1(\u_cpu.ALU.u_wallace._4237_ ),
    .Y(\u_cpu.ALU.Product_Wallace[8] ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5326_  (.A(\u_cpu.ALU.u_wallace._4215_ ),
    .B(\u_cpu.ALU.u_wallace._2494_ ),
    .C(\u_cpu.ALU.u_wallace._3317_ ),
    .Y(\u_cpu.ALU.u_wallace._4258_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5327_  (.A(\u_cpu.ALU.u_wallace._4226_ ),
    .B(\u_cpu.ALU.u_wallace._4258_ ),
    .Y(\u_cpu.ALU.u_wallace._4269_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._5328_  (.A1(\u_cpu.ALU.u_wallace._3985_ ),
    .A2(\u_cpu.ALU.u_wallace._4095_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3952_ ),
    .Y(\u_cpu.ALU.u_wallace._4280_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5329_  (.A(\u_cpu.ALU.SrcB[9] ),
    .X(\u_cpu.ALU.u_wallace._4291_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5330_  (.A(\u_cpu.ALU.u_wallace._4291_ ),
    .X(\u_cpu.ALU.u_wallace._4302_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5331_  (.A(\u_cpu.ALU.u_wallace._4302_ ),
    .X(\u_cpu.ALU.u_wallace._4313_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5332_  (.A1(\u_cpu.ALU.u_wallace._0272_ ),
    .A2(\u_cpu.ALU.u_wallace._4029_ ),
    .B1(\u_cpu.ALU.u_wallace._4313_ ),
    .B2(\u_cpu.ALU.u_wallace._1070_ ),
    .Y(\u_cpu.ALU.u_wallace._4324_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5333_  (.A(\u_cpu.ALU.u_wallace._0108_ ),
    .B(\u_cpu.ALU.u_wallace._0162_ ),
    .C(\u_cpu.ALU.u_wallace._4029_ ),
    .D(\u_cpu.ALU.u_wallace._4313_ ),
    .X(\u_cpu.ALU.u_wallace._4335_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5334_  (.A(\u_cpu.ALU.u_wallace._4324_ ),
    .B(\u_cpu.ALU.u_wallace._4335_ ),
    .Y(\u_cpu.ALU.u_wallace._4346_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5335_  (.A1(\u_cpu.ALU.u_wallace._3569_ ),
    .A2(\u_cpu.ALU.u_wallace._3930_ ),
    .B1(\u_cpu.ALU.u_wallace._4346_ ),
    .X(\u_cpu.ALU.u_wallace._4357_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5336_  (.A(\u_cpu.ALU.u_wallace._3569_ ),
    .B(\u_cpu.ALU.u_wallace._3930_ ),
    .C(\u_cpu.ALU.u_wallace._4346_ ),
    .Y(\u_cpu.ALU.u_wallace._4368_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5337_  (.A(\u_cpu.ALU.u_wallace._2900_ ),
    .B(\u_cpu.ALU.u_wallace._3700_ ),
    .C(\u_cpu.ALU.u_wallace._3711_ ),
    .X(\u_cpu.ALU.u_wallace._4379_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._5338_  (.A1(\u_cpu.ALU.u_wallace._3667_ ),
    .A2(\u_cpu.ALU.u_wallace._3766_ ),
    .A3(\u_cpu.ALU.u_wallace._3799_ ),
    .B1(\u_cpu.ALU.u_wallace._4379_ ),
    .X(\u_cpu.ALU.u_wallace._4390_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5339_  (.A(\u_cpu.ALU.SrcA[9] ),
    .X(\u_cpu.ALU.u_wallace._4401_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5340_  (.A(\u_cpu.ALU.u_wallace._4401_ ),
    .X(\u_cpu.ALU.u_wallace._4412_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5341_  (.A1(\u_cpu.ALU.u_wallace._2856_ ),
    .A2(\u_cpu.ALU.u_wallace._2549_ ),
    .B1(\u_cpu.ALU.u_wallace._4412_ ),
    .B2(\u_cpu.ALU.u_wallace._2747_ ),
    .Y(\u_cpu.ALU.u_wallace._4423_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5342_  (.A(\u_cpu.ALU.u_wallace._1760_ ),
    .X(\u_cpu.ALU.u_wallace._4431_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5343_  (.A(\u_cpu.ALU.u_wallace._4401_ ),
    .X(\u_cpu.ALU.u_wallace._4439_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5344_  (.A(\u_cpu.ALU.u_wallace._1749_ ),
    .B(\u_cpu.ALU.u_wallace._4431_ ),
    .C(\u_cpu.ALU.u_wallace._1278_ ),
    .D(\u_cpu.ALU.u_wallace._4439_ ),
    .Y(\u_cpu.ALU.u_wallace._4442_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._5345_  (.A_N(\u_cpu.ALU.u_wallace._4423_ ),
    .B(\u_cpu.ALU.u_wallace._4442_ ),
    .C(\u_cpu.ALU.u_wallace._3656_ ),
    .Y(\u_cpu.ALU.u_wallace._4443_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5346_  (.A(\u_cpu.ALU.SrcA[9] ),
    .X(\u_cpu.ALU.u_wallace._4444_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5347_  (.A(\u_cpu.ALU.u_wallace._0862_ ),
    .B(\u_cpu.ALU.u_wallace._3678_ ),
    .C(\u_cpu.ALU.u_wallace._0764_ ),
    .D(\u_cpu.ALU.u_wallace._4444_ ),
    .X(\u_cpu.ALU.u_wallace._4445_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5348_  (.A1(\u_cpu.ALU.u_wallace._4423_ ),
    .A2(\u_cpu.ALU.u_wallace._4445_ ),
    .B1(\u_cpu.ALU.u_wallace._3711_ ),
    .Y(\u_cpu.ALU.u_wallace._4446_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5349_  (.A(\u_cpu.ALU.SrcA[7] ),
    .X(\u_cpu.ALU.u_wallace._4447_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5350_  (.A1(\u_cpu.ALU.u_wallace._3689_ ),
    .A2(\u_cpu.ALU.u_wallace._0479_ ),
    .B1(\u_cpu.ALU.u_wallace._0490_ ),
    .B2(\u_cpu.ALU.u_wallace._4447_ ),
    .Y(\u_cpu.ALU.u_wallace._4448_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5351_  (.A(\u_cpu.ALU.SrcA[8] ),
    .X(\u_cpu.ALU.u_wallace._4449_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5352_  (.A(\u_cpu.ALU.SrcA[7] ),
    .X(\u_cpu.ALU.u_wallace._4450_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5353_  (.A(\u_cpu.ALU.u_wallace._4449_ ),
    .B(\u_cpu.ALU.u_wallace._4450_ ),
    .C(\u_cpu.ALU.u_wallace._1957_ ),
    .D(\u_cpu.ALU.u_wallace._1968_ ),
    .Y(\u_cpu.ALU.u_wallace._4451_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5354_  (.A(\u_cpu.ALU.u_wallace._2834_ ),
    .X(\u_cpu.ALU.u_wallace._4452_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._5355_  (.A_N(\u_cpu.ALU.u_wallace._4448_ ),
    .B(\u_cpu.ALU.u_wallace._4451_ ),
    .C(\u_cpu.ALU.u_wallace._4452_ ),
    .D(\u_cpu.ALU.u_wallace._0468_ ),
    .Y(\u_cpu.ALU.u_wallace._4453_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._5356_  (.A(\u_cpu.ALU.u_wallace._1782_ ),
    .Y(\u_cpu.ALU.u_wallace._4454_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5357_  (.A(\u_cpu.ALU.u_wallace._3689_ ),
    .B(\u_cpu.ALU.u_wallace._2790_ ),
    .C(\u_cpu.ALU.u_wallace._0479_ ),
    .D(\u_cpu.ALU.u_wallace._1914_ ),
    .X(\u_cpu.ALU.u_wallace._4455_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5358_  (.A1(\u_cpu.ALU.u_wallace._4454_ ),
    .A2(\u_cpu.ALU.u_wallace._1892_ ),
    .B1(\u_cpu.ALU.u_wallace._4448_ ),
    .B2(\u_cpu.ALU.u_wallace._4455_ ),
    .Y(\u_cpu.ALU.u_wallace._4456_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5359_  (.A1(\u_cpu.ALU.u_wallace._4443_ ),
    .A2(\u_cpu.ALU.u_wallace._4446_ ),
    .B1(\u_cpu.ALU.u_wallace._4453_ ),
    .B2(\u_cpu.ALU.u_wallace._4456_ ),
    .X(\u_cpu.ALU.u_wallace._4457_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5360_  (.A(\u_cpu.ALU.u_wallace._4443_ ),
    .B(\u_cpu.ALU.u_wallace._4446_ ),
    .C(\u_cpu.ALU.u_wallace._4453_ ),
    .D(\u_cpu.ALU.u_wallace._4456_ ),
    .Y(\u_cpu.ALU.u_wallace._4458_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5361_  (.A(\u_cpu.ALU.u_wallace._4390_ ),
    .B(\u_cpu.ALU.u_wallace._4457_ ),
    .C(\u_cpu.ALU.u_wallace._4458_ ),
    .Y(\u_cpu.ALU.u_wallace._4459_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5362_  (.A1(\u_cpu.ALU.u_wallace._4443_ ),
    .A2(\u_cpu.ALU.u_wallace._4446_ ),
    .B1(\u_cpu.ALU.u_wallace._4453_ ),
    .B2(\u_cpu.ALU.u_wallace._4456_ ),
    .Y(\u_cpu.ALU.u_wallace._4460_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5363_  (.A(\u_cpu.ALU.u_wallace._4443_ ),
    .B(\u_cpu.ALU.u_wallace._4446_ ),
    .C(\u_cpu.ALU.u_wallace._4453_ ),
    .D(\u_cpu.ALU.u_wallace._4456_ ),
    .X(\u_cpu.ALU.u_wallace._4461_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._5364_  (.A1(\u_cpu.ALU.u_wallace._4460_ ),
    .A2(\u_cpu.ALU.u_wallace._4461_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4390_ ),
    .Y(\u_cpu.ALU.u_wallace._4462_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5365_  (.A(\u_cpu.ALU.u_wallace._0731_ ),
    .X(\u_cpu.ALU.u_wallace._4463_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5366_  (.A(\u_cpu.ALU.u_wallace._3415_ ),
    .B(\u_cpu.ALU.u_wallace._3481_ ),
    .C(\u_cpu.ALU.u_wallace._4463_ ),
    .X(\u_cpu.ALU.u_wallace._4464_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5367_  (.A(\u_cpu.ALU.u_wallace._1125_ ),
    .B(\u_cpu.ALU.u_wallace._1180_ ),
    .C(\u_cpu.ALU.u_wallace._2045_ ),
    .D(\u_cpu.ALU.u_wallace._2056_ ),
    .Y(\u_cpu.ALU.u_wallace._4465_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5368_  (.A(\u_cpu.ALU.u_wallace._4465_ ),
    .B(\u_cpu.ALU.u_wallace._2626_ ),
    .C(\u_cpu.ALU.u_wallace._0359_ ),
    .Y(\u_cpu.ALU.u_wallace._4466_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5369_  (.A(\u_cpu.ALU.SrcB[4] ),
    .X(\u_cpu.ALU.u_wallace._4467_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5370_  (.A1(\u_cpu.ALU.u_wallace._2955_ ),
    .A2(\u_cpu.ALU.u_wallace._4467_ ),
    .B1(\u_cpu.ALU.u_wallace._2078_ ),
    .B2(\u_cpu.ALU.u_wallace._2922_ ),
    .Y(\u_cpu.ALU.u_wallace._4468_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5371_  (.A1(\u_cpu.ALU.u_wallace._3755_ ),
    .A2(\u_cpu.ALU.u_wallace._3733_ ),
    .B1(\u_cpu.ALU.u_wallace._3788_ ),
    .Y(\u_cpu.ALU.u_wallace._4469_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._5372_  (.A(\u_cpu.ALU.SrcB[7] ),
    .Y(\u_cpu.ALU.u_wallace._4470_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5373_  (.A(\u_cpu.ALU.u_wallace._4470_ ),
    .X(\u_cpu.ALU.u_wallace._4471_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5374_  (.A(\u_cpu.ALU.u_wallace._1311_ ),
    .B(\u_cpu.ALU.u_wallace._0895_ ),
    .C(\u_cpu.ALU.u_wallace._2144_ ),
    .D(\u_cpu.ALU.u_wallace._2538_ ),
    .X(\u_cpu.ALU.u_wallace._4472_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5375_  (.A1(\u_cpu.ALU.u_wallace._0403_ ),
    .A2(\u_cpu.ALU.u_wallace._4471_ ),
    .B1(\u_cpu.ALU.u_wallace._4468_ ),
    .B2(\u_cpu.ALU.u_wallace._4472_ ),
    .Y(\u_cpu.ALU.u_wallace._4473_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5376_  (.A1(\u_cpu.ALU.u_wallace._4466_ ),
    .A2(\u_cpu.ALU.u_wallace._4468_ ),
    .B1(\u_cpu.ALU.u_wallace._4469_ ),
    .C1(\u_cpu.ALU.u_wallace._4473_ ),
    .Y(\u_cpu.ALU.u_wallace._4474_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5377_  (.A1(\u_cpu.ALU.u_wallace._1979_ ),
    .A2(\u_cpu.ALU.u_wallace._2571_ ),
    .B1(\u_cpu.ALU.u_wallace._2582_ ),
    .B2(\u_cpu.ALU.u_wallace._1267_ ),
    .X(\u_cpu.ALU.u_wallace._4475_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5378_  (.A(\u_cpu.ALU.u_wallace._4475_ ),
    .B(\u_cpu.ALU.u_wallace._4465_ ),
    .C(\u_cpu.ALU.u_wallace._0359_ ),
    .D(\u_cpu.ALU.u_wallace._2604_ ),
    .Y(\u_cpu.ALU.u_wallace._4476_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5379_  (.A1(\u_cpu.ALU.u_wallace._4476_ ),
    .A2(\u_cpu.ALU.u_wallace._4473_ ),
    .B1(\u_cpu.ALU.u_wallace._4469_ ),
    .X(\u_cpu.ALU.u_wallace._4477_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5380_  (.A1(\u_cpu.ALU.u_wallace._3360_ ),
    .A2(\u_cpu.ALU.u_wallace._4464_ ),
    .B1(\u_cpu.ALU.u_wallace._4474_ ),
    .C1(\u_cpu.ALU.u_wallace._4477_ ),
    .X(\u_cpu.ALU.u_wallace._4478_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5381_  (.A1(\u_cpu.ALU.u_wallace._4466_ ),
    .A2(\u_cpu.ALU.u_wallace._4468_ ),
    .B1(\u_cpu.ALU.u_wallace._4469_ ),
    .C1(\u_cpu.ALU.u_wallace._4473_ ),
    .X(\u_cpu.ALU.u_wallace._4479_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5382_  (.A1(\u_cpu.ALU.u_wallace._4476_ ),
    .A2(\u_cpu.ALU.u_wallace._4473_ ),
    .B1(\u_cpu.ALU.u_wallace._4469_ ),
    .Y(\u_cpu.ALU.u_wallace._4480_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU.u_wallace._5383_  (.A1_N(\u_cpu.ALU.u_wallace._3371_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3415_ ),
    .B1(\u_cpu.ALU.u_wallace._1037_ ),
    .B2(\u_cpu.ALU.u_wallace._3393_ ),
    .X(\u_cpu.ALU.u_wallace._4481_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._5384_  (.A1(\u_cpu.ALU.u_wallace._4479_ ),
    .A2(\u_cpu.ALU.u_wallace._4480_ ),
    .B1(\u_cpu.ALU.u_wallace._4481_ ),
    .X(\u_cpu.ALU.u_wallace._4482_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5385_  (.A1_N(\u_cpu.ALU.u_wallace._4459_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4462_ ),
    .B1(\u_cpu.ALU.u_wallace._4478_ ),
    .B2(\u_cpu.ALU.u_wallace._4482_ ),
    .Y(\u_cpu.ALU.u_wallace._4483_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5386_  (.A1(\u_cpu.ALU.u_wallace._3360_ ),
    .A2(\u_cpu.ALU.u_wallace._4464_ ),
    .B1(\u_cpu.ALU.u_wallace._4479_ ),
    .B2(\u_cpu.ALU.u_wallace._4480_ ),
    .Y(\u_cpu.ALU.u_wallace._4484_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5387_  (.A(\u_cpu.ALU.u_wallace._4477_ ),
    .B(\u_cpu.ALU.u_wallace._4481_ ),
    .C(\u_cpu.ALU.u_wallace._4474_ ),
    .Y(\u_cpu.ALU.u_wallace._4485_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5388_  (.A(\u_cpu.ALU.u_wallace._4484_ ),
    .B(\u_cpu.ALU.u_wallace._4485_ ),
    .Y(\u_cpu.ALU.u_wallace._4486_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5389_  (.A(\u_cpu.ALU.u_wallace._4459_ ),
    .B(\u_cpu.ALU.u_wallace._4462_ ),
    .C(\u_cpu.ALU.u_wallace._4486_ ),
    .Y(\u_cpu.ALU.u_wallace._4487_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5390_  (.A1(\u_cpu.ALU.u_wallace._3930_ ),
    .A2(\u_cpu.ALU.u_wallace._3470_ ),
    .B1(\u_cpu.ALU.u_wallace._3514_ ),
    .C1(\u_cpu.ALU.u_wallace._3908_ ),
    .Y(\u_cpu.ALU.u_wallace._4488_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5391_  (.A(\u_cpu.ALU.u_wallace._3865_ ),
    .B(\u_cpu.ALU.u_wallace._4488_ ),
    .Y(\u_cpu.ALU.u_wallace._4489_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5392_  (.A1(\u_cpu.ALU.u_wallace._4483_ ),
    .A2(\u_cpu.ALU.u_wallace._4487_ ),
    .B1(\u_cpu.ALU.u_wallace._4489_ ),
    .Y(\u_cpu.ALU.u_wallace._4490_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5393_  (.A1(\u_cpu.ALU.u_wallace._4357_ ),
    .A2(\u_cpu.ALU.u_wallace._4368_ ),
    .B1(\u_cpu.ALU.u_wallace._4490_ ),
    .Y(\u_cpu.ALU.u_wallace._4491_ ));
 sky130_fd_sc_hd__a32oi_2 \u_cpu.ALU.u_wallace._5394_  (.A1(\u_cpu.ALU.u_wallace._4459_ ),
    .A2(\u_cpu.ALU.u_wallace._4462_ ),
    .A3(\u_cpu.ALU.u_wallace._4486_ ),
    .B1(\u_cpu.ALU.u_wallace._4488_ ),
    .B2(\u_cpu.ALU.u_wallace._3865_ ),
    .Y(\u_cpu.ALU.u_wallace._4492_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5395_  (.A(\u_cpu.ALU.u_wallace._4492_ ),
    .B(\u_cpu.ALU.u_wallace._4483_ ),
    .Y(\u_cpu.ALU.u_wallace._4493_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._5396_  (.A(\u_cpu.ALU.u_wallace._4357_ ),
    .B(\u_cpu.ALU.u_wallace._4368_ ),
    .X(\u_cpu.ALU.u_wallace._4494_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._5397_  (.A(\u_cpu.ALU.u_wallace._4494_ ),
    .Y(\u_cpu.ALU.u_wallace._4495_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5398_  (.A1(\u_cpu.ALU.u_wallace._4483_ ),
    .A2(\u_cpu.ALU.u_wallace._4492_ ),
    .B1(\u_cpu.ALU.u_wallace._4490_ ),
    .Y(\u_cpu.ALU.u_wallace._4496_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5399_  (.A1_N(\u_cpu.ALU.u_wallace._4491_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4493_ ),
    .B1(\u_cpu.ALU.u_wallace._4495_ ),
    .B2(\u_cpu.ALU.u_wallace._4496_ ),
    .Y(\u_cpu.ALU.u_wallace._4497_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._5400_  (.A1(\u_cpu.ALU.u_wallace._4497_ ),
    .A2(\u_cpu.ALU.u_wallace._4280_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4051_ ),
    .Y(\u_cpu.ALU.u_wallace._4498_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5401_  (.A1(\u_cpu.ALU.u_wallace._4280_ ),
    .A2(\u_cpu.ALU.u_wallace._4497_ ),
    .B1(\u_cpu.ALU.u_wallace._4498_ ),
    .Y(\u_cpu.ALU.u_wallace._4499_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._5402_  (.A1(\u_cpu.ALU.u_wallace._4483_ ),
    .A2(\u_cpu.ALU.u_wallace._4492_ ),
    .B1(\u_cpu.ALU.u_wallace._4494_ ),
    .C1(\u_cpu.ALU.u_wallace._4490_ ),
    .X(\u_cpu.ALU.u_wallace._4500_ ));
 sky130_fd_sc_hd__a21bo_2 \u_cpu.ALU.u_wallace._5403_  (.A1(\u_cpu.ALU.u_wallace._4095_ ),
    .A2(\u_cpu.ALU.u_wallace._3985_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3952_ ),
    .X(\u_cpu.ALU.u_wallace._4501_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5404_  (.A1(\u_cpu.ALU.u_wallace._4495_ ),
    .A2(\u_cpu.ALU.u_wallace._4496_ ),
    .B1(\u_cpu.ALU.u_wallace._4500_ ),
    .C1(\u_cpu.ALU.u_wallace._4501_ ),
    .Y(\u_cpu.ALU.u_wallace._4502_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.ALU.u_wallace._5405_  (.A1(\u_cpu.ALU.u_wallace._4357_ ),
    .A2(\u_cpu.ALU.u_wallace._4368_ ),
    .B1(\u_cpu.ALU.u_wallace._4483_ ),
    .B2(\u_cpu.ALU.u_wallace._4492_ ),
    .C1(\u_cpu.ALU.u_wallace._4490_ ),
    .Y(\u_cpu.ALU.u_wallace._4503_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5406_  (.A1(\u_cpu.ALU.u_wallace._4483_ ),
    .A2(\u_cpu.ALU.u_wallace._4487_ ),
    .B1(\u_cpu.ALU.u_wallace._4489_ ),
    .X(\u_cpu.ALU.u_wallace._4504_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5407_  (.A1(\u_cpu.ALU.u_wallace._4493_ ),
    .A2(\u_cpu.ALU.u_wallace._4504_ ),
    .B1(\u_cpu.ALU.u_wallace._4495_ ),
    .Y(\u_cpu.ALU.u_wallace._4505_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5408_  (.A1(\u_cpu.ALU.u_wallace._4503_ ),
    .A2(\u_cpu.ALU.u_wallace._4505_ ),
    .B1(\u_cpu.ALU.u_wallace._4280_ ),
    .Y(\u_cpu.ALU.u_wallace._4506_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._5409_  (.A1(\u_cpu.ALU.u_wallace._4062_ ),
    .A2(\u_cpu.ALU.u_wallace._4073_ ),
    .A3(\u_cpu.ALU.u_wallace._2670_ ),
    .B1(\u_cpu.ALU.u_wallace._2703_ ),
    .X(\u_cpu.ALU.u_wallace._4507_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5410_  (.A1_N(\u_cpu.ALU.u_wallace._4502_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4506_ ),
    .B1(\u_cpu.ALU.u_wallace._4040_ ),
    .B2(\u_cpu.ALU.u_wallace._4507_ ),
    .Y(\u_cpu.ALU.u_wallace._4508_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._5411_  (.A1(\u_cpu.ALU.u_wallace._4172_ ),
    .A2(\u_cpu.ALU.u_wallace._3328_ ),
    .B1(\u_cpu.ALU.u_wallace._4128_ ),
    .C1(\u_cpu.ALU.u_wallace._4499_ ),
    .D1(\u_cpu.ALU.u_wallace._4508_ ),
    .Y(\u_cpu.ALU.u_wallace._4509_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5412_  (.A(\u_cpu.ALU.u_wallace._4139_ ),
    .B(\u_cpu.ALU.u_wallace._3251_ ),
    .Y(\u_cpu.ALU.u_wallace._4510_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5413_  (.A1(\u_cpu.ALU.u_wallace._4128_ ),
    .A2(\u_cpu.ALU.u_wallace._4510_ ),
    .B1(\u_cpu.ALU.u_wallace._4499_ ),
    .B2(\u_cpu.ALU.u_wallace._4508_ ),
    .X(\u_cpu.ALU.u_wallace._4511_ ));
 sky130_fd_sc_hd__or4_2 \u_cpu.ALU.u_wallace._5414_  (.A(\u_cpu.ALU.u_wallace._3262_ ),
    .B(\u_cpu.ALU.u_wallace._3295_ ),
    .C(\u_cpu.ALU.u_wallace._4161_ ),
    .D(\u_cpu.ALU.u_wallace._4172_ ),
    .X(\u_cpu.ALU.u_wallace._4512_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5415_  (.A1(\u_cpu.ALU.u_wallace._4509_ ),
    .A2(\u_cpu.ALU.u_wallace._4511_ ),
    .B1(\u_cpu.ALU.u_wallace._4512_ ),
    .Y(\u_cpu.ALU.u_wallace._4513_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5416_  (.A(\u_cpu.ALU.u_wallace._4512_ ),
    .B(\u_cpu.ALU.u_wallace._4509_ ),
    .C(\u_cpu.ALU.u_wallace._4511_ ),
    .Y(\u_cpu.ALU.u_wallace._4514_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.ALU.u_wallace._5417_  (.A_N(\u_cpu.ALU.u_wallace._4513_ ),
    .B(\u_cpu.ALU.u_wallace._4514_ ),
    .X(\u_cpu.ALU.u_wallace._4515_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._5418_  (.A(\u_cpu.ALU.u_wallace._4269_ ),
    .B(\u_cpu.ALU.u_wallace._4515_ ),
    .X(\u_cpu.ALU.Product_Wallace[9] ));
 sky130_fd_sc_hd__a32oi_2 \u_cpu.ALU.u_wallace._5419_  (.A1(\u_cpu.ALU.u_wallace._4512_ ),
    .A2(\u_cpu.ALU.u_wallace._4509_ ),
    .A3(\u_cpu.ALU.u_wallace._4511_ ),
    .B1(\u_cpu.ALU.u_wallace._4258_ ),
    .B2(\u_cpu.ALU.u_wallace._4226_ ),
    .Y(\u_cpu.ALU.u_wallace._4516_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5420_  (.A(\u_cpu.ALU.u_wallace._4513_ ),
    .B(\u_cpu.ALU.u_wallace._4516_ ),
    .Y(\u_cpu.ALU.u_wallace._4517_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5421_  (.A1(\u_cpu.ALU.u_wallace._4502_ ),
    .A2(\u_cpu.ALU.u_wallace._4506_ ),
    .B1(\u_cpu.ALU.u_wallace._4051_ ),
    .Y(\u_cpu.ALU.u_wallace._4518_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._5422_  (.A1(\u_cpu.ALU.u_wallace._4502_ ),
    .A2(\u_cpu.ALU.u_wallace._4498_ ),
    .B1(\u_cpu.ALU.u_wallace._4510_ ),
    .C1(\u_cpu.ALU.u_wallace._4518_ ),
    .X(\u_cpu.ALU.u_wallace._4519_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5423_  (.A(\u_cpu.ALU.u_wallace._4128_ ),
    .B(\u_cpu.ALU.u_wallace._4518_ ),
    .Y(\u_cpu.ALU.u_wallace._4520_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU.u_wallace._5424_  (.A1(\u_cpu.ALU.u_wallace._3569_ ),
    .A2(\u_cpu.ALU.u_wallace._3930_ ),
    .B1(\u_cpu.ALU.u_wallace._4324_ ),
    .C1(\u_cpu.ALU.u_wallace._4335_ ),
    .Y(\u_cpu.ALU.u_wallace._4521_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5425_  (.A1(\u_cpu.ALU.u_wallace._4324_ ),
    .A2(\u_cpu.ALU.u_wallace._4335_ ),
    .B1(\u_cpu.ALU.u_wallace._3569_ ),
    .C1(\u_cpu.ALU.u_wallace._3930_ ),
    .X(\u_cpu.ALU.u_wallace._4522_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5426_  (.A1_N(\u_cpu.ALU.u_wallace._4493_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4504_ ),
    .B1(\u_cpu.ALU.u_wallace._4521_ ),
    .B2(\u_cpu.ALU.u_wallace._4522_ ),
    .Y(\u_cpu.ALU.u_wallace._4523_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5427_  (.A(\u_cpu.ALU.u_wallace._4501_ ),
    .B(\u_cpu.ALU.u_wallace._4500_ ),
    .C(\u_cpu.ALU.u_wallace._4523_ ),
    .X(\u_cpu.ALU.u_wallace._4524_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5428_  (.A1(\u_cpu.ALU.u_wallace._4051_ ),
    .A2(\u_cpu.ALU.u_wallace._4506_ ),
    .B1(\u_cpu.ALU.u_wallace._4524_ ),
    .Y(\u_cpu.ALU.u_wallace._4525_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5429_  (.A(\u_cpu.ALU.u_wallace._4489_ ),
    .B(\u_cpu.ALU.u_wallace._4483_ ),
    .C(\u_cpu.ALU.u_wallace._4487_ ),
    .X(\u_cpu.ALU.u_wallace._4526_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5430_  (.A(\u_cpu.ALU.u_wallace._0600_ ),
    .X(\u_cpu.ALU.u_wallace._4527_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5431_  (.A1(\u_cpu.ALU.u_wallace._3832_ ),
    .A2(\u_cpu.ALU.u_wallace._2045_ ),
    .B1(\u_cpu.ALU.u_wallace._1552_ ),
    .B2(\u_cpu.ALU.u_wallace._1125_ ),
    .X(\u_cpu.ALU.u_wallace._4528_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5432_  (.A(\u_cpu.ALU.u_wallace._1114_ ),
    .X(\u_cpu.ALU.u_wallace._4529_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5433_  (.A(\u_cpu.ALU.u_wallace._1848_ ),
    .B(\u_cpu.ALU.u_wallace._4529_ ),
    .C(\u_cpu.ALU.u_wallace._1530_ ),
    .D(\u_cpu.ALU.u_wallace._1552_ ),
    .Y(\u_cpu.ALU.u_wallace._4530_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5434_  (.A1(\u_cpu.ALU.u_wallace._4527_ ),
    .A2(\u_cpu.ALU.u_wallace._2604_ ),
    .B1(\u_cpu.ALU.u_wallace._4528_ ),
    .B2(\u_cpu.ALU.u_wallace._4530_ ),
    .Y(\u_cpu.ALU.u_wallace._4531_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5435_  (.A1(\u_cpu.ALU.u_wallace._3777_ ),
    .A2(\u_cpu.ALU.u_wallace._2045_ ),
    .B1(\u_cpu.ALU.u_wallace._2056_ ),
    .B2(\u_cpu.ALU.u_wallace._1125_ ),
    .Y(\u_cpu.ALU.u_wallace._4532_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5436_  (.A(\u_cpu.ALU.u_wallace._1421_ ),
    .B(\u_cpu.ALU.u_wallace._3404_ ),
    .Y(\u_cpu.ALU.u_wallace._4533_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5437_  (.A(\u_cpu.ALU.u_wallace._3777_ ),
    .B(\u_cpu.ALU.u_wallace._1979_ ),
    .C(\u_cpu.ALU.u_wallace._2571_ ),
    .D(\u_cpu.ALU.u_wallace._2078_ ),
    .X(\u_cpu.ALU.u_wallace._4534_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._5438_  (.A(\u_cpu.ALU.u_wallace._4532_ ),
    .B(\u_cpu.ALU.u_wallace._4533_ ),
    .C(\u_cpu.ALU.u_wallace._4534_ ),
    .Y(\u_cpu.ALU.u_wallace._4535_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5439_  (.A(\u_cpu.ALU.u_wallace._1848_ ),
    .B(\u_cpu.ALU.u_wallace._0753_ ),
    .Y(\u_cpu.ALU.u_wallace._4536_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5440_  (.A1(\u_cpu.ALU.u_wallace._4536_ ),
    .A2(\u_cpu.ALU.u_wallace._4448_ ),
    .B1(\u_cpu.ALU.u_wallace._4451_ ),
    .Y(\u_cpu.ALU.u_wallace._4537_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._5441_  (.A1(\u_cpu.ALU.u_wallace._4531_ ),
    .A2(\u_cpu.ALU.u_wallace._4535_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4537_ ),
    .Y(\u_cpu.ALU.u_wallace._4538_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5442_  (.A(\u_cpu.ALU.u_wallace._4470_ ),
    .X(\u_cpu.ALU.u_wallace._4539_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5443_  (.A1(\u_cpu.ALU.u_wallace._0621_ ),
    .A2(\u_cpu.ALU.u_wallace._4539_ ),
    .B1(\u_cpu.ALU.u_wallace._4532_ ),
    .B2(\u_cpu.ALU.u_wallace._4534_ ),
    .Y(\u_cpu.ALU.u_wallace._4540_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5444_  (.A(\u_cpu.ALU.u_wallace._1421_ ),
    .X(\u_cpu.ALU.u_wallace._4541_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5445_  (.A(\u_cpu.ALU.u_wallace._3404_ ),
    .X(\u_cpu.ALU.u_wallace._4542_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5446_  (.A(\u_cpu.ALU.u_wallace._4528_ ),
    .B(\u_cpu.ALU.u_wallace._4530_ ),
    .C(\u_cpu.ALU.u_wallace._4541_ ),
    .D(\u_cpu.ALU.u_wallace._4542_ ),
    .Y(\u_cpu.ALU.u_wallace._4543_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5447_  (.A(\u_cpu.ALU.u_wallace._4537_ ),
    .B(\u_cpu.ALU.u_wallace._4540_ ),
    .C(\u_cpu.ALU.u_wallace._4543_ ),
    .Y(\u_cpu.ALU.u_wallace._4544_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5448_  (.A(\u_cpu.ALU.u_wallace._0512_ ),
    .X(\u_cpu.ALU.u_wallace._4545_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._5449_  (.A1(\u_cpu.ALU.u_wallace._4475_ ),
    .A2(\u_cpu.ALU.u_wallace._4542_ ),
    .A3(\u_cpu.ALU.u_wallace._4545_ ),
    .B1(\u_cpu.ALU.u_wallace._4472_ ),
    .X(\u_cpu.ALU.u_wallace._4546_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5450_  (.A1(\u_cpu.ALU.u_wallace._4538_ ),
    .A2(\u_cpu.ALU.u_wallace._4544_ ),
    .B1(\u_cpu.ALU.u_wallace._4546_ ),
    .X(\u_cpu.ALU.u_wallace._4547_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5451_  (.A(\u_cpu.ALU.u_wallace._4537_ ),
    .B(\u_cpu.ALU.u_wallace._4540_ ),
    .Y(\u_cpu.ALU.u_wallace._4548_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5452_  (.A1(\u_cpu.ALU.u_wallace._4535_ ),
    .A2(\u_cpu.ALU.u_wallace._4548_ ),
    .B1(\u_cpu.ALU.u_wallace._4538_ ),
    .C1(\u_cpu.ALU.u_wallace._4546_ ),
    .Y(\u_cpu.ALU.u_wallace._4549_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5453_  (.A(\u_cpu.ALU.SrcA[10] ),
    .X(\u_cpu.ALU.u_wallace._4550_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5454_  (.A(\u_cpu.ALU.u_wallace._4550_ ),
    .X(\u_cpu.ALU.u_wallace._4551_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5455_  (.A1(\u_cpu.ALU.u_wallace._1771_ ),
    .A2(\u_cpu.ALU.u_wallace._2922_ ),
    .B1(\u_cpu.ALU.u_wallace._4551_ ),
    .B2(\u_cpu.ALU.u_wallace._1749_ ),
    .Y(\u_cpu.ALU.u_wallace._4552_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5456_  (.A(\u_cpu.ALU.SrcA[10] ),
    .X(\u_cpu.ALU.u_wallace._4553_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5457_  (.A(\u_cpu.ALU.u_wallace._4553_ ),
    .X(\u_cpu.ALU.u_wallace._4554_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._5458_  (.A1(\u_cpu.ALU.u_wallace._2757_ ),
    .A2(\u_cpu.ALU.u_wallace._2779_ ),
    .A3(\u_cpu.ALU.u_wallace._0906_ ),
    .A4(\u_cpu.ALU.u_wallace._4554_ ),
    .B1(\u_cpu.ALU.u_wallace._4442_ ),
    .X(\u_cpu.ALU.u_wallace._4555_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5459_  (.A(\u_cpu.ALU.SrcA[4] ),
    .X(\u_cpu.ALU.u_wallace._4556_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5460_  (.A(\u_cpu.ALU.SrcA[10] ),
    .X(\u_cpu.ALU.u_wallace._4557_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5461_  (.A(\u_cpu.ALU.u_wallace._2747_ ),
    .B(\u_cpu.ALU.u_wallace._2856_ ),
    .C(\u_cpu.ALU.u_wallace._4556_ ),
    .D(\u_cpu.ALU.u_wallace._4557_ ),
    .X(\u_cpu.ALU.u_wallace._4558_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5462_  (.A1(\u_cpu.ALU.u_wallace._4552_ ),
    .A2(\u_cpu.ALU.u_wallace._4558_ ),
    .B1(\u_cpu.ALU.u_wallace._4442_ ),
    .Y(\u_cpu.ALU.u_wallace._4559_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5463_  (.A1(\u_cpu.ALU.u_wallace._3623_ ),
    .A2(\u_cpu.ALU.u_wallace._1968_ ),
    .B1(\u_cpu.ALU.u_wallace._4439_ ),
    .B2(\u_cpu.ALU.u_wallace._1957_ ),
    .Y(\u_cpu.ALU.u_wallace._4560_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5464_  (.A(\u_cpu.ALU.SrcA[8] ),
    .X(\u_cpu.ALU.u_wallace._4561_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5465_  (.A(\u_cpu.ALU.u_wallace._4401_ ),
    .X(\u_cpu.ALU.u_wallace._4562_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5466_  (.A(\u_cpu.ALU.u_wallace._4561_ ),
    .B(\u_cpu.ALU.u_wallace._0206_ ),
    .C(\u_cpu.ALU.u_wallace._0490_ ),
    .D(\u_cpu.ALU.u_wallace._4562_ ),
    .X(\u_cpu.ALU.u_wallace._4563_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5467_  (.A(\u_cpu.ALU.u_wallace._3821_ ),
    .B(\u_cpu.ALU.u_wallace._0753_ ),
    .Y(\u_cpu.ALU.u_wallace._4564_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5468_  (.A1(\u_cpu.ALU.u_wallace._4560_ ),
    .A2(\u_cpu.ALU.u_wallace._4563_ ),
    .B1(\u_cpu.ALU.u_wallace._4564_ ),
    .Y(\u_cpu.ALU.u_wallace._4565_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5469_  (.A1(\u_cpu.ALU.u_wallace._3623_ ),
    .A2(\u_cpu.ALU.u_wallace._1968_ ),
    .B1(\u_cpu.ALU.u_wallace._4439_ ),
    .B2(\u_cpu.ALU.u_wallace._1957_ ),
    .X(\u_cpu.ALU.u_wallace._4566_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5470_  (.A(\u_cpu.ALU.u_wallace._4401_ ),
    .X(\u_cpu.ALU.u_wallace._4567_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5471_  (.A(\u_cpu.ALU.u_wallace._4449_ ),
    .B(\u_cpu.ALU.u_wallace._0523_ ),
    .C(\u_cpu.ALU.u_wallace._1169_ ),
    .D(\u_cpu.ALU.u_wallace._4567_ ),
    .Y(\u_cpu.ALU.u_wallace._4568_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5472_  (.A(\u_cpu.ALU.u_wallace._4566_ ),
    .B(\u_cpu.ALU.u_wallace._4568_ ),
    .C(\u_cpu.ALU.u_wallace._2801_ ),
    .D(\u_cpu.ALU.u_wallace._0578_ ),
    .Y(\u_cpu.ALU.u_wallace._4569_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._5473_  (.A1(\u_cpu.ALU.u_wallace._4552_ ),
    .A2(\u_cpu.ALU.u_wallace._4555_ ),
    .B1(\u_cpu.ALU.u_wallace._4559_ ),
    .C1(\u_cpu.ALU.u_wallace._4565_ ),
    .D1(\u_cpu.ALU.u_wallace._4569_ ),
    .X(\u_cpu.ALU.u_wallace._4570_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5474_  (.A1(\u_cpu.ALU.u_wallace._2779_ ),
    .A2(\u_cpu.ALU.u_wallace._1180_ ),
    .B1(\u_cpu.ALU.u_wallace._4554_ ),
    .B2(\u_cpu.ALU.u_wallace._0873_ ),
    .X(\u_cpu.ALU.u_wallace._4571_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5475_  (.A(\u_cpu.ALU.u_wallace._2757_ ),
    .B(\u_cpu.ALU.u_wallace._2779_ ),
    .C(\u_cpu.ALU.u_wallace._0906_ ),
    .D(\u_cpu.ALU.u_wallace._4554_ ),
    .Y(\u_cpu.ALU.u_wallace._4572_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._5476_  (.A(\u_cpu.ALU.u_wallace._4401_ ),
    .Y(\u_cpu.ALU.u_wallace._4573_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5477_  (.A(\u_cpu.ALU.u_wallace._4923_ ),
    .B(\u_cpu.ALU.u_wallace._4573_ ),
    .Y(\u_cpu.ALU.u_wallace._4574_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._5478_  (.A(\u_cpu.ALU.u_wallace._2779_ ),
    .B(\u_cpu.ALU.u_wallace._1191_ ),
    .X(\u_cpu.ALU.u_wallace._4575_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5479_  (.A(\u_cpu.ALU.u_wallace._4571_ ),
    .B(\u_cpu.ALU.u_wallace._4572_ ),
    .C(\u_cpu.ALU.u_wallace._4574_ ),
    .D(\u_cpu.ALU.u_wallace._4575_ ),
    .Y(\u_cpu.ALU.u_wallace._4576_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5480_  (.A1(\u_cpu.ALU.u_wallace._4565_ ),
    .A2(\u_cpu.ALU.u_wallace._4569_ ),
    .B1(\u_cpu.ALU.u_wallace._4559_ ),
    .B2(\u_cpu.ALU.u_wallace._4576_ ),
    .Y(\u_cpu.ALU.u_wallace._4577_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._5481_  (.A(\u_cpu.ALU.u_wallace._3711_ ),
    .B(\u_cpu.ALU.u_wallace._4423_ ),
    .C(\u_cpu.ALU.u_wallace._4445_ ),
    .Y(\u_cpu.ALU.u_wallace._4578_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._5482_  (.A1(\u_cpu.ALU.u_wallace._4446_ ),
    .A2(\u_cpu.ALU.u_wallace._4453_ ),
    .A3(\u_cpu.ALU.u_wallace._4456_ ),
    .B1(\u_cpu.ALU.u_wallace._4578_ ),
    .X(\u_cpu.ALU.u_wallace._4579_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._5483_  (.A1(\u_cpu.ALU.u_wallace._4570_ ),
    .A2(\u_cpu.ALU.u_wallace._4577_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4579_ ),
    .Y(\u_cpu.ALU.u_wallace._4580_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._5484_  (.A1(\u_cpu.ALU.u_wallace._4552_ ),
    .A2(\u_cpu.ALU.u_wallace._4555_ ),
    .B1(\u_cpu.ALU.u_wallace._4559_ ),
    .C1(\u_cpu.ALU.u_wallace._4565_ ),
    .D1(\u_cpu.ALU.u_wallace._4569_ ),
    .Y(\u_cpu.ALU.u_wallace._4581_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5485_  (.A1(\u_cpu.ALU.u_wallace._4565_ ),
    .A2(\u_cpu.ALU.u_wallace._4569_ ),
    .B1(\u_cpu.ALU.u_wallace._4559_ ),
    .B2(\u_cpu.ALU.u_wallace._4576_ ),
    .X(\u_cpu.ALU.u_wallace._4582_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5486_  (.A(\u_cpu.ALU.u_wallace._4581_ ),
    .B(\u_cpu.ALU.u_wallace._4582_ ),
    .C(\u_cpu.ALU.u_wallace._4579_ ),
    .Y(\u_cpu.ALU.u_wallace._4583_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5487_  (.A1(\u_cpu.ALU.u_wallace._4547_ ),
    .A2(\u_cpu.ALU.u_wallace._4549_ ),
    .B1(\u_cpu.ALU.u_wallace._4580_ ),
    .B2(\u_cpu.ALU.u_wallace._4583_ ),
    .Y(\u_cpu.ALU.u_wallace._4584_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5488_  (.A1(\u_cpu.ALU.u_wallace._4570_ ),
    .A2(\u_cpu.ALU.u_wallace._4577_ ),
    .B1(\u_cpu.ALU.u_wallace._4443_ ),
    .C1(\u_cpu.ALU.u_wallace._4458_ ),
    .X(\u_cpu.ALU.u_wallace._4585_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5489_  (.A(\u_cpu.ALU.u_wallace._4537_ ),
    .B(\u_cpu.ALU.u_wallace._4540_ ),
    .C(\u_cpu.ALU.u_wallace._4543_ ),
    .X(\u_cpu.ALU.u_wallace._4586_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5490_  (.A(\u_cpu.ALU.u_wallace._4546_ ),
    .B(\u_cpu.ALU.u_wallace._4538_ ),
    .Y(\u_cpu.ALU.u_wallace._4587_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5491_  (.A1(\u_cpu.ALU.u_wallace._4586_ ),
    .A2(\u_cpu.ALU.u_wallace._4587_ ),
    .B1(\u_cpu.ALU.u_wallace._4583_ ),
    .C1(\u_cpu.ALU.u_wallace._4547_ ),
    .Y(\u_cpu.ALU.u_wallace._4588_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5492_  (.A(\u_cpu.ALU.u_wallace._4390_ ),
    .B(\u_cpu.ALU.u_wallace._4458_ ),
    .Y(\u_cpu.ALU.u_wallace._4589_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5493_  (.A1_N(\u_cpu.ALU.u_wallace._4462_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4486_ ),
    .B1(\u_cpu.ALU.u_wallace._4460_ ),
    .B2(\u_cpu.ALU.u_wallace._4589_ ),
    .Y(\u_cpu.ALU.u_wallace._4590_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5494_  (.A1(\u_cpu.ALU.u_wallace._4585_ ),
    .A2(\u_cpu.ALU.u_wallace._4588_ ),
    .B1(\u_cpu.ALU.u_wallace._4590_ ),
    .Y(\u_cpu.ALU.u_wallace._4591_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._5495_  (.A1(\u_cpu.ALU.u_wallace._4587_ ),
    .A2(\u_cpu.ALU.u_wallace._4586_ ),
    .B1(\u_cpu.ALU.u_wallace._4547_ ),
    .C1(\u_cpu.ALU.u_wallace._4580_ ),
    .D1(\u_cpu.ALU.u_wallace._4583_ ),
    .X(\u_cpu.ALU.u_wallace._4592_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._5496_  (.A1(\u_cpu.ALU.u_wallace._4584_ ),
    .A2(\u_cpu.ALU.u_wallace._4592_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4590_ ),
    .Y(\u_cpu.ALU.u_wallace._4593_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5497_  (.A(\u_cpu.ALU.SrcB[8] ),
    .X(\u_cpu.ALU.u_wallace._4594_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5498_  (.A(\u_cpu.ALU.SrcB[9] ),
    .X(\u_cpu.ALU.u_wallace._4595_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5499_  (.A1(\u_cpu.ALU.u_wallace._0512_ ),
    .A2(\u_cpu.ALU.u_wallace._4594_ ),
    .B1(\u_cpu.ALU.u_wallace._4595_ ),
    .B2(\u_cpu.ALU.u_wallace._0250_ ),
    .X(\u_cpu.ALU.u_wallace._4596_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5500_  (.A(\u_cpu.ALU.u_wallace._0392_ ),
    .X(\u_cpu.ALU.u_wallace._4597_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5501_  (.A(\u_cpu.ALU.SrcB[9] ),
    .X(\u_cpu.ALU.u_wallace._4598_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5502_  (.A(\u_cpu.ALU.u_wallace._4598_ ),
    .X(\u_cpu.ALU.u_wallace._4599_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5503_  (.A(\u_cpu.ALU.u_wallace._4597_ ),
    .B(\u_cpu.ALU.u_wallace._0151_ ),
    .C(\u_cpu.ALU.u_wallace._4018_ ),
    .D(\u_cpu.ALU.u_wallace._4599_ ),
    .Y(\u_cpu.ALU.u_wallace._4600_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._5504_  (.A(\u_cpu.ALU.SrcB[10] ),
    .Y(\u_cpu.ALU.u_wallace._4601_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5505_  (.A(\u_cpu.ALU.u_wallace._4601_ ),
    .X(\u_cpu.ALU.u_wallace._4602_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU.u_wallace._5506_  (.A1_N(\u_cpu.ALU.u_wallace._4596_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4600_ ),
    .B1(\u_cpu.ALU.u_wallace._0032_ ),
    .B2(\u_cpu.ALU.u_wallace._4602_ ),
    .X(\u_cpu.ALU.u_wallace._4603_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5507_  (.A(\u_cpu.ALU.SrcB[10] ),
    .X(\u_cpu.ALU.u_wallace._4604_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5508_  (.A(\u_cpu.ALU.u_wallace._4604_ ),
    .X(\u_cpu.ALU.u_wallace._4605_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5509_  (.A(\u_cpu.ALU.u_wallace._4596_ ),
    .B(\u_cpu.ALU.u_wallace._4600_ ),
    .C(\u_cpu.ALU.u_wallace._1070_ ),
    .D(\u_cpu.ALU.u_wallace._4605_ ),
    .X(\u_cpu.ALU.u_wallace._4606_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5510_  (.A(\u_cpu.ALU.u_wallace._0108_ ),
    .B(\u_cpu.ALU.u_wallace._0162_ ),
    .C(\u_cpu.ALU.u_wallace._4029_ ),
    .D(\u_cpu.ALU.u_wallace._4313_ ),
    .Y(\u_cpu.ALU.u_wallace._4607_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5511_  (.A1(\u_cpu.ALU.u_wallace._4603_ ),
    .A2(\u_cpu.ALU.u_wallace._4606_ ),
    .B1(\u_cpu.ALU.u_wallace._4607_ ),
    .Y(\u_cpu.ALU.u_wallace._4608_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5512_  (.A(\u_cpu.ALU.SrcB[10] ),
    .X(\u_cpu.ALU.u_wallace._4609_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5513_  (.A(\u_cpu.ALU.u_wallace._4609_ ),
    .X(\u_cpu.ALU.u_wallace._4610_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5514_  (.A(\u_cpu.ALU.u_wallace._4600_ ),
    .B(\u_cpu.ALU.u_wallace._4610_ ),
    .C(\u_cpu.ALU.u_wallace._0994_ ),
    .X(\u_cpu.ALU.u_wallace._4611_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._5515_  (.A1(\u_cpu.ALU.u_wallace._4611_ ),
    .A2(\u_cpu.ALU.u_wallace._4596_ ),
    .B1(\u_cpu.ALU.u_wallace._4607_ ),
    .C1(\u_cpu.ALU.u_wallace._4603_ ),
    .X(\u_cpu.ALU.u_wallace._4612_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5516_  (.A1(\u_cpu.ALU.u_wallace._4479_ ),
    .A2(\u_cpu.ALU.u_wallace._4478_ ),
    .B1(\u_cpu.ALU.u_wallace._4608_ ),
    .C1(\u_cpu.ALU.u_wallace._4612_ ),
    .X(\u_cpu.ALU.u_wallace._4613_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5517_  (.A1(\u_cpu.ALU.u_wallace._3360_ ),
    .A2(\u_cpu.ALU.u_wallace._4464_ ),
    .B1(\u_cpu.ALU.u_wallace._4474_ ),
    .C1(\u_cpu.ALU.u_wallace._4477_ ),
    .Y(\u_cpu.ALU.u_wallace._4614_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5518_  (.A(\u_cpu.ALU.u_wallace._4608_ ),
    .B(\u_cpu.ALU.u_wallace._4612_ ),
    .Y(\u_cpu.ALU.u_wallace._4615_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5519_  (.A(\u_cpu.ALU.u_wallace._4474_ ),
    .B(\u_cpu.ALU.u_wallace._4614_ ),
    .C(\u_cpu.ALU.u_wallace._4615_ ),
    .X(\u_cpu.ALU.u_wallace._4616_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5520_  (.A(\u_cpu.ALU.u_wallace._4613_ ),
    .B(\u_cpu.ALU.u_wallace._4616_ ),
    .Y(\u_cpu.ALU.u_wallace._4617_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5521_  (.A1(\u_cpu.ALU.u_wallace._4584_ ),
    .A2(\u_cpu.ALU.u_wallace._4591_ ),
    .B1(\u_cpu.ALU.u_wallace._4593_ ),
    .C1(\u_cpu.ALU.u_wallace._4617_ ),
    .Y(\u_cpu.ALU.u_wallace._4618_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5522_  (.A1(\u_cpu.ALU.u_wallace._4547_ ),
    .A2(\u_cpu.ALU.u_wallace._4549_ ),
    .B1(\u_cpu.ALU.u_wallace._4580_ ),
    .B2(\u_cpu.ALU.u_wallace._4583_ ),
    .X(\u_cpu.ALU.u_wallace._4619_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5523_  (.A1(\u_cpu.ALU.u_wallace._4585_ ),
    .A2(\u_cpu.ALU.u_wallace._4588_ ),
    .B1(\u_cpu.ALU.u_wallace._4619_ ),
    .C1(\u_cpu.ALU.u_wallace._4590_ ),
    .Y(\u_cpu.ALU.u_wallace._4620_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5524_  (.A1_N(\u_cpu.ALU.u_wallace._4620_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4593_ ),
    .B1(\u_cpu.ALU.u_wallace._4613_ ),
    .B2(\u_cpu.ALU.u_wallace._4616_ ),
    .Y(\u_cpu.ALU.u_wallace._4621_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5525_  (.A1(\u_cpu.ALU.u_wallace._4526_ ),
    .A2(\u_cpu.ALU.u_wallace._4491_ ),
    .B1(\u_cpu.ALU.u_wallace._4618_ ),
    .C1(\u_cpu.ALU.u_wallace._4621_ ),
    .X(\u_cpu.ALU.u_wallace._4622_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5526_  (.A1(\u_cpu.ALU.u_wallace._4494_ ),
    .A2(\u_cpu.ALU.u_wallace._4490_ ),
    .B1(\u_cpu.ALU.u_wallace._4493_ ),
    .Y(\u_cpu.ALU.u_wallace._4623_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5527_  (.A1(\u_cpu.ALU.u_wallace._4618_ ),
    .A2(\u_cpu.ALU.u_wallace._4621_ ),
    .B1(\u_cpu.ALU.u_wallace._4623_ ),
    .Y(\u_cpu.ALU.u_wallace._4624_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5528_  (.A1(\u_cpu.ALU.u_wallace._4622_ ),
    .A2(\u_cpu.ALU.u_wallace._4624_ ),
    .B1(\u_cpu.ALU.u_wallace._4521_ ),
    .Y(\u_cpu.ALU.u_wallace._4625_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._5529_  (.A1(\u_cpu.ALU.u_wallace._3569_ ),
    .A2(\u_cpu.ALU.u_wallace._3930_ ),
    .B1(\u_cpu.ALU.u_wallace._4324_ ),
    .C1(\u_cpu.ALU.u_wallace._4335_ ),
    .X(\u_cpu.ALU.u_wallace._4626_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5530_  (.A1(\u_cpu.ALU.u_wallace._4526_ ),
    .A2(\u_cpu.ALU.u_wallace._4491_ ),
    .B1(\u_cpu.ALU.u_wallace._4618_ ),
    .C1(\u_cpu.ALU.u_wallace._4621_ ),
    .Y(\u_cpu.ALU.u_wallace._4627_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5531_  (.A1(\u_cpu.ALU.u_wallace._4618_ ),
    .A2(\u_cpu.ALU.u_wallace._4621_ ),
    .B1(\u_cpu.ALU.u_wallace._4623_ ),
    .X(\u_cpu.ALU.u_wallace._4628_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5532_  (.A(\u_cpu.ALU.u_wallace._4626_ ),
    .B(\u_cpu.ALU.u_wallace._4627_ ),
    .C(\u_cpu.ALU.u_wallace._4628_ ),
    .Y(\u_cpu.ALU.u_wallace._4629_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5533_  (.A(\u_cpu.ALU.u_wallace._4525_ ),
    .B(\u_cpu.ALU.u_wallace._4625_ ),
    .C(\u_cpu.ALU.u_wallace._4629_ ),
    .Y(\u_cpu.ALU.u_wallace._4630_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5534_  (.A(\u_cpu.ALU.u_wallace._4628_ ),
    .B(\u_cpu.ALU.u_wallace._4521_ ),
    .Y(\u_cpu.ALU.u_wallace._4631_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5535_  (.A1(\u_cpu.ALU.u_wallace._4622_ ),
    .A2(\u_cpu.ALU.u_wallace._4624_ ),
    .B1(\u_cpu.ALU.u_wallace._4626_ ),
    .Y(\u_cpu.ALU.u_wallace._4632_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._5536_  (.A1(\u_cpu.ALU.u_wallace._4524_ ),
    .A2(\u_cpu.ALU.u_wallace._4498_ ),
    .B1(\u_cpu.ALU.u_wallace._4622_ ),
    .B2(\u_cpu.ALU.u_wallace._4631_ ),
    .C1(\u_cpu.ALU.u_wallace._4632_ ),
    .Y(\u_cpu.ALU.u_wallace._4633_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5537_  (.A1(\u_cpu.ALU.u_wallace._4520_ ),
    .A2(\u_cpu.ALU.u_wallace._4499_ ),
    .B1(\u_cpu.ALU.u_wallace._4630_ ),
    .B2(\u_cpu.ALU.u_wallace._4633_ ),
    .Y(\u_cpu.ALU.u_wallace._4634_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5538_  (.A(\u_cpu.ALU.u_wallace._4520_ ),
    .B(\u_cpu.ALU.u_wallace._4630_ ),
    .C(\u_cpu.ALU.u_wallace._4499_ ),
    .X(\u_cpu.ALU.u_wallace._4635_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5539_  (.A(\u_cpu.ALU.u_wallace._4634_ ),
    .B(\u_cpu.ALU.u_wallace._4635_ ),
    .Y(\u_cpu.ALU.u_wallace._4636_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._5540_  (.A(\u_cpu.ALU.u_wallace._4519_ ),
    .B(\u_cpu.ALU.u_wallace._4636_ ),
    .X(\u_cpu.ALU.u_wallace._4637_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._5541_  (.A(\u_cpu.ALU.u_wallace._4517_ ),
    .B(\u_cpu.ALU.u_wallace._4637_ ),
    .X(\u_cpu.ALU.Product_Wallace[10] ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5542_  (.A(\u_cpu.ALU.u_wallace._4630_ ),
    .B(\u_cpu.ALU.u_wallace._4633_ ),
    .Y(\u_cpu.ALU.u_wallace._4638_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5543_  (.A(\u_cpu.ALU.u_wallace._4499_ ),
    .B(\u_cpu.ALU.u_wallace._4508_ ),
    .C(\u_cpu.ALU.u_wallace._4161_ ),
    .Y(\u_cpu.ALU.u_wallace._4639_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5544_  (.A1(\u_cpu.ALU.u_wallace._4626_ ),
    .A2(\u_cpu.ALU.u_wallace._4624_ ),
    .B1(\u_cpu.ALU.u_wallace._4627_ ),
    .Y(\u_cpu.ALU.u_wallace._4640_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5545_  (.A1_N(\u_cpu.ALU.u_wallace._4617_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4593_ ),
    .B1(\u_cpu.ALU.u_wallace._4591_ ),
    .B2(\u_cpu.ALU.u_wallace._4584_ ),
    .Y(\u_cpu.ALU.u_wallace._4641_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5546_  (.A(\u_cpu.ALU.SrcA[10] ),
    .X(\u_cpu.ALU.u_wallace._4642_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5547_  (.A(\u_cpu.ALU.u_wallace._4642_ ),
    .X(\u_cpu.ALU.u_wallace._4643_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5548_  (.A(\u_cpu.ALU.u_wallace._2747_ ),
    .B(\u_cpu.ALU.u_wallace._2856_ ),
    .C(\u_cpu.ALU.u_wallace._4556_ ),
    .X(\u_cpu.ALU.u_wallace._4644_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5549_  (.A(\u_cpu.ALU.u_wallace._1760_ ),
    .X(\u_cpu.ALU.u_wallace._4645_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5550_  (.A(\u_cpu.ALU.SrcA[11] ),
    .X(\u_cpu.ALU.u_wallace._4646_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5551_  (.A(\u_cpu.ALU.u_wallace._4646_ ),
    .X(\u_cpu.ALU.u_wallace._4647_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5552_  (.A1(\u_cpu.ALU.u_wallace._4645_ ),
    .A2(\u_cpu.ALU.u_wallace._2955_ ),
    .B1(\u_cpu.ALU.u_wallace._4647_ ),
    .B2(\u_cpu.ALU.u_wallace._0075_ ),
    .Y(\u_cpu.ALU.u_wallace._4648_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5553_  (.A(\u_cpu.ALU.SrcB[6] ),
    .X(\u_cpu.ALU.u_wallace._4649_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5554_  (.A(\u_cpu.ALU.SrcA[11] ),
    .X(\u_cpu.ALU.u_wallace._4650_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5555_  (.A(\u_cpu.ALU.u_wallace._0064_ ),
    .B(\u_cpu.ALU.u_wallace._4649_ ),
    .C(\u_cpu.ALU.u_wallace._1114_ ),
    .D(\u_cpu.ALU.u_wallace._4650_ ),
    .X(\u_cpu.ALU.u_wallace._4651_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5556_  (.A1_N(\u_cpu.ALU.u_wallace._4643_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4644_ ),
    .B1(\u_cpu.ALU.u_wallace._4648_ ),
    .B2(\u_cpu.ALU.u_wallace._4651_ ),
    .Y(\u_cpu.ALU.u_wallace._4652_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5557_  (.A(\u_cpu.ALU.u_wallace._4646_ ),
    .X(\u_cpu.ALU.u_wallace._4653_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5558_  (.A(\u_cpu.ALU.u_wallace._1749_ ),
    .B(\u_cpu.ALU.u_wallace._1771_ ),
    .C(\u_cpu.ALU.u_wallace._1979_ ),
    .D(\u_cpu.ALU.u_wallace._4653_ ),
    .Y(\u_cpu.ALU.u_wallace._4654_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._5559_  (.A_N(\u_cpu.ALU.u_wallace._4648_ ),
    .B(\u_cpu.ALU.u_wallace._4654_ ),
    .C(\u_cpu.ALU.u_wallace._4558_ ),
    .Y(\u_cpu.ALU.u_wallace._4655_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5560_  (.A1(\u_cpu.ALU.u_wallace._0807_ ),
    .A2(\u_cpu.ALU.u_wallace._4401_ ),
    .B1(\u_cpu.ALU.u_wallace._4553_ ),
    .B2(\u_cpu.ALU.u_wallace._1903_ ),
    .Y(\u_cpu.ALU.u_wallace._4656_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5561_  (.A(\u_cpu.ALU.u_wallace._0195_ ),
    .X(\u_cpu.ALU.u_wallace._4657_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5562_  (.A(\u_cpu.ALU.u_wallace._0282_ ),
    .X(\u_cpu.ALU.u_wallace._4658_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5563_  (.A(\u_cpu.ALU.u_wallace._4657_ ),
    .B(\u_cpu.ALU.u_wallace._4658_ ),
    .C(\u_cpu.ALU.u_wallace._4412_ ),
    .D(\u_cpu.ALU.u_wallace._4642_ ),
    .Y(\u_cpu.ALU.u_wallace._4659_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5564_  (.A(\u_cpu.ALU.u_wallace._3645_ ),
    .X(\u_cpu.ALU.u_wallace._4660_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5565_  (.A(\u_cpu.ALU.u_wallace._4660_ ),
    .X(\u_cpu.ALU.u_wallace._4661_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5566_  (.A(\u_cpu.ALU.u_wallace._0457_ ),
    .X(\u_cpu.ALU.u_wallace._4662_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5567_  (.A(\u_cpu.ALU.u_wallace._4662_ ),
    .X(\u_cpu.ALU.u_wallace._4663_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._5568_  (.A_N(\u_cpu.ALU.u_wallace._4656_ ),
    .B(\u_cpu.ALU.u_wallace._4659_ ),
    .C(\u_cpu.ALU.u_wallace._4661_ ),
    .D(\u_cpu.ALU.u_wallace._4663_ ),
    .Y(\u_cpu.ALU.u_wallace._4664_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5569_  (.A(\u_cpu.ALU.u_wallace._0206_ ),
    .B(\u_cpu.ALU.u_wallace._0490_ ),
    .C(\u_cpu.ALU.u_wallace._4444_ ),
    .D(\u_cpu.ALU.u_wallace._4557_ ),
    .X(\u_cpu.ALU.u_wallace._4665_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5570_  (.A(\u_cpu.ALU.u_wallace._4449_ ),
    .B(\u_cpu.ALU.u_wallace._0753_ ),
    .Y(\u_cpu.ALU.u_wallace._4666_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5571_  (.A1(\u_cpu.ALU.u_wallace._4656_ ),
    .A2(\u_cpu.ALU.u_wallace._4665_ ),
    .B1(\u_cpu.ALU.u_wallace._4666_ ),
    .Y(\u_cpu.ALU.u_wallace._4667_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5572_  (.A1(\u_cpu.ALU.u_wallace._4652_ ),
    .A2(\u_cpu.ALU.u_wallace._4655_ ),
    .B1(\u_cpu.ALU.u_wallace._4664_ ),
    .B2(\u_cpu.ALU.u_wallace._4667_ ),
    .Y(\u_cpu.ALU.u_wallace._4668_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5573_  (.A(\u_cpu.ALU.u_wallace._4561_ ),
    .X(\u_cpu.ALU.u_wallace._4669_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5574_  (.A(\u_cpu.ALU.u_wallace._4659_ ),
    .B(\u_cpu.ALU.u_wallace._0468_ ),
    .C(\u_cpu.ALU.u_wallace._4669_ ),
    .Y(\u_cpu.ALU.u_wallace._4670_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._5575_  (.A1(\u_cpu.ALU.u_wallace._4670_ ),
    .A2(\u_cpu.ALU.u_wallace._4656_ ),
    .B1(\u_cpu.ALU.u_wallace._4655_ ),
    .C1(\u_cpu.ALU.u_wallace._4652_ ),
    .D1(\u_cpu.ALU.u_wallace._4667_ ),
    .X(\u_cpu.ALU.u_wallace._4671_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._5576_  (.A1(\u_cpu.ALU.u_wallace._4552_ ),
    .A2(\u_cpu.ALU.u_wallace._4555_ ),
    .B1(\u_cpu.ALU.u_wallace._4668_ ),
    .B2(\u_cpu.ALU.u_wallace._4671_ ),
    .C1(\u_cpu.ALU.u_wallace._4581_ ),
    .X(\u_cpu.ALU.u_wallace._4672_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5577_  (.A(\u_cpu.ALU.u_wallace._4445_ ),
    .B(\u_cpu.ALU.u_wallace._4571_ ),
    .C(\u_cpu.ALU.u_wallace._4572_ ),
    .X(\u_cpu.ALU.u_wallace._4673_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._5578_  (.A1(\u_cpu.ALU.u_wallace._4565_ ),
    .A2(\u_cpu.ALU.u_wallace._4569_ ),
    .A3(\u_cpu.ALU.u_wallace._4559_ ),
    .B1(\u_cpu.ALU.u_wallace._4673_ ),
    .Y(\u_cpu.ALU.u_wallace._4674_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5579_  (.A(\u_cpu.ALU.u_wallace._4656_ ),
    .B(\u_cpu.ALU.u_wallace._4670_ ),
    .Y(\u_cpu.ALU.u_wallace._4675_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._5580_  (.A(\u_cpu.ALU.SrcA[8] ),
    .Y(\u_cpu.ALU.u_wallace._4676_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5581_  (.A(\u_cpu.ALU.u_wallace._4676_ ),
    .X(\u_cpu.ALU.u_wallace._4677_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5582_  (.A(\u_cpu.ALU.u_wallace._1224_ ),
    .X(\u_cpu.ALU.u_wallace._4678_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._5583_  (.A1(\u_cpu.ALU.u_wallace._4677_ ),
    .A2(\u_cpu.ALU.u_wallace._4678_ ),
    .B1(\u_cpu.ALU.u_wallace._4656_ ),
    .B2(\u_cpu.ALU.u_wallace._4665_ ),
    .X(\u_cpu.ALU.u_wallace._4679_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5584_  (.A1_N(\u_cpu.ALU.u_wallace._4652_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4655_ ),
    .B1(\u_cpu.ALU.u_wallace._4675_ ),
    .B2(\u_cpu.ALU.u_wallace._4679_ ),
    .Y(\u_cpu.ALU.u_wallace._4680_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._5585_  (.A1(\u_cpu.ALU.u_wallace._4670_ ),
    .A2(\u_cpu.ALU.u_wallace._4656_ ),
    .B1(\u_cpu.ALU.u_wallace._4655_ ),
    .C1(\u_cpu.ALU.u_wallace._4652_ ),
    .D1(\u_cpu.ALU.u_wallace._4667_ ),
    .Y(\u_cpu.ALU.u_wallace._4681_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5586_  (.A(\u_cpu.ALU.u_wallace._4680_ ),
    .B(\u_cpu.ALU.u_wallace._4681_ ),
    .Y(\u_cpu.ALU.u_wallace._4682_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5587_  (.A(\u_cpu.ALU.u_wallace._4528_ ),
    .B(\u_cpu.ALU.u_wallace._4542_ ),
    .C(\u_cpu.ALU.u_wallace._4541_ ),
    .X(\u_cpu.ALU.u_wallace._4683_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5588_  (.A1(\u_cpu.ALU.u_wallace._4450_ ),
    .A2(\u_cpu.ALU.u_wallace._4467_ ),
    .B1(\u_cpu.ALU.u_wallace._2078_ ),
    .B2(\u_cpu.ALU.u_wallace._1793_ ),
    .X(\u_cpu.ALU.u_wallace._4684_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5589_  (.A(\u_cpu.ALU.u_wallace._2725_ ),
    .B(\u_cpu.ALU.u_wallace._3777_ ),
    .C(\u_cpu.ALU.u_wallace._2571_ ),
    .D(\u_cpu.ALU.u_wallace._2582_ ),
    .Y(\u_cpu.ALU.u_wallace._4685_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._5590_  (.A(\u_cpu.ALU.u_wallace._1267_ ),
    .B(\u_cpu.ALU.SrcB[7] ),
    .X(\u_cpu.ALU.u_wallace._4686_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5591_  (.A(\u_cpu.ALU.u_wallace._4684_ ),
    .B(\u_cpu.ALU.u_wallace._4685_ ),
    .C(\u_cpu.ALU.u_wallace._4686_ ),
    .X(\u_cpu.ALU.u_wallace._4687_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5592_  (.A(\u_cpu.ALU.u_wallace._4564_ ),
    .B(\u_cpu.ALU.u_wallace._4560_ ),
    .Y(\u_cpu.ALU.u_wallace._4688_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5593_  (.A1(\u_cpu.ALU.u_wallace._3821_ ),
    .A2(\u_cpu.ALU.u_wallace._2155_ ),
    .B1(\u_cpu.ALU.u_wallace._2187_ ),
    .B2(\u_cpu.ALU.u_wallace._1848_ ),
    .Y(\u_cpu.ALU.u_wallace._4689_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5594_  (.A(\u_cpu.ALU.u_wallace._4450_ ),
    .B(\u_cpu.ALU.u_wallace._1793_ ),
    .C(\u_cpu.ALU.u_wallace._2571_ ),
    .D(\u_cpu.ALU.u_wallace._2078_ ),
    .X(\u_cpu.ALU.u_wallace._4690_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5595_  (.A1(\u_cpu.ALU.u_wallace._0939_ ),
    .A2(\u_cpu.ALU.u_wallace._4471_ ),
    .B1(\u_cpu.ALU.u_wallace._4689_ ),
    .B2(\u_cpu.ALU.u_wallace._4690_ ),
    .Y(\u_cpu.ALU.u_wallace._4691_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5596_  (.A1(\u_cpu.ALU.u_wallace._4563_ ),
    .A2(\u_cpu.ALU.u_wallace._4688_ ),
    .B1(\u_cpu.ALU.u_wallace._4691_ ),
    .Y(\u_cpu.ALU.u_wallace._4692_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5597_  (.A1(\u_cpu.ALU.u_wallace._4684_ ),
    .A2(\u_cpu.ALU.u_wallace._4685_ ),
    .B1(\u_cpu.ALU.u_wallace._4686_ ),
    .Y(\u_cpu.ALU.u_wallace._4693_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._5598_  (.A1(\u_cpu.ALU.u_wallace._4560_ ),
    .A2(\u_cpu.ALU.u_wallace._4564_ ),
    .B1(\u_cpu.ALU.u_wallace._4693_ ),
    .B2(\u_cpu.ALU.u_wallace._4687_ ),
    .C1(\u_cpu.ALU.u_wallace._4568_ ),
    .Y(\u_cpu.ALU.u_wallace._4694_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._5599_  (.A1(\u_cpu.ALU.u_wallace._4534_ ),
    .A2(\u_cpu.ALU.u_wallace._4683_ ),
    .B1(\u_cpu.ALU.u_wallace._4687_ ),
    .B2(\u_cpu.ALU.u_wallace._4692_ ),
    .C1(\u_cpu.ALU.u_wallace._4694_ ),
    .Y(\u_cpu.ALU.u_wallace._4695_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5600_  (.A(\u_cpu.ALU.u_wallace._4684_ ),
    .B(\u_cpu.ALU.u_wallace._4685_ ),
    .C(\u_cpu.ALU.u_wallace._0917_ ),
    .D(\u_cpu.ALU.u_wallace._3481_ ),
    .Y(\u_cpu.ALU.u_wallace._4696_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5601_  (.A1(\u_cpu.ALU.u_wallace._4563_ ),
    .A2(\u_cpu.ALU.u_wallace._4688_ ),
    .B1(\u_cpu.ALU.u_wallace._4696_ ),
    .C1(\u_cpu.ALU.u_wallace._4691_ ),
    .X(\u_cpu.ALU.u_wallace._4697_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5602_  (.A(\u_cpu.ALU.u_wallace._2725_ ),
    .X(\u_cpu.ALU.u_wallace._4698_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._5603_  (.A1(\u_cpu.ALU.u_wallace._4566_ ),
    .A2(\u_cpu.ALU.u_wallace._0983_ ),
    .A3(\u_cpu.ALU.u_wallace._4698_ ),
    .B1(\u_cpu.ALU.u_wallace._4563_ ),
    .X(\u_cpu.ALU.u_wallace._4699_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5604_  (.A1(\u_cpu.ALU.u_wallace._4696_ ),
    .A2(\u_cpu.ALU.u_wallace._4691_ ),
    .B1(\u_cpu.ALU.u_wallace._4699_ ),
    .Y(\u_cpu.ALU.u_wallace._4700_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._5605_  (.A1(\u_cpu.ALU.u_wallace._0621_ ),
    .A2(\u_cpu.ALU.u_wallace._4539_ ),
    .A3(\u_cpu.ALU.u_wallace._4532_ ),
    .B1(\u_cpu.ALU.u_wallace._4530_ ),
    .X(\u_cpu.ALU.u_wallace._4701_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5606_  (.A1(\u_cpu.ALU.u_wallace._4697_ ),
    .A2(\u_cpu.ALU.u_wallace._4700_ ),
    .B1(\u_cpu.ALU.u_wallace._4701_ ),
    .Y(\u_cpu.ALU.u_wallace._4702_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5607_  (.A1(\u_cpu.ALU.u_wallace._4674_ ),
    .A2(\u_cpu.ALU.u_wallace._4682_ ),
    .B1(\u_cpu.ALU.u_wallace._4695_ ),
    .C1(\u_cpu.ALU.u_wallace._4702_ ),
    .Y(\u_cpu.ALU.u_wallace._4703_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5608_  (.A(\u_cpu.ALU.u_wallace._4581_ ),
    .B(\u_cpu.ALU.u_wallace._4582_ ),
    .C(\u_cpu.ALU.u_wallace._4579_ ),
    .X(\u_cpu.ALU.u_wallace._4704_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5609_  (.A1(\u_cpu.ALU.u_wallace._4587_ ),
    .A2(\u_cpu.ALU.u_wallace._4586_ ),
    .B1(\u_cpu.ALU.u_wallace._4547_ ),
    .C1(\u_cpu.ALU.u_wallace._4580_ ),
    .X(\u_cpu.ALU.u_wallace._4705_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._5610_  (.A1(\u_cpu.ALU.u_wallace._4565_ ),
    .A2(\u_cpu.ALU.u_wallace._4569_ ),
    .A3(\u_cpu.ALU.u_wallace._4559_ ),
    .B1(\u_cpu.ALU.u_wallace._4673_ ),
    .X(\u_cpu.ALU.u_wallace._4706_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5611_  (.A(\u_cpu.ALU.u_wallace._4706_ ),
    .B(\u_cpu.ALU.u_wallace._4680_ ),
    .C(\u_cpu.ALU.u_wallace._4681_ ),
    .Y(\u_cpu.ALU.u_wallace._4707_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5612_  (.A1(\u_cpu.ALU.u_wallace._4668_ ),
    .A2(\u_cpu.ALU.u_wallace._4671_ ),
    .B1(\u_cpu.ALU.u_wallace._4674_ ),
    .Y(\u_cpu.ALU.u_wallace._4708_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._5613_  (.A1(\u_cpu.ALU.u_wallace._4534_ ),
    .A2(\u_cpu.ALU.u_wallace._4683_ ),
    .B1(\u_cpu.ALU.u_wallace._4687_ ),
    .B2(\u_cpu.ALU.u_wallace._4692_ ),
    .C1(\u_cpu.ALU.u_wallace._4694_ ),
    .X(\u_cpu.ALU.u_wallace._4709_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._5614_  (.A1(\u_cpu.ALU.u_wallace._4697_ ),
    .A2(\u_cpu.ALU.u_wallace._4700_ ),
    .B1(\u_cpu.ALU.u_wallace._4701_ ),
    .X(\u_cpu.ALU.u_wallace._4710_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5615_  (.A1_N(\u_cpu.ALU.u_wallace._4707_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4708_ ),
    .B1(\u_cpu.ALU.u_wallace._4709_ ),
    .B2(\u_cpu.ALU.u_wallace._4710_ ),
    .Y(\u_cpu.ALU.u_wallace._4711_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._5616_  (.A1(\u_cpu.ALU.u_wallace._4672_ ),
    .A2(\u_cpu.ALU.u_wallace._4703_ ),
    .B1(\u_cpu.ALU.u_wallace._4704_ ),
    .B2(\u_cpu.ALU.u_wallace._4705_ ),
    .C1(\u_cpu.ALU.u_wallace._4711_ ),
    .Y(\u_cpu.ALU.u_wallace._4712_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5617_  (.A1(\u_cpu.ALU.u_wallace._4672_ ),
    .A2(\u_cpu.ALU.u_wallace._4703_ ),
    .B1(\u_cpu.ALU.u_wallace._4711_ ),
    .Y(\u_cpu.ALU.u_wallace._4713_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._5618_  (.A1(\u_cpu.ALU.u_wallace._4547_ ),
    .A2(\u_cpu.ALU.u_wallace._4549_ ),
    .A3(\u_cpu.ALU.u_wallace._4580_ ),
    .B1(\u_cpu.ALU.u_wallace._4704_ ),
    .Y(\u_cpu.ALU.u_wallace._4714_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5619_  (.A(\u_cpu.ALU.u_wallace._4713_ ),
    .B(\u_cpu.ALU.u_wallace._4714_ ),
    .Y(\u_cpu.ALU.u_wallace._4715_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5620_  (.A(\u_cpu.ALU.SrcB[8] ),
    .X(\u_cpu.ALU.u_wallace._4716_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5621_  (.A(\u_cpu.ALU.u_wallace._4716_ ),
    .X(\u_cpu.ALU.u_wallace._4717_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5622_  (.A(\u_cpu.ALU.u_wallace._0731_ ),
    .B(\u_cpu.ALU.u_wallace._4609_ ),
    .Y(\u_cpu.ALU.u_wallace._4718_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._5623_  (.A1(\u_cpu.ALU.u_wallace._4545_ ),
    .A2(\u_cpu.ALU.u_wallace._4527_ ),
    .A3(\u_cpu.ALU.u_wallace._4717_ ),
    .A4(\u_cpu.ALU.u_wallace._4313_ ),
    .B1(\u_cpu.ALU.u_wallace._4718_ ),
    .X(\u_cpu.ALU.u_wallace._4719_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5624_  (.A(\u_cpu.ALU.SrcB[8] ),
    .X(\u_cpu.ALU.u_wallace._4720_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5625_  (.A1(\u_cpu.ALU.u_wallace._1278_ ),
    .A2(\u_cpu.ALU.u_wallace._4720_ ),
    .B1(\u_cpu.ALU.u_wallace._4595_ ),
    .B2(\u_cpu.ALU.u_wallace._0348_ ),
    .Y(\u_cpu.ALU.u_wallace._4721_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5626_  (.A(\u_cpu.ALU.u_wallace._0446_ ),
    .B(\u_cpu.ALU.u_wallace._4604_ ),
    .Y(\u_cpu.ALU.u_wallace._4722_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5627_  (.A1(\u_cpu.ALU.u_wallace._4597_ ),
    .A2(\u_cpu.ALU.u_wallace._4717_ ),
    .B1(\u_cpu.ALU.u_wallace._4599_ ),
    .B2(\u_cpu.ALU.u_wallace._1454_ ),
    .Y(\u_cpu.ALU.u_wallace._4723_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5628_  (.A1(\u_cpu.ALU.u_wallace._4722_ ),
    .A2(\u_cpu.ALU.u_wallace._4723_ ),
    .B1(\u_cpu.ALU.u_wallace._4600_ ),
    .Y(\u_cpu.ALU.u_wallace._4724_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5629_  (.A(\u_cpu.ALU.u_wallace._0512_ ),
    .B(\u_cpu.ALU.u_wallace._1191_ ),
    .C(\u_cpu.ALU.u_wallace._4594_ ),
    .D(\u_cpu.ALU.u_wallace._4595_ ),
    .X(\u_cpu.ALU.u_wallace._4725_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5630_  (.A1(\u_cpu.ALU.u_wallace._4721_ ),
    .A2(\u_cpu.ALU.u_wallace._4725_ ),
    .B1(\u_cpu.ALU.u_wallace._4718_ ),
    .Y(\u_cpu.ALU.u_wallace._4726_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5631_  (.A1(\u_cpu.ALU.u_wallace._4719_ ),
    .A2(\u_cpu.ALU.u_wallace._4721_ ),
    .B1(\u_cpu.ALU.u_wallace._4724_ ),
    .C1(\u_cpu.ALU.u_wallace._4726_ ),
    .X(\u_cpu.ALU.u_wallace._4727_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5632_  (.A(\u_cpu.ALU.u_wallace._1410_ ),
    .B(\u_cpu.ALU.u_wallace._1421_ ),
    .C(\u_cpu.ALU.u_wallace._4018_ ),
    .D(\u_cpu.ALU.u_wallace._4302_ ),
    .Y(\u_cpu.ALU.u_wallace._4728_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._5633_  (.A_N(\u_cpu.ALU.u_wallace._4721_ ),
    .B(\u_cpu.ALU.u_wallace._4728_ ),
    .C(\u_cpu.ALU.u_wallace._0162_ ),
    .D(\u_cpu.ALU.u_wallace._4610_ ),
    .Y(\u_cpu.ALU.u_wallace._4729_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5634_  (.A1(\u_cpu.ALU.u_wallace._4726_ ),
    .A2(\u_cpu.ALU.u_wallace._4729_ ),
    .B1(\u_cpu.ALU.u_wallace._4724_ ),
    .X(\u_cpu.ALU.u_wallace._4730_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5635_  (.A(\u_cpu.ALU.SrcB[11] ),
    .X(\u_cpu.ALU.u_wallace._4731_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5636_  (.A(\u_cpu.ALU.u_wallace._4731_ ),
    .X(\u_cpu.ALU.u_wallace._4732_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5637_  (.A(\u_cpu.ALU.u_wallace._4732_ ),
    .X(\u_cpu.ALU.u_wallace._4733_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5638_  (.A(\u_cpu.ALU.u_wallace._4730_ ),
    .B(\u_cpu.ALU.u_wallace._4733_ ),
    .C(\u_cpu.ALU.u_wallace._3996_ ),
    .Y(\u_cpu.ALU.u_wallace._4734_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5639_  (.A1(\u_cpu.ALU.u_wallace._4535_ ),
    .A2(\u_cpu.ALU.u_wallace._4548_ ),
    .B1(\u_cpu.ALU.u_wallace._4538_ ),
    .C1(\u_cpu.ALU.u_wallace._4546_ ),
    .X(\u_cpu.ALU.u_wallace._4735_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5640_  (.A1(\u_cpu.ALU.u_wallace._4719_ ),
    .A2(\u_cpu.ALU.u_wallace._4721_ ),
    .B1(\u_cpu.ALU.u_wallace._4724_ ),
    .C1(\u_cpu.ALU.u_wallace._4726_ ),
    .Y(\u_cpu.ALU.u_wallace._4736_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5641_  (.A1(\u_cpu.ALU.u_wallace._3996_ ),
    .A2(\u_cpu.ALU.u_wallace._4733_ ),
    .B1(\u_cpu.ALU.u_wallace._4736_ ),
    .B2(\u_cpu.ALU.u_wallace._4730_ ),
    .X(\u_cpu.ALU.u_wallace._4737_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._5642_  (.A1(\u_cpu.ALU.u_wallace._4727_ ),
    .A2(\u_cpu.ALU.u_wallace._4734_ ),
    .B1(\u_cpu.ALU.u_wallace._4586_ ),
    .B2(\u_cpu.ALU.u_wallace._4735_ ),
    .C1(\u_cpu.ALU.u_wallace._4737_ ),
    .Y(\u_cpu.ALU.u_wallace._4738_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5643_  (.A1(\u_cpu.ALU.u_wallace._4546_ ),
    .A2(\u_cpu.ALU.u_wallace._4538_ ),
    .B1(\u_cpu.ALU.u_wallace._4586_ ),
    .Y(\u_cpu.ALU.u_wallace._4739_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5644_  (.A1(\u_cpu.ALU.u_wallace._4726_ ),
    .A2(\u_cpu.ALU.u_wallace._4729_ ),
    .B1(\u_cpu.ALU.u_wallace._4724_ ),
    .Y(\u_cpu.ALU.u_wallace._4740_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5645_  (.A1(\u_cpu.ALU.u_wallace._4727_ ),
    .A2(\u_cpu.ALU.u_wallace._4740_ ),
    .B1(\u_cpu.ALU.u_wallace._0129_ ),
    .C1(\u_cpu.ALU.u_wallace._4733_ ),
    .Y(\u_cpu.ALU.u_wallace._4741_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5646_  (.A(\u_cpu.ALU.u_wallace._3996_ ),
    .B(\u_cpu.ALU.u_wallace._4733_ ),
    .Y(\u_cpu.ALU.u_wallace._4742_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5647_  (.A(\u_cpu.ALU.u_wallace._4742_ ),
    .B(\u_cpu.ALU.u_wallace._4736_ ),
    .C(\u_cpu.ALU.u_wallace._4730_ ),
    .Y(\u_cpu.ALU.u_wallace._4743_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5648_  (.A(\u_cpu.ALU.u_wallace._4739_ ),
    .B(\u_cpu.ALU.u_wallace._4741_ ),
    .C(\u_cpu.ALU.u_wallace._4743_ ),
    .Y(\u_cpu.ALU.u_wallace._4744_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU.u_wallace._5649_  (.A1(\u_cpu.ALU.u_wallace._4611_ ),
    .A2(\u_cpu.ALU.u_wallace._4596_ ),
    .B1(\u_cpu.ALU.u_wallace._4607_ ),
    .C1(\u_cpu.ALU.u_wallace._4603_ ),
    .Y(\u_cpu.ALU.u_wallace._4745_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5650_  (.A(\u_cpu.ALU.u_wallace._4738_ ),
    .B(\u_cpu.ALU.u_wallace._4744_ ),
    .C(\u_cpu.ALU.u_wallace._4745_ ),
    .X(\u_cpu.ALU.u_wallace._4746_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5651_  (.A1(\u_cpu.ALU.u_wallace._4738_ ),
    .A2(\u_cpu.ALU.u_wallace._4744_ ),
    .B1(\u_cpu.ALU.u_wallace._4745_ ),
    .Y(\u_cpu.ALU.u_wallace._4747_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5652_  (.A1_N(\u_cpu.ALU.u_wallace._4712_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4715_ ),
    .B1(\u_cpu.ALU.u_wallace._4746_ ),
    .B2(\u_cpu.ALU.u_wallace._4747_ ),
    .Y(\u_cpu.ALU.u_wallace._4748_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._5653_  (.A1(\u_cpu.ALU.u_wallace._4739_ ),
    .A2(\u_cpu.ALU.u_wallace._4741_ ),
    .A3(\u_cpu.ALU.u_wallace._4743_ ),
    .B1(\u_cpu.ALU.u_wallace._4612_ ),
    .Y(\u_cpu.ALU.u_wallace._4749_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5654_  (.A(\u_cpu.ALU.u_wallace._4749_ ),
    .B(\u_cpu.ALU.u_wallace._4738_ ),
    .Y(\u_cpu.ALU.u_wallace._4750_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5655_  (.A1(\u_cpu.ALU.u_wallace._4738_ ),
    .A2(\u_cpu.ALU.u_wallace._4744_ ),
    .B1(\u_cpu.ALU.u_wallace._4745_ ),
    .X(\u_cpu.ALU.u_wallace._4751_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5656_  (.A(\u_cpu.ALU.u_wallace._4712_ ),
    .B(\u_cpu.ALU.u_wallace._4715_ ),
    .C(\u_cpu.ALU.u_wallace._4750_ ),
    .D(\u_cpu.ALU.u_wallace._4751_ ),
    .Y(\u_cpu.ALU.u_wallace._4752_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5657_  (.A(\u_cpu.ALU.u_wallace._4641_ ),
    .B(\u_cpu.ALU.u_wallace._4748_ ),
    .C(\u_cpu.ALU.u_wallace._4752_ ),
    .Y(\u_cpu.ALU.u_wallace._4753_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5658_  (.A1(\u_cpu.ALU.u_wallace._4748_ ),
    .A2(\u_cpu.ALU.u_wallace._4752_ ),
    .B1(\u_cpu.ALU.u_wallace._4641_ ),
    .X(\u_cpu.ALU.u_wallace._4754_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._5659_  (.A1(\u_cpu.ALU.u_wallace._4481_ ),
    .A2(\u_cpu.ALU.u_wallace._4480_ ),
    .B1(\u_cpu.ALU.u_wallace._4474_ ),
    .X(\u_cpu.ALU.u_wallace._4755_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5660_  (.A1_N(\u_cpu.ALU.u_wallace._4753_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4754_ ),
    .B1(\u_cpu.ALU.u_wallace._4755_ ),
    .B2(\u_cpu.ALU.u_wallace._4615_ ),
    .Y(\u_cpu.ALU.u_wallace._4756_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5661_  (.A(\u_cpu.ALU.u_wallace._4754_ ),
    .B(\u_cpu.ALU.u_wallace._4613_ ),
    .C(\u_cpu.ALU.u_wallace._4753_ ),
    .Y(\u_cpu.ALU.u_wallace._4757_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5662_  (.A(\u_cpu.ALU.u_wallace._4640_ ),
    .B(\u_cpu.ALU.u_wallace._4756_ ),
    .C(\u_cpu.ALU.u_wallace._4757_ ),
    .Y(\u_cpu.ALU.u_wallace._4758_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5663_  (.A1(\u_cpu.ALU.u_wallace._4756_ ),
    .A2(\u_cpu.ALU.u_wallace._4757_ ),
    .B1(\u_cpu.ALU.u_wallace._4640_ ),
    .X(\u_cpu.ALU.u_wallace._4759_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._5664_  (.A1(\u_cpu.ALU.u_wallace._4638_ ),
    .A2(\u_cpu.ALU.u_wallace._4639_ ),
    .B1(\u_cpu.ALU.u_wallace._4758_ ),
    .C1(\u_cpu.ALU.u_wallace._4759_ ),
    .D1(\u_cpu.ALU.u_wallace._4633_ ),
    .Y(\u_cpu.ALU.u_wallace._4760_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._5665_  (.A1(\u_cpu.ALU.u_wallace._4525_ ),
    .A2(\u_cpu.ALU.u_wallace._4625_ ),
    .A3(\u_cpu.ALU.u_wallace._4629_ ),
    .B1(\u_cpu.ALU.u_wallace._4639_ ),
    .X(\u_cpu.ALU.u_wallace._4761_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5666_  (.A1(\u_cpu.ALU.u_wallace._4633_ ),
    .A2(\u_cpu.ALU.u_wallace._4761_ ),
    .B1(\u_cpu.ALU.u_wallace._4758_ ),
    .B2(\u_cpu.ALU.u_wallace._4759_ ),
    .X(\u_cpu.ALU.u_wallace._4762_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5667_  (.A(\u_cpu.ALU.u_wallace._4139_ ),
    .B(\u_cpu.ALU.u_wallace._4499_ ),
    .C(\u_cpu.ALU.u_wallace._4508_ ),
    .D(\u_cpu.ALU.u_wallace._3251_ ),
    .X(\u_cpu.ALU.u_wallace._4763_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5668_  (.A1(\u_cpu.ALU.u_wallace._4513_ ),
    .A2(\u_cpu.ALU.u_wallace._4516_ ),
    .B1(\u_cpu.ALU.u_wallace._4763_ ),
    .B2(\u_cpu.ALU.u_wallace._4636_ ),
    .Y(\u_cpu.ALU.u_wallace._4764_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5669_  (.A1(\u_cpu.ALU.u_wallace._4638_ ),
    .A2(\u_cpu.ALU.u_wallace._4639_ ),
    .B1(\u_cpu.ALU.u_wallace._4519_ ),
    .X(\u_cpu.ALU.u_wallace._4765_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5670_  (.A1(\u_cpu.ALU.u_wallace._4760_ ),
    .A2(\u_cpu.ALU.u_wallace._4762_ ),
    .B1(\u_cpu.ALU.u_wallace._4764_ ),
    .B2(\u_cpu.ALU.u_wallace._4765_ ),
    .Y(\u_cpu.ALU.u_wallace._4766_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5671_  (.A(\u_cpu.ALU.u_wallace._4765_ ),
    .B(\u_cpu.ALU.u_wallace._4760_ ),
    .C(\u_cpu.ALU.u_wallace._4762_ ),
    .D(\u_cpu.ALU.u_wallace._4764_ ),
    .X(\u_cpu.ALU.u_wallace._4767_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5672_  (.A(\u_cpu.ALU.u_wallace._4766_ ),
    .B(\u_cpu.ALU.u_wallace._4767_ ),
    .Y(\u_cpu.ALU.Product_Wallace[11] ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5673_  (.A1(\u_cpu.ALU.u_wallace._4756_ ),
    .A2(\u_cpu.ALU.u_wallace._4757_ ),
    .B1(\u_cpu.ALU.u_wallace._4640_ ),
    .Y(\u_cpu.ALU.u_wallace._4768_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._5674_  (.A1(\u_cpu.ALU.u_wallace._4641_ ),
    .A2(\u_cpu.ALU.u_wallace._4748_ ),
    .A3(\u_cpu.ALU.u_wallace._4752_ ),
    .B1(\u_cpu.ALU.u_wallace._4754_ ),
    .B2(\u_cpu.ALU.u_wallace._4613_ ),
    .X(\u_cpu.ALU.u_wallace._4769_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._5675_  (.A(\u_cpu.ALU.u_wallace._4738_ ),
    .B(\u_cpu.ALU.u_wallace._4750_ ),
    .X(\u_cpu.ALU.u_wallace._4770_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._5676_  (.A1(\u_cpu.ALU.u_wallace._4672_ ),
    .A2(\u_cpu.ALU.u_wallace._4703_ ),
    .B1(\u_cpu.ALU.u_wallace._4704_ ),
    .B2(\u_cpu.ALU.u_wallace._4705_ ),
    .C1(\u_cpu.ALU.u_wallace._4711_ ),
    .X(\u_cpu.ALU.u_wallace._4771_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.ALU.u_wallace._5677_  (.A1(\u_cpu.ALU.u_wallace._4738_ ),
    .A2(\u_cpu.ALU.u_wallace._4749_ ),
    .B1(\u_cpu.ALU.u_wallace._4713_ ),
    .B2(\u_cpu.ALU.u_wallace._4714_ ),
    .C1(\u_cpu.ALU.u_wallace._4747_ ),
    .Y(\u_cpu.ALU.u_wallace._4772_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5678_  (.A1(\u_cpu.ALU.u_wallace._4576_ ),
    .A2(\u_cpu.ALU.u_wallace._4581_ ),
    .B1(\u_cpu.ALU.u_wallace._4682_ ),
    .Y(\u_cpu.ALU.u_wallace._4773_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5679_  (.A1(\u_cpu.ALU.u_wallace._4534_ ),
    .A2(\u_cpu.ALU.u_wallace._4683_ ),
    .B1(\u_cpu.ALU.u_wallace._4697_ ),
    .B2(\u_cpu.ALU.u_wallace._4700_ ),
    .Y(\u_cpu.ALU.u_wallace._4774_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5680_  (.A1(\u_cpu.ALU.u_wallace._4563_ ),
    .A2(\u_cpu.ALU.u_wallace._4688_ ),
    .B1(\u_cpu.ALU.u_wallace._4696_ ),
    .C1(\u_cpu.ALU.u_wallace._4691_ ),
    .Y(\u_cpu.ALU.u_wallace._4775_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._5681_  (.A1(\u_cpu.ALU.u_wallace._4533_ ),
    .A2(\u_cpu.ALU.u_wallace._4532_ ),
    .B1(\u_cpu.ALU.u_wallace._4530_ ),
    .C1(\u_cpu.ALU.u_wallace._4775_ ),
    .D1(\u_cpu.ALU.u_wallace._4694_ ),
    .Y(\u_cpu.ALU.u_wallace._4776_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5682_  (.A1(\u_cpu.ALU.u_wallace._4674_ ),
    .A2(\u_cpu.ALU.u_wallace._4682_ ),
    .B1(\u_cpu.ALU.u_wallace._4774_ ),
    .B2(\u_cpu.ALU.u_wallace._4776_ ),
    .Y(\u_cpu.ALU.u_wallace._4777_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5683_  (.A1(\u_cpu.ALU.u_wallace._4670_ ),
    .A2(\u_cpu.ALU.u_wallace._4656_ ),
    .B1(\u_cpu.ALU.u_wallace._4652_ ),
    .C1(\u_cpu.ALU.u_wallace._4667_ ),
    .Y(\u_cpu.ALU.u_wallace._4778_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5684_  (.A(\u_cpu.ALU.u_wallace._4655_ ),
    .B(\u_cpu.ALU.u_wallace._4778_ ),
    .Y(\u_cpu.ALU.u_wallace._4779_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5685_  (.A(\u_cpu.ALU.u_wallace._1957_ ),
    .B(\u_cpu.ALU.u_wallace._4658_ ),
    .C(\u_cpu.ALU.u_wallace._4642_ ),
    .D(\u_cpu.ALU.u_wallace._4647_ ),
    .Y(\u_cpu.ALU.u_wallace._4780_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5686_  (.A1(\u_cpu.ALU.u_wallace._0490_ ),
    .A2(\u_cpu.ALU.u_wallace._4557_ ),
    .B1(\u_cpu.ALU.u_wallace._4647_ ),
    .B2(\u_cpu.ALU.u_wallace._0206_ ),
    .X(\u_cpu.ALU.u_wallace._4781_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5687_  (.A1_N(\u_cpu.ALU.u_wallace._4780_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4781_ ),
    .B1(\u_cpu.ALU.u_wallace._1892_ ),
    .B2(\u_cpu.ALU.u_wallace._4573_ ),
    .Y(\u_cpu.ALU.u_wallace._4782_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5688_  (.A(\u_cpu.ALU.u_wallace._4562_ ),
    .X(\u_cpu.ALU.u_wallace._4783_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5689_  (.A(\u_cpu.ALU.u_wallace._4781_ ),
    .B(\u_cpu.ALU.u_wallace._4783_ ),
    .C(\u_cpu.ALU.u_wallace._0468_ ),
    .D(\u_cpu.ALU.u_wallace._4780_ ),
    .Y(\u_cpu.ALU.u_wallace._4784_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5690_  (.A(\u_cpu.ALU.SrcA[12] ),
    .X(\u_cpu.ALU.u_wallace._4785_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5691_  (.A1(\u_cpu.ALU.u_wallace._4645_ ),
    .A2(\u_cpu.ALU.u_wallace._2834_ ),
    .B1(\u_cpu.ALU.u_wallace._4785_ ),
    .B2(\u_cpu.ALU.u_wallace._2747_ ),
    .Y(\u_cpu.ALU.u_wallace._4786_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5692_  (.A(\u_cpu.ALU.SrcA[12] ),
    .X(\u_cpu.ALU.u_wallace._4787_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5693_  (.A(\u_cpu.ALU.u_wallace._1859_ ),
    .B(\u_cpu.ALU.u_wallace._1826_ ),
    .C(\u_cpu.ALU.u_wallace._3832_ ),
    .D(\u_cpu.ALU.u_wallace._4787_ ),
    .Y(\u_cpu.ALU.u_wallace._4788_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._5694_  (.A_N(\u_cpu.ALU.u_wallace._4786_ ),
    .B(\u_cpu.ALU.u_wallace._4788_ ),
    .C(\u_cpu.ALU.u_wallace._4651_ ),
    .Y(\u_cpu.ALU.u_wallace._4789_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5695_  (.A(\u_cpu.ALU.SrcA[12] ),
    .X(\u_cpu.ALU.u_wallace._4790_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5696_  (.A(\u_cpu.ALU.u_wallace._0064_ ),
    .B(\u_cpu.ALU.u_wallace._4649_ ),
    .C(\u_cpu.ALU.u_wallace._1782_ ),
    .D(\u_cpu.ALU.u_wallace._4790_ ),
    .X(\u_cpu.ALU.u_wallace._4791_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5697_  (.A1(\u_cpu.ALU.u_wallace._4786_ ),
    .A2(\u_cpu.ALU.u_wallace._4791_ ),
    .B1(\u_cpu.ALU.u_wallace._4654_ ),
    .Y(\u_cpu.ALU.u_wallace._4792_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5698_  (.A1(\u_cpu.ALU.u_wallace._4782_ ),
    .A2(\u_cpu.ALU.u_wallace._4784_ ),
    .B1(\u_cpu.ALU.u_wallace._4789_ ),
    .B2(\u_cpu.ALU.u_wallace._4792_ ),
    .X(\u_cpu.ALU.u_wallace._4793_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5699_  (.A(\u_cpu.ALU.u_wallace._4650_ ),
    .X(\u_cpu.ALU.u_wallace._4794_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5700_  (.A1(\u_cpu.ALU.u_wallace._1169_ ),
    .A2(\u_cpu.ALU.u_wallace._4551_ ),
    .B1(\u_cpu.ALU.u_wallace._4794_ ),
    .B2(\u_cpu.ALU.u_wallace._0523_ ),
    .Y(\u_cpu.ALU.u_wallace._4795_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5701_  (.A(\u_cpu.ALU.u_wallace._1914_ ),
    .X(\u_cpu.ALU.u_wallace._4796_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5702_  (.A(\u_cpu.ALU.u_wallace._4646_ ),
    .X(\u_cpu.ALU.u_wallace._4797_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5703_  (.A(\u_cpu.ALU.u_wallace._4797_ ),
    .X(\u_cpu.ALU.u_wallace._4798_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5704_  (.A(\u_cpu.ALU.u_wallace._0753_ ),
    .B(\u_cpu.ALU.u_wallace._4567_ ),
    .Y(\u_cpu.ALU.u_wallace._4799_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._5705_  (.A1(\u_cpu.ALU.u_wallace._0217_ ),
    .A2(\u_cpu.ALU.u_wallace._4796_ ),
    .A3(\u_cpu.ALU.u_wallace._4643_ ),
    .A4(\u_cpu.ALU.u_wallace._4798_ ),
    .B1(\u_cpu.ALU.u_wallace._4799_ ),
    .X(\u_cpu.ALU.u_wallace._4800_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._5706_  (.A1(\u_cpu.ALU.u_wallace._4795_ ),
    .A2(\u_cpu.ALU.u_wallace._4800_ ),
    .B1(\u_cpu.ALU.u_wallace._4789_ ),
    .C1(\u_cpu.ALU.u_wallace._4792_ ),
    .D1(\u_cpu.ALU.u_wallace._4782_ ),
    .Y(\u_cpu.ALU.u_wallace._4801_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5707_  (.A(\u_cpu.ALU.u_wallace._4779_ ),
    .B(\u_cpu.ALU.u_wallace._4793_ ),
    .C(\u_cpu.ALU.u_wallace._4801_ ),
    .Y(\u_cpu.ALU.u_wallace._4802_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5708_  (.A1(\u_cpu.ALU.u_wallace._4782_ ),
    .A2(\u_cpu.ALU.u_wallace._4784_ ),
    .B1(\u_cpu.ALU.u_wallace._4789_ ),
    .B2(\u_cpu.ALU.u_wallace._4792_ ),
    .Y(\u_cpu.ALU.u_wallace._4803_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._5709_  (.A1(\u_cpu.ALU.u_wallace._4795_ ),
    .A2(\u_cpu.ALU.u_wallace._4800_ ),
    .B1(\u_cpu.ALU.u_wallace._4789_ ),
    .C1(\u_cpu.ALU.u_wallace._4792_ ),
    .D1(\u_cpu.ALU.u_wallace._4782_ ),
    .X(\u_cpu.ALU.u_wallace._4804_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._5710_  (.A1(\u_cpu.ALU.u_wallace._4572_ ),
    .A2(\u_cpu.ALU.u_wallace._4648_ ),
    .A3(\u_cpu.ALU.u_wallace._4651_ ),
    .B1(\u_cpu.ALU.u_wallace._4778_ ),
    .X(\u_cpu.ALU.u_wallace._4805_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5711_  (.A1(\u_cpu.ALU.u_wallace._4803_ ),
    .A2(\u_cpu.ALU.u_wallace._4804_ ),
    .B1(\u_cpu.ALU.u_wallace._4805_ ),
    .Y(\u_cpu.ALU.u_wallace._4806_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5712_  (.A(\u_cpu.ALU.u_wallace._4684_ ),
    .B(\u_cpu.ALU.u_wallace._4686_ ),
    .Y(\u_cpu.ALU.u_wallace._4807_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._5713_  (.A1(\u_cpu.ALU.u_wallace._4677_ ),
    .A2(\u_cpu.ALU.u_wallace._1892_ ),
    .A3(\u_cpu.ALU.u_wallace._4656_ ),
    .B1(\u_cpu.ALU.u_wallace._4659_ ),
    .X(\u_cpu.ALU.u_wallace._4808_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5714_  (.A1(\u_cpu.ALU.u_wallace._3689_ ),
    .A2(\u_cpu.ALU.u_wallace._2144_ ),
    .B1(\u_cpu.ALU.u_wallace._1497_ ),
    .B2(\u_cpu.ALU.u_wallace._4447_ ),
    .X(\u_cpu.ALU.u_wallace._4809_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5715_  (.A(\u_cpu.ALU.u_wallace._3623_ ),
    .B(\u_cpu.ALU.u_wallace._4450_ ),
    .C(\u_cpu.ALU.u_wallace._2571_ ),
    .D(\u_cpu.ALU.u_wallace._2078_ ),
    .Y(\u_cpu.ALU.u_wallace._4810_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5716_  (.A(\u_cpu.ALU.u_wallace._4809_ ),
    .B(\u_cpu.ALU.u_wallace._4810_ ),
    .C(\u_cpu.ALU.u_wallace._1322_ ),
    .D(\u_cpu.ALU.u_wallace._2626_ ),
    .Y(\u_cpu.ALU.u_wallace._4811_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._5717_  (.A(\u_cpu.ALU.SrcA[5] ),
    .Y(\u_cpu.ALU.u_wallace._4812_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5718_  (.A(\u_cpu.ALU.u_wallace._4812_ ),
    .X(\u_cpu.ALU.u_wallace._4813_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5719_  (.A1(\u_cpu.ALU.u_wallace._4561_ ),
    .A2(\u_cpu.ALU.u_wallace._1465_ ),
    .B1(\u_cpu.ALU.u_wallace._2582_ ),
    .B2(\u_cpu.ALU.u_wallace._4450_ ),
    .Y(\u_cpu.ALU.u_wallace._4814_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5720_  (.A(\u_cpu.ALU.u_wallace._3645_ ),
    .B(\u_cpu.ALU.u_wallace._2878_ ),
    .C(\u_cpu.ALU.u_wallace._1026_ ),
    .D(\u_cpu.ALU.u_wallace._1541_ ),
    .X(\u_cpu.ALU.u_wallace._4815_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5721_  (.A1(\u_cpu.ALU.u_wallace._4813_ ),
    .A2(\u_cpu.ALU.u_wallace._4471_ ),
    .B1(\u_cpu.ALU.u_wallace._4814_ ),
    .B2(\u_cpu.ALU.u_wallace._4815_ ),
    .Y(\u_cpu.ALU.u_wallace._4816_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5722_  (.A(\u_cpu.ALU.u_wallace._4811_ ),
    .B(\u_cpu.ALU.u_wallace._4816_ ),
    .Y(\u_cpu.ALU.u_wallace._4817_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5723_  (.A(\u_cpu.ALU.u_wallace._4666_ ),
    .B(\u_cpu.ALU.u_wallace._4656_ ),
    .Y(\u_cpu.ALU.u_wallace._4818_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5724_  (.A1(\u_cpu.ALU.u_wallace._4665_ ),
    .A2(\u_cpu.ALU.u_wallace._4818_ ),
    .B1(\u_cpu.ALU.u_wallace._4811_ ),
    .C1(\u_cpu.ALU.u_wallace._4816_ ),
    .X(\u_cpu.ALU.u_wallace._4819_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.ALU.u_wallace._5725_  (.A1(\u_cpu.ALU.u_wallace._4685_ ),
    .A2(\u_cpu.ALU.u_wallace._4807_ ),
    .B1(\u_cpu.ALU.u_wallace._4808_ ),
    .B2(\u_cpu.ALU.u_wallace._4817_ ),
    .C1(\u_cpu.ALU.u_wallace._4819_ ),
    .Y(\u_cpu.ALU.u_wallace._4820_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5726_  (.A1(\u_cpu.ALU.u_wallace._4665_ ),
    .A2(\u_cpu.ALU.u_wallace._4818_ ),
    .B1(\u_cpu.ALU.u_wallace._4811_ ),
    .C1(\u_cpu.ALU.u_wallace._4816_ ),
    .Y(\u_cpu.ALU.u_wallace._4821_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5727_  (.A1(\u_cpu.ALU.u_wallace._4666_ ),
    .A2(\u_cpu.ALU.u_wallace._4656_ ),
    .B1(\u_cpu.ALU.u_wallace._4659_ ),
    .Y(\u_cpu.ALU.u_wallace._4822_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5728_  (.A1(\u_cpu.ALU.u_wallace._4811_ ),
    .A2(\u_cpu.ALU.u_wallace._4816_ ),
    .B1(\u_cpu.ALU.u_wallace._4822_ ),
    .X(\u_cpu.ALU.u_wallace._4823_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._5729_  (.A1(\u_cpu.ALU.u_wallace._4684_ ),
    .A2(\u_cpu.ALU.u_wallace._4542_ ),
    .A3(\u_cpu.ALU.u_wallace._0917_ ),
    .B1(\u_cpu.ALU.u_wallace._4690_ ),
    .X(\u_cpu.ALU.u_wallace._4824_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5730_  (.A1(\u_cpu.ALU.u_wallace._4821_ ),
    .A2(\u_cpu.ALU.u_wallace._4823_ ),
    .B1(\u_cpu.ALU.u_wallace._4824_ ),
    .Y(\u_cpu.ALU.u_wallace._4825_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5731_  (.A1_N(\u_cpu.ALU.u_wallace._4802_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4806_ ),
    .B1(\u_cpu.ALU.u_wallace._4820_ ),
    .B2(\u_cpu.ALU.u_wallace._4825_ ),
    .Y(\u_cpu.ALU.u_wallace._4826_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5732_  (.A1(\u_cpu.ALU.u_wallace._4685_ ),
    .A2(\u_cpu.ALU.u_wallace._4807_ ),
    .B1(\u_cpu.ALU.u_wallace._4817_ ),
    .B2(\u_cpu.ALU.u_wallace._4808_ ),
    .Y(\u_cpu.ALU.u_wallace._4827_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5733_  (.A1(\u_cpu.ALU.u_wallace._4808_ ),
    .A2(\u_cpu.ALU.u_wallace._4817_ ),
    .B1(\u_cpu.ALU.u_wallace._4827_ ),
    .Y(\u_cpu.ALU.u_wallace._4828_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5734_  (.A1(\u_cpu.ALU.u_wallace._4811_ ),
    .A2(\u_cpu.ALU.u_wallace._4816_ ),
    .B1(\u_cpu.ALU.u_wallace._4822_ ),
    .Y(\u_cpu.ALU.u_wallace._4829_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._5735_  (.A1(\u_cpu.ALU.u_wallace._4819_ ),
    .A2(\u_cpu.ALU.u_wallace._4829_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4824_ ),
    .Y(\u_cpu.ALU.u_wallace._4830_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5736_  (.A(\u_cpu.ALU.u_wallace._4802_ ),
    .B(\u_cpu.ALU.u_wallace._4806_ ),
    .C(\u_cpu.ALU.u_wallace._4828_ ),
    .D(\u_cpu.ALU.u_wallace._4830_ ),
    .Y(\u_cpu.ALU.u_wallace._4831_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5737_  (.A1(\u_cpu.ALU.u_wallace._4773_ ),
    .A2(\u_cpu.ALU.u_wallace._4777_ ),
    .B1(\u_cpu.ALU.u_wallace._4826_ ),
    .C1(\u_cpu.ALU.u_wallace._4831_ ),
    .X(\u_cpu.ALU.u_wallace._4832_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._5738_  (.A1(\u_cpu.ALU.u_wallace._4708_ ),
    .A2(\u_cpu.ALU.u_wallace._4695_ ),
    .A3(\u_cpu.ALU.u_wallace._4702_ ),
    .B1(\u_cpu.ALU.u_wallace._4773_ ),
    .X(\u_cpu.ALU.u_wallace._4833_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5739_  (.A1(\u_cpu.ALU.u_wallace._4826_ ),
    .A2(\u_cpu.ALU.u_wallace._4831_ ),
    .B1(\u_cpu.ALU.u_wallace._4833_ ),
    .Y(\u_cpu.ALU.u_wallace._4834_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5740_  (.A1(\u_cpu.ALU.u_wallace._4701_ ),
    .A2(\u_cpu.ALU.u_wallace._4700_ ),
    .B1(\u_cpu.ALU.u_wallace._4775_ ),
    .Y(\u_cpu.ALU.u_wallace._4835_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5741_  (.A(\u_cpu.ALU.SrcB[11] ),
    .X(\u_cpu.ALU.u_wallace._4836_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5742_  (.A(\u_cpu.ALU.u_wallace._4836_ ),
    .X(\u_cpu.ALU.u_wallace._4837_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5743_  (.A(\u_cpu.ALU.SrcB[12] ),
    .X(\u_cpu.ALU.u_wallace._4838_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5744_  (.A(\u_cpu.ALU.u_wallace._0021_ ),
    .B(\u_cpu.ALU.u_wallace._0731_ ),
    .C(\u_cpu.ALU.u_wallace._4837_ ),
    .D(\u_cpu.ALU.u_wallace._4838_ ),
    .X(\u_cpu.ALU.u_wallace._4839_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5745_  (.A(\u_cpu.ALU.u_wallace._4836_ ),
    .X(\u_cpu.ALU.u_wallace._4840_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5746_  (.A(\u_cpu.ALU.SrcB[12] ),
    .X(\u_cpu.ALU.u_wallace._4841_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5747_  (.A(\u_cpu.ALU.u_wallace._4841_ ),
    .X(\u_cpu.ALU.u_wallace._4842_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5748_  (.A1(\u_cpu.ALU.u_wallace._1454_ ),
    .A2(\u_cpu.ALU.u_wallace._4840_ ),
    .B1(\u_cpu.ALU.u_wallace._4842_ ),
    .B2(\u_cpu.ALU.u_wallace._0021_ ),
    .Y(\u_cpu.ALU.u_wallace._4843_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU.u_wallace._5749_  (.A(\u_cpu.ALU.u_wallace._4839_ ),
    .B(\u_cpu.ALU.u_wallace._4843_ ),
    .X(\u_cpu.ALU.u_wallace._4844_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5750_  (.A(\u_cpu.ALU.u_wallace._1410_ ),
    .B(\u_cpu.ALU.u_wallace._4609_ ),
    .Y(\u_cpu.ALU.u_wallace._4845_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._5751_  (.A1(\u_cpu.ALU.u_wallace._2933_ ),
    .A2(\u_cpu.ALU.u_wallace._1421_ ),
    .A3(\u_cpu.ALU.u_wallace._4717_ ),
    .A4(\u_cpu.ALU.u_wallace._4599_ ),
    .B1(\u_cpu.ALU.u_wallace._4845_ ),
    .X(\u_cpu.ALU.u_wallace._4846_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5752_  (.A(\u_cpu.ALU.SrcB[8] ),
    .X(\u_cpu.ALU.u_wallace._4847_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5753_  (.A(\u_cpu.ALU.SrcB[9] ),
    .X(\u_cpu.ALU.u_wallace._4848_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5754_  (.A1(\u_cpu.ALU.u_wallace._4556_ ),
    .A2(\u_cpu.ALU.u_wallace._4847_ ),
    .B1(\u_cpu.ALU.u_wallace._4848_ ),
    .B2(\u_cpu.ALU.u_wallace._0600_ ),
    .Y(\u_cpu.ALU.u_wallace._4849_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5755_  (.A1(\u_cpu.ALU.u_wallace._4718_ ),
    .A2(\u_cpu.ALU.u_wallace._4721_ ),
    .B1(\u_cpu.ALU.u_wallace._4728_ ),
    .Y(\u_cpu.ALU.u_wallace._4850_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5756_  (.A(\u_cpu.ALU.u_wallace._1267_ ),
    .B(\u_cpu.ALU.u_wallace._1278_ ),
    .C(\u_cpu.ALU.u_wallace._4720_ ),
    .D(\u_cpu.ALU.u_wallace._4848_ ),
    .X(\u_cpu.ALU.u_wallace._4851_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5757_  (.A1(\u_cpu.ALU.u_wallace._0403_ ),
    .A2(\u_cpu.ALU.u_wallace._4602_ ),
    .B1(\u_cpu.ALU.u_wallace._4849_ ),
    .B2(\u_cpu.ALU.u_wallace._4851_ ),
    .Y(\u_cpu.ALU.u_wallace._4852_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5758_  (.A1(\u_cpu.ALU.u_wallace._4846_ ),
    .A2(\u_cpu.ALU.u_wallace._4849_ ),
    .B1(\u_cpu.ALU.u_wallace._4850_ ),
    .C1(\u_cpu.ALU.u_wallace._4852_ ),
    .Y(\u_cpu.ALU.u_wallace._4853_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5759_  (.A(\u_cpu.ALU.u_wallace._1180_ ),
    .B(\u_cpu.ALU.u_wallace._1191_ ),
    .C(\u_cpu.ALU.u_wallace._4594_ ),
    .D(\u_cpu.ALU.u_wallace._4595_ ),
    .Y(\u_cpu.ALU.u_wallace._4854_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._5760_  (.A_N(\u_cpu.ALU.u_wallace._4849_ ),
    .B(\u_cpu.ALU.u_wallace._4854_ ),
    .C(\u_cpu.ALU.u_wallace._4545_ ),
    .D(\u_cpu.ALU.u_wallace._4610_ ),
    .Y(\u_cpu.ALU.u_wallace._4855_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5761_  (.A1(\u_cpu.ALU.u_wallace._4852_ ),
    .A2(\u_cpu.ALU.u_wallace._4855_ ),
    .B1(\u_cpu.ALU.u_wallace._4850_ ),
    .X(\u_cpu.ALU.u_wallace._4856_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._5762_  (.A_N(\u_cpu.ALU.u_wallace._4844_ ),
    .B(\u_cpu.ALU.u_wallace._4853_ ),
    .C(\u_cpu.ALU.u_wallace._4856_ ),
    .Y(\u_cpu.ALU.u_wallace._4857_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5763_  (.A1(\u_cpu.ALU.u_wallace._4846_ ),
    .A2(\u_cpu.ALU.u_wallace._4849_ ),
    .B1(\u_cpu.ALU.u_wallace._4850_ ),
    .C1(\u_cpu.ALU.u_wallace._4852_ ),
    .X(\u_cpu.ALU.u_wallace._4858_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5764_  (.A1(\u_cpu.ALU.u_wallace._4852_ ),
    .A2(\u_cpu.ALU.u_wallace._4855_ ),
    .B1(\u_cpu.ALU.u_wallace._4850_ ),
    .Y(\u_cpu.ALU.u_wallace._4859_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5765_  (.A1(\u_cpu.ALU.u_wallace._4839_ ),
    .A2(\u_cpu.ALU.u_wallace._4843_ ),
    .B1(\u_cpu.ALU.u_wallace._4858_ ),
    .B2(\u_cpu.ALU.u_wallace._4859_ ),
    .Y(\u_cpu.ALU.u_wallace._4860_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5766_  (.A(\u_cpu.ALU.u_wallace._4835_ ),
    .B(\u_cpu.ALU.u_wallace._4857_ ),
    .C(\u_cpu.ALU.u_wallace._4860_ ),
    .X(\u_cpu.ALU.u_wallace._4861_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._5767_  (.A1(\u_cpu.ALU.u_wallace._4730_ ),
    .A2(\u_cpu.ALU.u_wallace._4733_ ),
    .A3(\u_cpu.ALU.u_wallace._3996_ ),
    .B1(\u_cpu.ALU.u_wallace._4727_ ),
    .X(\u_cpu.ALU.u_wallace._4862_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._5768_  (.A1(\u_cpu.ALU.u_wallace._4692_ ),
    .A2(\u_cpu.ALU.u_wallace._4687_ ),
    .B1(\u_cpu.ALU.u_wallace._4701_ ),
    .B2(\u_cpu.ALU.u_wallace._4700_ ),
    .X(\u_cpu.ALU.u_wallace._4863_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._5769_  (.A1(\u_cpu.ALU.u_wallace._4858_ ),
    .A2(\u_cpu.ALU.u_wallace._4859_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4844_ ),
    .Y(\u_cpu.ALU.u_wallace._4864_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5770_  (.A1(\u_cpu.ALU.u_wallace._4839_ ),
    .A2(\u_cpu.ALU.u_wallace._4843_ ),
    .B1(\u_cpu.ALU.u_wallace._4853_ ),
    .C1(\u_cpu.ALU.u_wallace._4856_ ),
    .Y(\u_cpu.ALU.u_wallace._4865_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5771_  (.A(\u_cpu.ALU.u_wallace._4863_ ),
    .B(\u_cpu.ALU.u_wallace._4864_ ),
    .C(\u_cpu.ALU.u_wallace._4865_ ),
    .Y(\u_cpu.ALU.u_wallace._4866_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5772_  (.A(\u_cpu.ALU.u_wallace._4862_ ),
    .B(\u_cpu.ALU.u_wallace._4866_ ),
    .Y(\u_cpu.ALU.u_wallace._4867_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5773_  (.A(\u_cpu.ALU.u_wallace._4835_ ),
    .B(\u_cpu.ALU.u_wallace._4857_ ),
    .C(\u_cpu.ALU.u_wallace._4860_ ),
    .Y(\u_cpu.ALU.u_wallace._4868_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5774_  (.A1(\u_cpu.ALU.u_wallace._4866_ ),
    .A2(\u_cpu.ALU.u_wallace._4868_ ),
    .B1(\u_cpu.ALU.u_wallace._4862_ ),
    .X(\u_cpu.ALU.u_wallace._4869_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5775_  (.A1(\u_cpu.ALU.u_wallace._4861_ ),
    .A2(\u_cpu.ALU.u_wallace._4867_ ),
    .B1(\u_cpu.ALU.u_wallace._4869_ ),
    .Y(\u_cpu.ALU.u_wallace._4870_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5776_  (.A1(\u_cpu.ALU.u_wallace._4832_ ),
    .A2(\u_cpu.ALU.u_wallace._4834_ ),
    .B1(\u_cpu.ALU.u_wallace._4870_ ),
    .Y(\u_cpu.ALU.u_wallace._4871_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5777_  (.A1(\u_cpu.ALU.u_wallace._4773_ ),
    .A2(\u_cpu.ALU.u_wallace._4777_ ),
    .B1(\u_cpu.ALU.u_wallace._4826_ ),
    .C1(\u_cpu.ALU.u_wallace._4831_ ),
    .Y(\u_cpu.ALU.u_wallace._4872_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._5778_  (.A1(\u_cpu.ALU.u_wallace._4826_ ),
    .A2(\u_cpu.ALU.u_wallace._4831_ ),
    .B1(\u_cpu.ALU.u_wallace._4773_ ),
    .C1(\u_cpu.ALU.u_wallace._4777_ ),
    .X(\u_cpu.ALU.u_wallace._4873_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._5779_  (.A1(\u_cpu.ALU.u_wallace._4867_ ),
    .A2(\u_cpu.ALU.u_wallace._4861_ ),
    .B1(\u_cpu.ALU.u_wallace._4869_ ),
    .C1(\u_cpu.ALU.u_wallace._4872_ ),
    .D1(\u_cpu.ALU.u_wallace._4873_ ),
    .Y(\u_cpu.ALU.u_wallace._4874_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5780_  (.A1(\u_cpu.ALU.u_wallace._4771_ ),
    .A2(\u_cpu.ALU.u_wallace._4772_ ),
    .B1(\u_cpu.ALU.u_wallace._4871_ ),
    .C1(\u_cpu.ALU.u_wallace._4874_ ),
    .Y(\u_cpu.ALU.u_wallace._4875_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._5781_  (.A1(\u_cpu.ALU.u_wallace._4715_ ),
    .A2(\u_cpu.ALU.u_wallace._4750_ ),
    .A3(\u_cpu.ALU.u_wallace._4751_ ),
    .B1(\u_cpu.ALU.u_wallace._4771_ ),
    .X(\u_cpu.ALU.u_wallace._4876_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5782_  (.A1(\u_cpu.ALU.u_wallace._4871_ ),
    .A2(\u_cpu.ALU.u_wallace._4874_ ),
    .B1(\u_cpu.ALU.u_wallace._4876_ ),
    .X(\u_cpu.ALU.u_wallace._4877_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._5783_  (.A_N(\u_cpu.ALU.u_wallace._4770_ ),
    .B(\u_cpu.ALU.u_wallace._4875_ ),
    .C(\u_cpu.ALU.u_wallace._4877_ ),
    .Y(\u_cpu.ALU.u_wallace._4878_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5784_  (.A1(\u_cpu.ALU.u_wallace._4771_ ),
    .A2(\u_cpu.ALU.u_wallace._4772_ ),
    .B1(\u_cpu.ALU.u_wallace._4871_ ),
    .C1(\u_cpu.ALU.u_wallace._4874_ ),
    .X(\u_cpu.ALU.u_wallace._4879_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5785_  (.A1(\u_cpu.ALU.u_wallace._4871_ ),
    .A2(\u_cpu.ALU.u_wallace._4874_ ),
    .B1(\u_cpu.ALU.u_wallace._4876_ ),
    .Y(\u_cpu.ALU.u_wallace._4880_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5786_  (.A1(\u_cpu.ALU.u_wallace._4879_ ),
    .A2(\u_cpu.ALU.u_wallace._4880_ ),
    .B1(\u_cpu.ALU.u_wallace._4770_ ),
    .Y(\u_cpu.ALU.u_wallace._4881_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5787_  (.A(\u_cpu.ALU.u_wallace._4769_ ),
    .B(\u_cpu.ALU.u_wallace._4878_ ),
    .C(\u_cpu.ALU.u_wallace._4881_ ),
    .Y(\u_cpu.ALU.u_wallace._4882_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5788_  (.A1(\u_cpu.ALU.u_wallace._4878_ ),
    .A2(\u_cpu.ALU.u_wallace._4881_ ),
    .B1(\u_cpu.ALU.u_wallace._4769_ ),
    .X(\u_cpu.ALU.u_wallace._4883_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._5789_  (.A1(\u_cpu.ALU.u_wallace._4633_ ),
    .A2(\u_cpu.ALU.u_wallace._4768_ ),
    .B1(\u_cpu.ALU.u_wallace._4882_ ),
    .C1(\u_cpu.ALU.u_wallace._4883_ ),
    .D1(\u_cpu.ALU.u_wallace._4758_ ),
    .Y(\u_cpu.ALU.u_wallace._4884_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5790_  (.A(\u_cpu.ALU.u_wallace._4769_ ),
    .B(\u_cpu.ALU.u_wallace._4878_ ),
    .C(\u_cpu.ALU.u_wallace._4881_ ),
    .X(\u_cpu.ALU.u_wallace._4885_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5791_  (.A1(\u_cpu.ALU.u_wallace._4878_ ),
    .A2(\u_cpu.ALU.u_wallace._4881_ ),
    .B1(\u_cpu.ALU.u_wallace._4769_ ),
    .Y(\u_cpu.ALU.u_wallace._4886_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5792_  (.A1(\u_cpu.ALU.u_wallace._4633_ ),
    .A2(\u_cpu.ALU.u_wallace._4768_ ),
    .B1(\u_cpu.ALU.u_wallace._4758_ ),
    .Y(\u_cpu.ALU.u_wallace._4887_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5793_  (.A1(\u_cpu.ALU.u_wallace._4885_ ),
    .A2(\u_cpu.ALU.u_wallace._4886_ ),
    .B1(\u_cpu.ALU.u_wallace._4887_ ),
    .Y(\u_cpu.ALU.u_wallace._4888_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5794_  (.A(\u_cpu.ALU.u_wallace._4635_ ),
    .B(\u_cpu.ALU.u_wallace._4758_ ),
    .C(\u_cpu.ALU.u_wallace._4759_ ),
    .Y(\u_cpu.ALU.u_wallace._4889_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5795_  (.A1(\u_cpu.ALU.u_wallace._4884_ ),
    .A2(\u_cpu.ALU.u_wallace._4888_ ),
    .B1(\u_cpu.ALU.u_wallace._4889_ ),
    .Y(\u_cpu.ALU.u_wallace._4890_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5796_  (.A(\u_cpu.ALU.u_wallace._4640_ ),
    .B(\u_cpu.ALU.u_wallace._4756_ ),
    .C(\u_cpu.ALU.u_wallace._4757_ ),
    .X(\u_cpu.ALU.u_wallace._4891_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU.u_wallace._5797_  (.A1(\u_cpu.ALU.u_wallace._4891_ ),
    .A2(\u_cpu.ALU.u_wallace._4768_ ),
    .A3(\u_cpu.ALU.u_wallace._4761_ ),
    .B1(\u_cpu.ALU.u_wallace._4884_ ),
    .C1(\u_cpu.ALU.u_wallace._4888_ ),
    .X(\u_cpu.ALU.u_wallace._4892_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5798_  (.A(\u_cpu.ALU.u_wallace._4890_ ),
    .B(\u_cpu.ALU.u_wallace._4892_ ),
    .Y(\u_cpu.ALU.u_wallace._4893_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._5799_  (.A(\u_cpu.ALU.u_wallace._4766_ ),
    .B(\u_cpu.ALU.u_wallace._4893_ ),
    .X(\u_cpu.ALU.Product_Wallace[12] ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5800_  (.A(\u_cpu.ALU.u_wallace._4838_ ),
    .X(\u_cpu.ALU.u_wallace._4894_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5801_  (.A(\u_cpu.ALU.u_wallace._0129_ ),
    .B(\u_cpu.ALU.u_wallace._0184_ ),
    .C(\u_cpu.ALU.u_wallace._4733_ ),
    .D(\u_cpu.ALU.u_wallace._4894_ ),
    .Y(\u_cpu.ALU.u_wallace._4895_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5802_  (.A1(\u_cpu.ALU.u_wallace._4868_ ),
    .A2(\u_cpu.ALU.u_wallace._4867_ ),
    .B1(\u_cpu.ALU.u_wallace._4895_ ),
    .Y(\u_cpu.ALU.u_wallace._4896_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5803_  (.A(\u_cpu.ALU.u_wallace._4895_ ),
    .B(\u_cpu.ALU.u_wallace._4868_ ),
    .C(\u_cpu.ALU.u_wallace._4867_ ),
    .X(\u_cpu.ALU.u_wallace._4897_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._5804_  (.A(\u_cpu.ALU.u_wallace._4654_ ),
    .B(\u_cpu.ALU.u_wallace._4786_ ),
    .C(\u_cpu.ALU.u_wallace._4791_ ),
    .Y(\u_cpu.ALU.u_wallace._4898_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._5805_  (.A1(\u_cpu.ALU.u_wallace._4782_ ),
    .A2(\u_cpu.ALU.u_wallace._4784_ ),
    .A3(\u_cpu.ALU.u_wallace._4792_ ),
    .B1(\u_cpu.ALU.u_wallace._4898_ ),
    .X(\u_cpu.ALU.u_wallace._4899_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5806_  (.A(\u_cpu.ALU.SrcA[12] ),
    .X(\u_cpu.ALU.u_wallace._4900_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5807_  (.A1(\u_cpu.ALU.u_wallace._1914_ ),
    .A2(\u_cpu.ALU.u_wallace._4797_ ),
    .B1(\u_cpu.ALU.u_wallace._4900_ ),
    .B2(\u_cpu.ALU.u_wallace._0479_ ),
    .Y(\u_cpu.ALU.u_wallace._4901_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5808_  (.A(\u_cpu.ALU.u_wallace._0523_ ),
    .B(\u_cpu.ALU.u_wallace._0545_ ),
    .C(\u_cpu.ALU.u_wallace._4653_ ),
    .D(\u_cpu.ALU.u_wallace._4787_ ),
    .Y(\u_cpu.ALU.u_wallace._4902_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._5809_  (.A_N(\u_cpu.ALU.u_wallace._4901_ ),
    .B(\u_cpu.ALU.u_wallace._4902_ ),
    .C(\u_cpu.ALU.u_wallace._4662_ ),
    .D(\u_cpu.ALU.u_wallace._4643_ ),
    .Y(\u_cpu.ALU.u_wallace._4903_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._5810_  (.A(\u_cpu.ALU.u_wallace._4557_ ),
    .Y(\u_cpu.ALU.u_wallace._4904_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5811_  (.A(\u_cpu.ALU.u_wallace._1903_ ),
    .B(\u_cpu.ALU.u_wallace._0807_ ),
    .C(\u_cpu.ALU.u_wallace._4650_ ),
    .D(\u_cpu.ALU.u_wallace._4790_ ),
    .X(\u_cpu.ALU.u_wallace._4905_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5812_  (.A1(\u_cpu.ALU.u_wallace._1224_ ),
    .A2(\u_cpu.ALU.u_wallace._4904_ ),
    .B1(\u_cpu.ALU.u_wallace._4901_ ),
    .B2(\u_cpu.ALU.u_wallace._4905_ ),
    .Y(\u_cpu.ALU.u_wallace._4906_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5813_  (.A(\u_cpu.ALU.SrcA[13] ),
    .X(\u_cpu.ALU.u_wallace._4907_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5814_  (.A1(\u_cpu.ALU.u_wallace._4645_ ),
    .A2(\u_cpu.ALU.u_wallace._4447_ ),
    .B1(\u_cpu.ALU.u_wallace._4907_ ),
    .B2(\u_cpu.ALU.u_wallace._0075_ ),
    .Y(\u_cpu.ALU.u_wallace._4908_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5815_  (.A(\u_cpu.ALU.SrcA[13] ),
    .X(\u_cpu.ALU.u_wallace._4909_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5816_  (.A(\u_cpu.ALU.u_wallace._2747_ ),
    .B(\u_cpu.ALU.u_wallace._2856_ ),
    .C(\u_cpu.ALU.u_wallace._2790_ ),
    .D(\u_cpu.ALU.u_wallace._4909_ ),
    .X(\u_cpu.ALU.u_wallace._4910_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._5817_  (.A(\u_cpu.ALU.u_wallace._4788_ ),
    .B(\u_cpu.ALU.u_wallace._4908_ ),
    .C(\u_cpu.ALU.u_wallace._4910_ ),
    .Y(\u_cpu.ALU.u_wallace._4911_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._5818_  (.A(\u_cpu.ALU.u_wallace._4900_ ),
    .Y(\u_cpu.ALU.u_wallace._4913_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5819_  (.A(\u_cpu.ALU.u_wallace._1826_ ),
    .B(\u_cpu.ALU.u_wallace._3832_ ),
    .Y(\u_cpu.ALU.u_wallace._4914_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.ALU.u_wallace._5820_  (.A1(\u_cpu.ALU.u_wallace._4923_ ),
    .A2(\u_cpu.ALU.u_wallace._4913_ ),
    .A3(\u_cpu.ALU.u_wallace._4914_ ),
    .B1(\u_cpu.ALU.u_wallace._4908_ ),
    .B2(\u_cpu.ALU.u_wallace._4910_ ),
    .X(\u_cpu.ALU.u_wallace._4915_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5821_  (.A1_N(\u_cpu.ALU.u_wallace._4903_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4906_ ),
    .B1(\u_cpu.ALU.u_wallace._4911_ ),
    .B2(\u_cpu.ALU.u_wallace._4915_ ),
    .Y(\u_cpu.ALU.u_wallace._4916_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5822_  (.A(\u_cpu.ALU.u_wallace._4790_ ),
    .X(\u_cpu.ALU.u_wallace._4917_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5823_  (.A(\u_cpu.ALU.u_wallace._0457_ ),
    .B(\u_cpu.ALU.u_wallace._4551_ ),
    .Y(\u_cpu.ALU.u_wallace._4918_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._5824_  (.A1(\u_cpu.ALU.u_wallace._0217_ ),
    .A2(\u_cpu.ALU.u_wallace._4796_ ),
    .A3(\u_cpu.ALU.u_wallace._4794_ ),
    .A4(\u_cpu.ALU.u_wallace._4917_ ),
    .B1(\u_cpu.ALU.u_wallace._4918_ ),
    .X(\u_cpu.ALU.u_wallace._4919_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5825_  (.A(\u_cpu.ALU.SrcA[13] ),
    .X(\u_cpu.ALU.u_wallace._4920_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5826_  (.A(\u_cpu.ALU.u_wallace._4920_ ),
    .X(\u_cpu.ALU.u_wallace._4921_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5827_  (.A(\u_cpu.ALU.u_wallace._1749_ ),
    .B(\u_cpu.ALU.u_wallace._4431_ ),
    .C(\u_cpu.ALU.u_wallace._4450_ ),
    .D(\u_cpu.ALU.u_wallace._4921_ ),
    .Y(\u_cpu.ALU.u_wallace._4922_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._5828_  (.A_N(\u_cpu.ALU.u_wallace._4908_ ),
    .B(\u_cpu.ALU.u_wallace._4922_ ),
    .C(\u_cpu.ALU.u_wallace._4791_ ),
    .Y(\u_cpu.ALU.u_wallace._4924_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5829_  (.A(\u_cpu.ALU.u_wallace._0873_ ),
    .B(\u_cpu.ALU.u_wallace._4917_ ),
    .Y(\u_cpu.ALU.u_wallace._4925_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5830_  (.A1(\u_cpu.ALU.u_wallace._4925_ ),
    .A2(\u_cpu.ALU.u_wallace._4914_ ),
    .B1(\u_cpu.ALU.u_wallace._4908_ ),
    .B2(\u_cpu.ALU.u_wallace._4910_ ),
    .Y(\u_cpu.ALU.u_wallace._4926_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._5831_  (.A1(\u_cpu.ALU.u_wallace._4901_ ),
    .A2(\u_cpu.ALU.u_wallace._4919_ ),
    .B1(\u_cpu.ALU.u_wallace._4906_ ),
    .C1(\u_cpu.ALU.u_wallace._4924_ ),
    .D1(\u_cpu.ALU.u_wallace._4926_ ),
    .Y(\u_cpu.ALU.u_wallace._4927_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5832_  (.A(\u_cpu.ALU.u_wallace._4899_ ),
    .B(\u_cpu.ALU.u_wallace._4916_ ),
    .C(\u_cpu.ALU.u_wallace._4927_ ),
    .Y(\u_cpu.ALU.u_wallace._4928_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5833_  (.A1(\u_cpu.ALU.u_wallace._4903_ ),
    .A2(\u_cpu.ALU.u_wallace._4906_ ),
    .B1(\u_cpu.ALU.u_wallace._4924_ ),
    .B2(\u_cpu.ALU.u_wallace._4926_ ),
    .Y(\u_cpu.ALU.u_wallace._4929_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._5834_  (.A1(\u_cpu.ALU.u_wallace._4901_ ),
    .A2(\u_cpu.ALU.u_wallace._4919_ ),
    .B1(\u_cpu.ALU.u_wallace._4906_ ),
    .C1(\u_cpu.ALU.u_wallace._4924_ ),
    .D1(\u_cpu.ALU.u_wallace._4926_ ),
    .X(\u_cpu.ALU.u_wallace._4930_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._5835_  (.A1(\u_cpu.ALU.u_wallace._4782_ ),
    .A2(\u_cpu.ALU.u_wallace._4784_ ),
    .A3(\u_cpu.ALU.u_wallace._4792_ ),
    .B1(\u_cpu.ALU.u_wallace._4898_ ),
    .Y(\u_cpu.ALU.u_wallace._4931_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5836_  (.A1(\u_cpu.ALU.u_wallace._4929_ ),
    .A2(\u_cpu.ALU.u_wallace._4930_ ),
    .B1(\u_cpu.ALU.u_wallace._4931_ ),
    .Y(\u_cpu.ALU.u_wallace._4932_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._5837_  (.A1(\u_cpu.ALU.u_wallace._4813_ ),
    .A2(\u_cpu.ALU.u_wallace._4539_ ),
    .A3(\u_cpu.ALU.u_wallace._4814_ ),
    .B1(\u_cpu.ALU.u_wallace._4810_ ),
    .X(\u_cpu.ALU.u_wallace._4933_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5838_  (.A(\u_cpu.ALU.u_wallace._0217_ ),
    .B(\u_cpu.ALU.u_wallace._4796_ ),
    .C(\u_cpu.ALU.u_wallace._4554_ ),
    .D(\u_cpu.ALU.u_wallace._4794_ ),
    .X(\u_cpu.ALU.u_wallace._0000_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5839_  (.A(\u_cpu.ALU.u_wallace._4799_ ),
    .B(\u_cpu.ALU.u_wallace._4795_ ),
    .Y(\u_cpu.ALU.u_wallace._0001_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5840_  (.A1(\u_cpu.ALU.u_wallace._4561_ ),
    .A2(\u_cpu.ALU.u_wallace._1497_ ),
    .B1(\u_cpu.ALU.u_wallace._4412_ ),
    .B2(\u_cpu.ALU.u_wallace._4467_ ),
    .X(\u_cpu.ALU.u_wallace._0002_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5841_  (.A(\u_cpu.ALU.u_wallace._4449_ ),
    .B(\u_cpu.ALU.u_wallace._2571_ ),
    .C(\u_cpu.ALU.u_wallace._2582_ ),
    .D(\u_cpu.ALU.u_wallace._4439_ ),
    .Y(\u_cpu.ALU.u_wallace._0003_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5842_  (.A(\u_cpu.ALU.u_wallace._0002_ ),
    .B(\u_cpu.ALU.u_wallace._0003_ ),
    .C(\u_cpu.ALU.u_wallace._4452_ ),
    .D(\u_cpu.ALU.u_wallace._2626_ ),
    .Y(\u_cpu.ALU.u_wallace._0004_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5843_  (.A1(\u_cpu.ALU.u_wallace._3623_ ),
    .A2(\u_cpu.ALU.u_wallace._2078_ ),
    .B1(\u_cpu.ALU.u_wallace._4439_ ),
    .B2(\u_cpu.ALU.u_wallace._2045_ ),
    .Y(\u_cpu.ALU.u_wallace._0005_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5844_  (.A(\u_cpu.ALU.u_wallace._3689_ ),
    .B(\u_cpu.ALU.u_wallace._1465_ ),
    .C(\u_cpu.ALU.u_wallace._2538_ ),
    .D(\u_cpu.ALU.u_wallace._4562_ ),
    .X(\u_cpu.ALU.u_wallace._0006_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5845_  (.A1(\u_cpu.ALU.u_wallace._4454_ ),
    .A2(\u_cpu.ALU.u_wallace._4471_ ),
    .B1(\u_cpu.ALU.u_wallace._0005_ ),
    .B2(\u_cpu.ALU.u_wallace._0006_ ),
    .Y(\u_cpu.ALU.u_wallace._0007_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5846_  (.A1(\u_cpu.ALU.u_wallace._0000_ ),
    .A2(\u_cpu.ALU.u_wallace._0001_ ),
    .B1(\u_cpu.ALU.u_wallace._0004_ ),
    .C1(\u_cpu.ALU.u_wallace._0007_ ),
    .X(\u_cpu.ALU.u_wallace._0008_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5847_  (.A1(\u_cpu.ALU.u_wallace._4799_ ),
    .A2(\u_cpu.ALU.u_wallace._4795_ ),
    .B1(\u_cpu.ALU.u_wallace._4780_ ),
    .Y(\u_cpu.ALU.u_wallace._0009_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5848_  (.A1(\u_cpu.ALU.u_wallace._0004_ ),
    .A2(\u_cpu.ALU.u_wallace._0007_ ),
    .B1(\u_cpu.ALU.u_wallace._0009_ ),
    .Y(\u_cpu.ALU.u_wallace._0011_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._5849_  (.A(\u_cpu.ALU.u_wallace._4933_ ),
    .B(\u_cpu.ALU.u_wallace._0008_ ),
    .C(\u_cpu.ALU.u_wallace._0011_ ),
    .Y(\u_cpu.ALU.u_wallace._0012_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5850_  (.A1(\u_cpu.ALU.u_wallace._0000_ ),
    .A2(\u_cpu.ALU.u_wallace._0001_ ),
    .B1(\u_cpu.ALU.u_wallace._0004_ ),
    .C1(\u_cpu.ALU.u_wallace._0007_ ),
    .Y(\u_cpu.ALU.u_wallace._0013_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5851_  (.A1(\u_cpu.ALU.u_wallace._0004_ ),
    .A2(\u_cpu.ALU.u_wallace._0007_ ),
    .B1(\u_cpu.ALU.u_wallace._0009_ ),
    .X(\u_cpu.ALU.u_wallace._0014_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5852_  (.A(\u_cpu.ALU.u_wallace._2604_ ),
    .X(\u_cpu.ALU.u_wallace._0015_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._5853_  (.A1(\u_cpu.ALU.u_wallace._4809_ ),
    .A2(\u_cpu.ALU.u_wallace._0015_ ),
    .A3(\u_cpu.ALU.u_wallace._1333_ ),
    .B1(\u_cpu.ALU.u_wallace._4815_ ),
    .X(\u_cpu.ALU.u_wallace._0016_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5854_  (.A1(\u_cpu.ALU.u_wallace._0013_ ),
    .A2(\u_cpu.ALU.u_wallace._0014_ ),
    .B1(\u_cpu.ALU.u_wallace._0016_ ),
    .Y(\u_cpu.ALU.u_wallace._0017_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._5855_  (.A1_N(\u_cpu.ALU.u_wallace._4928_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4932_ ),
    .B1(\u_cpu.ALU.u_wallace._0012_ ),
    .B2(\u_cpu.ALU.u_wallace._0017_ ),
    .Y(\u_cpu.ALU.u_wallace._0018_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5856_  (.A(\u_cpu.ALU.u_wallace._0016_ ),
    .B(\u_cpu.ALU.u_wallace._0013_ ),
    .C(\u_cpu.ALU.u_wallace._0014_ ),
    .Y(\u_cpu.ALU.u_wallace._0019_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5857_  (.A1(\u_cpu.ALU.u_wallace._0008_ ),
    .A2(\u_cpu.ALU.u_wallace._0011_ ),
    .B1(\u_cpu.ALU.u_wallace._4933_ ),
    .Y(\u_cpu.ALU.u_wallace._0020_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5858_  (.A(\u_cpu.ALU.u_wallace._4928_ ),
    .B(\u_cpu.ALU.u_wallace._4932_ ),
    .C(\u_cpu.ALU.u_wallace._0019_ ),
    .D(\u_cpu.ALU.u_wallace._0020_ ),
    .Y(\u_cpu.ALU.u_wallace._0022_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU.u_wallace._5859_  (.A1(\u_cpu.ALU.u_wallace._4655_ ),
    .A2(\u_cpu.ALU.u_wallace._4778_ ),
    .B1(\u_cpu.ALU.u_wallace._4803_ ),
    .C1(\u_cpu.ALU.u_wallace._4804_ ),
    .Y(\u_cpu.ALU.u_wallace._0023_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._5860_  (.A1(\u_cpu.ALU.u_wallace._4806_ ),
    .A2(\u_cpu.ALU.u_wallace._4828_ ),
    .A3(\u_cpu.ALU.u_wallace._4830_ ),
    .B1(\u_cpu.ALU.u_wallace._0023_ ),
    .X(\u_cpu.ALU.u_wallace._0024_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5861_  (.A1(\u_cpu.ALU.u_wallace._0018_ ),
    .A2(\u_cpu.ALU.u_wallace._0022_ ),
    .B1(\u_cpu.ALU.u_wallace._0024_ ),
    .Y(\u_cpu.ALU.u_wallace._0025_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._5862_  (.A1(\u_cpu.ALU.u_wallace._4665_ ),
    .A2(\u_cpu.ALU.u_wallace._4818_ ),
    .B1(\u_cpu.ALU.u_wallace._4816_ ),
    .X(\u_cpu.ALU.u_wallace._0026_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5863_  (.A1(\u_cpu.ALU.u_wallace._4811_ ),
    .A2(\u_cpu.ALU.u_wallace._0026_ ),
    .B1(\u_cpu.ALU.u_wallace._4823_ ),
    .B2(\u_cpu.ALU.u_wallace._4824_ ),
    .Y(\u_cpu.ALU.u_wallace._0027_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5864_  (.A(\u_cpu.ALU.SrcB[11] ),
    .X(\u_cpu.ALU.u_wallace._0028_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5865_  (.A(\u_cpu.ALU.SrcB[12] ),
    .X(\u_cpu.ALU.u_wallace._0029_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5866_  (.A(\u_cpu.ALU.u_wallace._0512_ ),
    .B(\u_cpu.ALU.u_wallace._0250_ ),
    .C(\u_cpu.ALU.u_wallace._0028_ ),
    .D(\u_cpu.ALU.u_wallace._0029_ ),
    .X(\u_cpu.ALU.u_wallace._0030_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5867_  (.A1(\u_cpu.ALU.u_wallace._4597_ ),
    .A2(\u_cpu.ALU.u_wallace._4840_ ),
    .B1(\u_cpu.ALU.u_wallace._4842_ ),
    .B2(\u_cpu.ALU.u_wallace._1454_ ),
    .Y(\u_cpu.ALU.u_wallace._0031_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5868_  (.A(\u_cpu.ALU.SrcB[13] ),
    .X(\u_cpu.ALU.u_wallace._0033_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5869_  (.A(\u_cpu.ALU.u_wallace._0033_ ),
    .X(\u_cpu.ALU.u_wallace._0034_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5870_  (.A1(\u_cpu.ALU.u_wallace._0030_ ),
    .A2(\u_cpu.ALU.u_wallace._0031_ ),
    .B1(\u_cpu.ALU.u_wallace._0108_ ),
    .C1(\u_cpu.ALU.u_wallace._0034_ ),
    .X(\u_cpu.ALU.u_wallace._0035_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._5871_  (.A(\u_cpu.ALU.SrcB[13] ),
    .Y(\u_cpu.ALU.u_wallace._0036_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5872_  (.A(\u_cpu.ALU.u_wallace._0036_ ),
    .X(\u_cpu.ALU.u_wallace._0037_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5873_  (.A(\u_cpu.ALU.u_wallace._4597_ ),
    .B(\u_cpu.ALU.u_wallace._0151_ ),
    .C(\u_cpu.ALU.u_wallace._4840_ ),
    .D(\u_cpu.ALU.u_wallace._4842_ ),
    .Y(\u_cpu.ALU.u_wallace._0038_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5874_  (.A1(\u_cpu.ALU.u_wallace._1410_ ),
    .A2(\u_cpu.ALU.u_wallace._4837_ ),
    .B1(\u_cpu.ALU.u_wallace._4838_ ),
    .B2(\u_cpu.ALU.u_wallace._0731_ ),
    .X(\u_cpu.ALU.u_wallace._0039_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5875_  (.A1(\u_cpu.ALU.u_wallace._0032_ ),
    .A2(\u_cpu.ALU.u_wallace._0037_ ),
    .B1(\u_cpu.ALU.u_wallace._0038_ ),
    .C1(\u_cpu.ALU.u_wallace._0039_ ),
    .X(\u_cpu.ALU.u_wallace._0040_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5876_  (.A(\u_cpu.ALU.SrcB[10] ),
    .X(\u_cpu.ALU.u_wallace._0041_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5877_  (.A(\u_cpu.ALU.u_wallace._1278_ ),
    .B(\u_cpu.ALU.u_wallace._0041_ ),
    .Y(\u_cpu.ALU.u_wallace._0042_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._5878_  (.A1(\u_cpu.ALU.u_wallace._4529_ ),
    .A2(\u_cpu.ALU.u_wallace._0906_ ),
    .A3(\u_cpu.ALU.u_wallace._4018_ ),
    .A4(\u_cpu.ALU.u_wallace._4302_ ),
    .B1(\u_cpu.ALU.u_wallace._0042_ ),
    .X(\u_cpu.ALU.u_wallace._0044_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5879_  (.A(\u_cpu.ALU.SrcB[9] ),
    .X(\u_cpu.ALU.u_wallace._0045_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5880_  (.A1(\u_cpu.ALU.u_wallace._2955_ ),
    .A2(\u_cpu.ALU.u_wallace._4847_ ),
    .B1(\u_cpu.ALU.u_wallace._0045_ ),
    .B2(\u_cpu.ALU.u_wallace._4556_ ),
    .Y(\u_cpu.ALU.u_wallace._0046_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5881_  (.A1(\u_cpu.ALU.u_wallace._4845_ ),
    .A2(\u_cpu.ALU.u_wallace._4849_ ),
    .B1(\u_cpu.ALU.u_wallace._4854_ ),
    .Y(\u_cpu.ALU.u_wallace._0047_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5882_  (.A(\u_cpu.ALU.u_wallace._1311_ ),
    .B(\u_cpu.ALU.u_wallace._4556_ ),
    .C(\u_cpu.ALU.u_wallace._4716_ ),
    .D(\u_cpu.ALU.u_wallace._4598_ ),
    .X(\u_cpu.ALU.u_wallace._0048_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5883_  (.A1(\u_cpu.ALU.u_wallace._0610_ ),
    .A2(\u_cpu.ALU.u_wallace._4601_ ),
    .B1(\u_cpu.ALU.u_wallace._0046_ ),
    .B2(\u_cpu.ALU.u_wallace._0048_ ),
    .Y(\u_cpu.ALU.u_wallace._0049_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5884_  (.A1(\u_cpu.ALU.u_wallace._0044_ ),
    .A2(\u_cpu.ALU.u_wallace._0046_ ),
    .B1(\u_cpu.ALU.u_wallace._0047_ ),
    .C1(\u_cpu.ALU.u_wallace._0049_ ),
    .X(\u_cpu.ALU.u_wallace._0050_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5885_  (.A(\u_cpu.ALU.u_wallace._4529_ ),
    .B(\u_cpu.ALU.u_wallace._1180_ ),
    .C(\u_cpu.ALU.u_wallace._4594_ ),
    .D(\u_cpu.ALU.u_wallace._4302_ ),
    .Y(\u_cpu.ALU.u_wallace._0051_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5886_  (.A(\u_cpu.ALU.u_wallace._0041_ ),
    .X(\u_cpu.ALU.u_wallace._0052_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._5887_  (.A_N(\u_cpu.ALU.u_wallace._0046_ ),
    .B(\u_cpu.ALU.u_wallace._0051_ ),
    .C(\u_cpu.ALU.u_wallace._4527_ ),
    .D(\u_cpu.ALU.u_wallace._0052_ ),
    .Y(\u_cpu.ALU.u_wallace._0053_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5888_  (.A1(\u_cpu.ALU.u_wallace._0053_ ),
    .A2(\u_cpu.ALU.u_wallace._0049_ ),
    .B1(\u_cpu.ALU.u_wallace._0047_ ),
    .Y(\u_cpu.ALU.u_wallace._0054_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5889_  (.A1(\u_cpu.ALU.u_wallace._0035_ ),
    .A2(\u_cpu.ALU.u_wallace._0040_ ),
    .B1(\u_cpu.ALU.u_wallace._0050_ ),
    .B2(\u_cpu.ALU.u_wallace._0054_ ),
    .Y(\u_cpu.ALU.u_wallace._0055_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._5890_  (.A1(\u_cpu.ALU.u_wallace._0032_ ),
    .A2(\u_cpu.ALU.u_wallace._0037_ ),
    .B1(\u_cpu.ALU.u_wallace._0030_ ),
    .B2(\u_cpu.ALU.u_wallace._0031_ ),
    .X(\u_cpu.ALU.u_wallace._0056_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5891_  (.A(\u_cpu.ALU.u_wallace._0033_ ),
    .X(\u_cpu.ALU.u_wallace._0057_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5892_  (.A(\u_cpu.ALU.u_wallace._0039_ ),
    .B(\u_cpu.ALU.u_wallace._0057_ ),
    .C(\u_cpu.ALU.u_wallace._0994_ ),
    .D(\u_cpu.ALU.u_wallace._0038_ ),
    .X(\u_cpu.ALU.u_wallace._0058_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5893_  (.A1(\u_cpu.ALU.u_wallace._0044_ ),
    .A2(\u_cpu.ALU.u_wallace._0046_ ),
    .B1(\u_cpu.ALU.u_wallace._0047_ ),
    .C1(\u_cpu.ALU.u_wallace._0049_ ),
    .Y(\u_cpu.ALU.u_wallace._0059_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5894_  (.A1(\u_cpu.ALU.u_wallace._0053_ ),
    .A2(\u_cpu.ALU.u_wallace._0049_ ),
    .B1(\u_cpu.ALU.u_wallace._0047_ ),
    .X(\u_cpu.ALU.u_wallace._0060_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5895_  (.A1(\u_cpu.ALU.u_wallace._0056_ ),
    .A2(\u_cpu.ALU.u_wallace._0058_ ),
    .B1(\u_cpu.ALU.u_wallace._0059_ ),
    .C1(\u_cpu.ALU.u_wallace._0060_ ),
    .Y(\u_cpu.ALU.u_wallace._0061_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5896_  (.A(\u_cpu.ALU.u_wallace._0027_ ),
    .B(\u_cpu.ALU.u_wallace._0055_ ),
    .C(\u_cpu.ALU.u_wallace._0061_ ),
    .Y(\u_cpu.ALU.u_wallace._0062_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5897_  (.A1(\u_cpu.ALU.u_wallace._0035_ ),
    .A2(\u_cpu.ALU.u_wallace._0040_ ),
    .B1(\u_cpu.ALU.u_wallace._0059_ ),
    .C1(\u_cpu.ALU.u_wallace._0060_ ),
    .Y(\u_cpu.ALU.u_wallace._0063_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5898_  (.A1(\u_cpu.ALU.u_wallace._0056_ ),
    .A2(\u_cpu.ALU.u_wallace._0058_ ),
    .B1(\u_cpu.ALU.u_wallace._0050_ ),
    .B2(\u_cpu.ALU.u_wallace._0054_ ),
    .Y(\u_cpu.ALU.u_wallace._0065_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5899_  (.A1(\u_cpu.ALU.u_wallace._4819_ ),
    .A2(\u_cpu.ALU.u_wallace._4827_ ),
    .B1(\u_cpu.ALU.u_wallace._0063_ ),
    .C1(\u_cpu.ALU.u_wallace._0065_ ),
    .Y(\u_cpu.ALU.u_wallace._0066_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5900_  (.A(\u_cpu.ALU.u_wallace._4844_ ),
    .B(\u_cpu.ALU.u_wallace._4859_ ),
    .Y(\u_cpu.ALU.u_wallace._0067_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._5901_  (.A1(\u_cpu.ALU.u_wallace._4850_ ),
    .A2(\u_cpu.ALU.u_wallace._4852_ ),
    .A3(\u_cpu.ALU.u_wallace._4855_ ),
    .B1(\u_cpu.ALU.u_wallace._0067_ ),
    .X(\u_cpu.ALU.u_wallace._0068_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5902_  (.A1(\u_cpu.ALU.u_wallace._0062_ ),
    .A2(\u_cpu.ALU.u_wallace._0066_ ),
    .B1(\u_cpu.ALU.u_wallace._0068_ ),
    .X(\u_cpu.ALU.u_wallace._0069_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5903_  (.A1(\u_cpu.ALU.u_wallace._4858_ ),
    .A2(\u_cpu.ALU.u_wallace._0067_ ),
    .B1(\u_cpu.ALU.u_wallace._0062_ ),
    .C1(\u_cpu.ALU.u_wallace._0066_ ),
    .Y(\u_cpu.ALU.u_wallace._0070_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5904_  (.A(\u_cpu.ALU.u_wallace._4899_ ),
    .B(\u_cpu.ALU.u_wallace._4916_ ),
    .C(\u_cpu.ALU.u_wallace._4927_ ),
    .X(\u_cpu.ALU.u_wallace._0071_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5905_  (.A(\u_cpu.ALU.u_wallace._0071_ ),
    .X(\u_cpu.ALU.u_wallace._0072_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5906_  (.A(\u_cpu.ALU.u_wallace._4932_ ),
    .B(\u_cpu.ALU.u_wallace._0019_ ),
    .C(\u_cpu.ALU.u_wallace._0020_ ),
    .Y(\u_cpu.ALU.u_wallace._0073_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5907_  (.A1(\u_cpu.ALU.u_wallace._4819_ ),
    .A2(\u_cpu.ALU.u_wallace._4829_ ),
    .B1(\u_cpu.ALU.u_wallace._4824_ ),
    .Y(\u_cpu.ALU.u_wallace._0074_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._5908_  (.A_N(\u_cpu.ALU.u_wallace._4824_ ),
    .B(\u_cpu.ALU.u_wallace._4821_ ),
    .C(\u_cpu.ALU.u_wallace._4823_ ),
    .Y(\u_cpu.ALU.u_wallace._0076_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5909_  (.A1(\u_cpu.ALU.u_wallace._4793_ ),
    .A2(\u_cpu.ALU.u_wallace._4801_ ),
    .B1(\u_cpu.ALU.u_wallace._4779_ ),
    .Y(\u_cpu.ALU.u_wallace._0077_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5910_  (.A1(\u_cpu.ALU.u_wallace._0074_ ),
    .A2(\u_cpu.ALU.u_wallace._0076_ ),
    .B1(\u_cpu.ALU.u_wallace._0077_ ),
    .Y(\u_cpu.ALU.u_wallace._0078_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._5911_  (.A1(\u_cpu.ALU.u_wallace._0072_ ),
    .A2(\u_cpu.ALU.u_wallace._0073_ ),
    .B1(\u_cpu.ALU.u_wallace._0023_ ),
    .B2(\u_cpu.ALU.u_wallace._0078_ ),
    .C1(\u_cpu.ALU.u_wallace._0018_ ),
    .Y(\u_cpu.ALU.u_wallace._0079_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5912_  (.A(\u_cpu.ALU.u_wallace._0069_ ),
    .B(\u_cpu.ALU.u_wallace._0070_ ),
    .C(\u_cpu.ALU.u_wallace._0079_ ),
    .Y(\u_cpu.ALU.u_wallace._0080_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5913_  (.A1(\u_cpu.ALU.u_wallace._0062_ ),
    .A2(\u_cpu.ALU.u_wallace._0066_ ),
    .B1(\u_cpu.ALU.u_wallace._0068_ ),
    .Y(\u_cpu.ALU.u_wallace._0081_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5914_  (.A1(\u_cpu.ALU.u_wallace._4858_ ),
    .A2(\u_cpu.ALU.u_wallace._0067_ ),
    .B1(\u_cpu.ALU.u_wallace._0062_ ),
    .C1(\u_cpu.ALU.u_wallace._0066_ ),
    .X(\u_cpu.ALU.u_wallace._0082_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._5915_  (.A1(\u_cpu.ALU.u_wallace._0072_ ),
    .A2(\u_cpu.ALU.u_wallace._0073_ ),
    .B1(\u_cpu.ALU.u_wallace._0023_ ),
    .B2(\u_cpu.ALU.u_wallace._0078_ ),
    .C1(\u_cpu.ALU.u_wallace._0018_ ),
    .X(\u_cpu.ALU.u_wallace._0083_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5916_  (.A1(\u_cpu.ALU.u_wallace._0081_ ),
    .A2(\u_cpu.ALU.u_wallace._0082_ ),
    .B1(\u_cpu.ALU.u_wallace._0083_ ),
    .B2(\u_cpu.ALU.u_wallace._0025_ ),
    .Y(\u_cpu.ALU.u_wallace._0084_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5917_  (.A1(\u_cpu.ALU.u_wallace._4834_ ),
    .A2(\u_cpu.ALU.u_wallace._4870_ ),
    .B1(\u_cpu.ALU.u_wallace._4872_ ),
    .Y(\u_cpu.ALU.u_wallace._0085_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5918_  (.A1(\u_cpu.ALU.u_wallace._0025_ ),
    .A2(\u_cpu.ALU.u_wallace._0080_ ),
    .B1(\u_cpu.ALU.u_wallace._0084_ ),
    .C1(\u_cpu.ALU.u_wallace._0085_ ),
    .X(\u_cpu.ALU.u_wallace._0087_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5919_  (.A(\u_cpu.ALU.u_wallace._0081_ ),
    .B(\u_cpu.ALU.u_wallace._0082_ ),
    .Y(\u_cpu.ALU.u_wallace._0088_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5920_  (.A1(\u_cpu.ALU.u_wallace._0018_ ),
    .A2(\u_cpu.ALU.u_wallace._0022_ ),
    .B1(\u_cpu.ALU.u_wallace._0024_ ),
    .X(\u_cpu.ALU.u_wallace._0089_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5921_  (.A(\u_cpu.ALU.u_wallace._0088_ ),
    .B(\u_cpu.ALU.u_wallace._0079_ ),
    .C(\u_cpu.ALU.u_wallace._0089_ ),
    .Y(\u_cpu.ALU.u_wallace._0090_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5922_  (.A1(\u_cpu.ALU.u_wallace._0084_ ),
    .A2(\u_cpu.ALU.u_wallace._0090_ ),
    .B1(\u_cpu.ALU.u_wallace._0085_ ),
    .Y(\u_cpu.ALU.u_wallace._0091_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5923_  (.A1(\u_cpu.ALU.u_wallace._4896_ ),
    .A2(\u_cpu.ALU.u_wallace._4897_ ),
    .B1(\u_cpu.ALU.u_wallace._0087_ ),
    .B2(\u_cpu.ALU.u_wallace._0091_ ),
    .Y(\u_cpu.ALU.u_wallace._0092_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU.u_wallace._5924_  (.A(\u_cpu.ALU.u_wallace._4896_ ),
    .B(\u_cpu.ALU.u_wallace._4897_ ),
    .X(\u_cpu.ALU.u_wallace._0093_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5925_  (.A1(\u_cpu.ALU.u_wallace._0025_ ),
    .A2(\u_cpu.ALU.u_wallace._0080_ ),
    .B1(\u_cpu.ALU.u_wallace._0084_ ),
    .C1(\u_cpu.ALU.u_wallace._0085_ ),
    .Y(\u_cpu.ALU.u_wallace._0094_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5926_  (.A1(\u_cpu.ALU.u_wallace._0084_ ),
    .A2(\u_cpu.ALU.u_wallace._0090_ ),
    .B1(\u_cpu.ALU.u_wallace._0085_ ),
    .X(\u_cpu.ALU.u_wallace._0095_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._5927_  (.A_N(\u_cpu.ALU.u_wallace._0093_ ),
    .B(\u_cpu.ALU.u_wallace._0094_ ),
    .C(\u_cpu.ALU.u_wallace._0095_ ),
    .Y(\u_cpu.ALU.u_wallace._0096_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5928_  (.A1(\u_cpu.ALU.u_wallace._4770_ ),
    .A2(\u_cpu.ALU.u_wallace._4880_ ),
    .B1(\u_cpu.ALU.u_wallace._4875_ ),
    .Y(\u_cpu.ALU.u_wallace._0098_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5929_  (.A1(\u_cpu.ALU.u_wallace._0092_ ),
    .A2(\u_cpu.ALU.u_wallace._0096_ ),
    .B1(\u_cpu.ALU.u_wallace._0098_ ),
    .X(\u_cpu.ALU.u_wallace._0099_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5930_  (.A(\u_cpu.ALU.u_wallace._0092_ ),
    .B(\u_cpu.ALU.u_wallace._0096_ ),
    .C(\u_cpu.ALU.u_wallace._0098_ ),
    .Y(\u_cpu.ALU.u_wallace._0100_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._5931_  (.A1(\u_cpu.ALU.u_wallace._4758_ ),
    .A2(\u_cpu.ALU.u_wallace._4886_ ),
    .B1(\u_cpu.ALU.u_wallace._0099_ ),
    .C1(\u_cpu.ALU.u_wallace._0100_ ),
    .D1(\u_cpu.ALU.u_wallace._4882_ ),
    .X(\u_cpu.ALU.u_wallace._0101_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5932_  (.A(\u_cpu.ALU.u_wallace._4891_ ),
    .B(\u_cpu.ALU.u_wallace._4883_ ),
    .Y(\u_cpu.ALU.u_wallace._0102_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5933_  (.A1(\u_cpu.ALU.u_wallace._0099_ ),
    .A2(\u_cpu.ALU.u_wallace._0100_ ),
    .B1(\u_cpu.ALU.u_wallace._0102_ ),
    .B2(\u_cpu.ALU.u_wallace._4882_ ),
    .Y(\u_cpu.ALU.u_wallace._0103_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5934_  (.A(\u_cpu.ALU.u_wallace._4633_ ),
    .B(\u_cpu.ALU.u_wallace._4768_ ),
    .Y(\u_cpu.ALU.u_wallace._0104_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5935_  (.A(\u_cpu.ALU.u_wallace._0104_ ),
    .B(\u_cpu.ALU.u_wallace._4882_ ),
    .C(\u_cpu.ALU.u_wallace._4883_ ),
    .D(\u_cpu.ALU.u_wallace._4758_ ),
    .Y(\u_cpu.ALU.u_wallace._0105_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._5936_  (.A1(\u_cpu.ALU.u_wallace._0101_ ),
    .A2(\u_cpu.ALU.u_wallace._0103_ ),
    .B1_N(\u_cpu.ALU.u_wallace._0105_ ),
    .Y(\u_cpu.ALU.u_wallace._0106_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5937_  (.A(\u_cpu.ALU.u_wallace._0099_ ),
    .B(\u_cpu.ALU.u_wallace._0100_ ),
    .Y(\u_cpu.ALU.u_wallace._0107_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._5938_  (.A1(\u_cpu.ALU.u_wallace._4891_ ),
    .A2(\u_cpu.ALU.u_wallace._4883_ ),
    .B1(\u_cpu.ALU.u_wallace._4885_ ),
    .C1(\u_cpu.ALU.u_wallace._0107_ ),
    .X(\u_cpu.ALU.u_wallace._0109_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5939_  (.A1(\u_cpu.ALU.u_wallace._0099_ ),
    .A2(\u_cpu.ALU.u_wallace._0100_ ),
    .B1(\u_cpu.ALU.u_wallace._0102_ ),
    .B2(\u_cpu.ALU.u_wallace._4882_ ),
    .X(\u_cpu.ALU.u_wallace._0110_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5940_  (.A(\u_cpu.ALU.u_wallace._0109_ ),
    .B(\u_cpu.ALU.u_wallace._0110_ ),
    .C(\u_cpu.ALU.u_wallace._0105_ ),
    .Y(\u_cpu.ALU.u_wallace._0111_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5941_  (.A(\u_cpu.ALU.u_wallace._0106_ ),
    .B(\u_cpu.ALU.u_wallace._0111_ ),
    .Y(\u_cpu.ALU.u_wallace._0112_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5942_  (.A1(\u_cpu.ALU.u_wallace._4766_ ),
    .A2(\u_cpu.ALU.u_wallace._4893_ ),
    .B1(\u_cpu.ALU.u_wallace._4890_ ),
    .Y(\u_cpu.ALU.u_wallace._0113_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._5943_  (.A(\u_cpu.ALU.u_wallace._0112_ ),
    .B(\u_cpu.ALU.u_wallace._0113_ ),
    .X(\u_cpu.ALU.Product_Wallace[13] ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._5944_  (.A1(\u_cpu.ALU.u_wallace._4769_ ),
    .A2(\u_cpu.ALU.u_wallace._4878_ ),
    .A3(\u_cpu.ALU.u_wallace._4881_ ),
    .B1(\u_cpu.ALU.u_wallace._0102_ ),
    .X(\u_cpu.ALU.u_wallace._0114_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5945_  (.A1(\u_cpu.ALU.u_wallace._0092_ ),
    .A2(\u_cpu.ALU.u_wallace._0096_ ),
    .B1(\u_cpu.ALU.u_wallace._0098_ ),
    .Y(\u_cpu.ALU.u_wallace._0115_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5946_  (.A1(\u_cpu.ALU.u_wallace._0093_ ),
    .A2(\u_cpu.ALU.u_wallace._0091_ ),
    .B1(\u_cpu.ALU.u_wallace._0094_ ),
    .Y(\u_cpu.ALU.u_wallace._0116_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5947_  (.A(\u_cpu.ALU.u_wallace._0057_ ),
    .X(\u_cpu.ALU.u_wallace._0117_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._5948_  (.A1(\u_cpu.ALU.u_wallace._0039_ ),
    .A2(\u_cpu.ALU.u_wallace._0117_ ),
    .A3(\u_cpu.ALU.u_wallace._1070_ ),
    .B1(\u_cpu.ALU.u_wallace._0030_ ),
    .X(\u_cpu.ALU.u_wallace._0119_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5949_  (.A(\u_cpu.ALU.SrcB[14] ),
    .X(\u_cpu.ALU.u_wallace._0120_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5950_  (.A(\u_cpu.ALU.u_wallace._0120_ ),
    .X(\u_cpu.ALU.u_wallace._0121_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5951_  (.A(\u_cpu.ALU.u_wallace._0121_ ),
    .X(\u_cpu.ALU.u_wallace._0122_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5952_  (.A(\u_cpu.ALU.u_wallace._0119_ ),
    .B(\u_cpu.ALU.u_wallace._0122_ ),
    .C(\u_cpu.ALU.u_wallace._3996_ ),
    .X(\u_cpu.ALU.u_wallace._0123_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5953_  (.A(\u_cpu.ALU.u_wallace._0036_ ),
    .X(\u_cpu.ALU.u_wallace._0124_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5954_  (.A(\u_cpu.ALU.u_wallace._0118_ ),
    .B(\u_cpu.ALU.u_wallace._0122_ ),
    .Y(\u_cpu.ALU.u_wallace._0125_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU.u_wallace._5955_  (.A1(\u_cpu.ALU.u_wallace._0043_ ),
    .A2(\u_cpu.ALU.u_wallace._0124_ ),
    .A3(\u_cpu.ALU.u_wallace._0031_ ),
    .B1(\u_cpu.ALU.u_wallace._0125_ ),
    .C1(\u_cpu.ALU.u_wallace._0038_ ),
    .X(\u_cpu.ALU.u_wallace._0126_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU.u_wallace._5956_  (.A(\u_cpu.ALU.u_wallace._0123_ ),
    .B(\u_cpu.ALU.u_wallace._0126_ ),
    .X(\u_cpu.ALU.u_wallace._0127_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5957_  (.A1(\u_cpu.ALU.u_wallace._0066_ ),
    .A2(\u_cpu.ALU.u_wallace._0070_ ),
    .B1(\u_cpu.ALU.u_wallace._0127_ ),
    .Y(\u_cpu.ALU.u_wallace._0128_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5958_  (.A1(\u_cpu.ALU.u_wallace._0123_ ),
    .A2(\u_cpu.ALU.u_wallace._0126_ ),
    .B1(\u_cpu.ALU.u_wallace._0066_ ),
    .C1(\u_cpu.ALU.u_wallace._0070_ ),
    .Y(\u_cpu.ALU.u_wallace._0130_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.ALU.u_wallace._5959_  (.A(\u_cpu.ALU.u_wallace._0128_ ),
    .B_N(\u_cpu.ALU.u_wallace._0130_ ),
    .X(\u_cpu.ALU.u_wallace._0131_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._5960_  (.A1(\u_cpu.ALU.u_wallace._4933_ ),
    .A2(\u_cpu.ALU.u_wallace._0011_ ),
    .B1(\u_cpu.ALU.u_wallace._0013_ ),
    .X(\u_cpu.ALU.u_wallace._0132_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5961_  (.A(\u_cpu.ALU.u_wallace._2922_ ),
    .B(\u_cpu.ALU.u_wallace._0041_ ),
    .Y(\u_cpu.ALU.u_wallace._0133_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._5962_  (.A1(\u_cpu.ALU.u_wallace._4452_ ),
    .A2(\u_cpu.ALU.u_wallace._4529_ ),
    .A3(\u_cpu.ALU.u_wallace._4018_ ),
    .A4(\u_cpu.ALU.u_wallace._4302_ ),
    .B1(\u_cpu.ALU.u_wallace._0133_ ),
    .X(\u_cpu.ALU.u_wallace._0134_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5963_  (.A1(\u_cpu.ALU.u_wallace._1837_ ),
    .A2(\u_cpu.ALU.u_wallace._4007_ ),
    .B1(\u_cpu.ALU.u_wallace._0045_ ),
    .B2(\u_cpu.ALU.u_wallace._1311_ ),
    .Y(\u_cpu.ALU.u_wallace._0135_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5964_  (.A1(\u_cpu.ALU.u_wallace._0042_ ),
    .A2(\u_cpu.ALU.u_wallace._0046_ ),
    .B1(\u_cpu.ALU.u_wallace._0051_ ),
    .Y(\u_cpu.ALU.u_wallace._0136_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5965_  (.A(\u_cpu.ALU.u_wallace._2834_ ),
    .B(\u_cpu.ALU.u_wallace._1311_ ),
    .C(\u_cpu.ALU.u_wallace._4716_ ),
    .D(\u_cpu.ALU.u_wallace._4598_ ),
    .X(\u_cpu.ALU.u_wallace._0137_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5966_  (.A1(\u_cpu.ALU.u_wallace._0135_ ),
    .A2(\u_cpu.ALU.u_wallace._0137_ ),
    .B1(\u_cpu.ALU.u_wallace._0133_ ),
    .Y(\u_cpu.ALU.u_wallace._0138_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._5967_  (.A1(\u_cpu.ALU.u_wallace._0134_ ),
    .A2(\u_cpu.ALU.u_wallace._0135_ ),
    .B1(\u_cpu.ALU.u_wallace._0136_ ),
    .C1(\u_cpu.ALU.u_wallace._0138_ ),
    .X(\u_cpu.ALU.u_wallace._0139_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5968_  (.A(\u_cpu.ALU.u_wallace._3832_ ),
    .B(\u_cpu.ALU.u_wallace._1125_ ),
    .C(\u_cpu.ALU.u_wallace._4594_ ),
    .D(\u_cpu.ALU.u_wallace._4302_ ),
    .Y(\u_cpu.ALU.u_wallace._0141_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._5969_  (.A_N(\u_cpu.ALU.u_wallace._0135_ ),
    .B(\u_cpu.ALU.u_wallace._0141_ ),
    .C(\u_cpu.ALU.u_wallace._2933_ ),
    .D(\u_cpu.ALU.u_wallace._0052_ ),
    .Y(\u_cpu.ALU.u_wallace._0142_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5970_  (.A1(\u_cpu.ALU.u_wallace._0138_ ),
    .A2(\u_cpu.ALU.u_wallace._0142_ ),
    .B1(\u_cpu.ALU.u_wallace._0136_ ),
    .Y(\u_cpu.ALU.u_wallace._0143_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._5971_  (.A(\u_cpu.ALU.SrcB[12] ),
    .X(\u_cpu.ALU.u_wallace._0144_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5972_  (.A1(\u_cpu.ALU.u_wallace._0600_ ),
    .A2(\u_cpu.ALU.u_wallace._4731_ ),
    .B1(\u_cpu.ALU.u_wallace._0144_ ),
    .B2(\u_cpu.ALU.u_wallace._0348_ ),
    .X(\u_cpu.ALU.u_wallace._0145_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5973_  (.A(\u_cpu.ALU.u_wallace._1410_ ),
    .B(\u_cpu.ALU.u_wallace._1191_ ),
    .C(\u_cpu.ALU.u_wallace._4837_ ),
    .D(\u_cpu.ALU.u_wallace._0029_ ),
    .Y(\u_cpu.ALU.u_wallace._0146_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5974_  (.A1(\u_cpu.ALU.u_wallace._4463_ ),
    .A2(\u_cpu.ALU.u_wallace._0057_ ),
    .B1(\u_cpu.ALU.u_wallace._0145_ ),
    .B2(\u_cpu.ALU.u_wallace._0146_ ),
    .Y(\u_cpu.ALU.u_wallace._0147_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5975_  (.A(\u_cpu.ALU.u_wallace._0145_ ),
    .B(\u_cpu.ALU.u_wallace._0146_ ),
    .C(\u_cpu.ALU.u_wallace._0261_ ),
    .D(\u_cpu.ALU.u_wallace._0057_ ),
    .X(\u_cpu.ALU.u_wallace._0148_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._5976_  (.A(\u_cpu.ALU.u_wallace._0147_ ),
    .B(\u_cpu.ALU.u_wallace._0148_ ),
    .Y(\u_cpu.ALU.u_wallace._0149_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5977_  (.A1(\u_cpu.ALU.u_wallace._0139_ ),
    .A2(\u_cpu.ALU.u_wallace._0143_ ),
    .B1(\u_cpu.ALU.u_wallace._0149_ ),
    .Y(\u_cpu.ALU.u_wallace._0150_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5978_  (.A1(\u_cpu.ALU.u_wallace._0134_ ),
    .A2(\u_cpu.ALU.u_wallace._0135_ ),
    .B1(\u_cpu.ALU.u_wallace._0136_ ),
    .C1(\u_cpu.ALU.u_wallace._0138_ ),
    .Y(\u_cpu.ALU.u_wallace._0152_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._5979_  (.A1(\u_cpu.ALU.u_wallace._0138_ ),
    .A2(\u_cpu.ALU.u_wallace._0142_ ),
    .B1(\u_cpu.ALU.u_wallace._0136_ ),
    .X(\u_cpu.ALU.u_wallace._0153_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._5980_  (.A1(\u_cpu.ALU.u_wallace._0147_ ),
    .A2(\u_cpu.ALU.u_wallace._0148_ ),
    .B1(\u_cpu.ALU.u_wallace._0152_ ),
    .C1(\u_cpu.ALU.u_wallace._0153_ ),
    .Y(\u_cpu.ALU.u_wallace._0154_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5981_  (.A(\u_cpu.ALU.u_wallace._0132_ ),
    .B(\u_cpu.ALU.u_wallace._0150_ ),
    .C(\u_cpu.ALU.u_wallace._0154_ ),
    .Y(\u_cpu.ALU.u_wallace._0155_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5982_  (.A1(\u_cpu.ALU.u_wallace._4933_ ),
    .A2(\u_cpu.ALU.u_wallace._0011_ ),
    .B1(\u_cpu.ALU.u_wallace._0013_ ),
    .Y(\u_cpu.ALU.u_wallace._0156_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5983_  (.A(\u_cpu.ALU.u_wallace._0153_ ),
    .B(\u_cpu.ALU.u_wallace._0149_ ),
    .C(\u_cpu.ALU.u_wallace._0152_ ),
    .Y(\u_cpu.ALU.u_wallace._0157_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5984_  (.A1(\u_cpu.ALU.u_wallace._0147_ ),
    .A2(\u_cpu.ALU.u_wallace._0148_ ),
    .B1(\u_cpu.ALU.u_wallace._0139_ ),
    .B2(\u_cpu.ALU.u_wallace._0143_ ),
    .Y(\u_cpu.ALU.u_wallace._0158_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5985_  (.A(\u_cpu.ALU.u_wallace._0156_ ),
    .B(\u_cpu.ALU.u_wallace._0157_ ),
    .C(\u_cpu.ALU.u_wallace._0158_ ),
    .Y(\u_cpu.ALU.u_wallace._0159_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.ALU.u_wallace._5986_  (.A1(\u_cpu.ALU.u_wallace._0056_ ),
    .A2(\u_cpu.ALU.u_wallace._0058_ ),
    .A3(\u_cpu.ALU.u_wallace._0054_ ),
    .B1(\u_cpu.ALU.u_wallace._0059_ ),
    .Y(\u_cpu.ALU.u_wallace._0160_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._5987_  (.A1(\u_cpu.ALU.u_wallace._0155_ ),
    .A2(\u_cpu.ALU.u_wallace._0159_ ),
    .B1(\u_cpu.ALU.u_wallace._0160_ ),
    .Y(\u_cpu.ALU.u_wallace._0161_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._5988_  (.A(\u_cpu.ALU.u_wallace._0160_ ),
    .B(\u_cpu.ALU.u_wallace._0155_ ),
    .C(\u_cpu.ALU.u_wallace._0159_ ),
    .X(\u_cpu.ALU.u_wallace._0163_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._5989_  (.A(\u_cpu.ALU.u_wallace._4916_ ),
    .B(\u_cpu.ALU.u_wallace._4927_ ),
    .Y(\u_cpu.ALU.u_wallace._0164_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._5990_  (.A1(\u_cpu.ALU.u_wallace._0008_ ),
    .A2(\u_cpu.ALU.u_wallace._0011_ ),
    .B1(\u_cpu.ALU.u_wallace._0016_ ),
    .Y(\u_cpu.ALU.u_wallace._0165_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._5991_  (.A(\u_cpu.ALU.u_wallace._0014_ ),
    .B(\u_cpu.ALU.u_wallace._4933_ ),
    .C(\u_cpu.ALU.u_wallace._0013_ ),
    .Y(\u_cpu.ALU.u_wallace._0166_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5992_  (.A1(\u_cpu.ALU.u_wallace._4931_ ),
    .A2(\u_cpu.ALU.u_wallace._0164_ ),
    .B1(\u_cpu.ALU.u_wallace._0165_ ),
    .B2(\u_cpu.ALU.u_wallace._0166_ ),
    .Y(\u_cpu.ALU.u_wallace._0167_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._5993_  (.A1(\u_cpu.ALU.u_wallace._4903_ ),
    .A2(\u_cpu.ALU.u_wallace._4906_ ),
    .A3(\u_cpu.ALU.u_wallace._4926_ ),
    .B1(\u_cpu.ALU.u_wallace._4911_ ),
    .X(\u_cpu.ALU.u_wallace._0168_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._5994_  (.A(\u_cpu.ALU.u_wallace._4797_ ),
    .Y(\u_cpu.ALU.u_wallace._0169_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._5995_  (.A1(\u_cpu.ALU.u_wallace._0282_ ),
    .A2(\u_cpu.ALU.SrcA[12] ),
    .B1(\u_cpu.ALU.SrcA[13] ),
    .B2(\u_cpu.ALU.u_wallace._0195_ ),
    .Y(\u_cpu.ALU.u_wallace._0170_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._5996_  (.A(\u_cpu.ALU.u_wallace._1903_ ),
    .B(\u_cpu.ALU.u_wallace._0807_ ),
    .C(\u_cpu.ALU.u_wallace._4790_ ),
    .D(\u_cpu.ALU.u_wallace._4920_ ),
    .X(\u_cpu.ALU.u_wallace._0171_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._5997_  (.A1(\u_cpu.ALU.u_wallace._1224_ ),
    .A2(\u_cpu.ALU.u_wallace._0169_ ),
    .B1(\u_cpu.ALU.u_wallace._0170_ ),
    .B2(\u_cpu.ALU.u_wallace._0171_ ),
    .Y(\u_cpu.ALU.u_wallace._0172_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._5998_  (.A1(\u_cpu.ALU.u_wallace._1968_ ),
    .A2(\u_cpu.ALU.u_wallace._4785_ ),
    .B1(\u_cpu.ALU.u_wallace._4907_ ),
    .B2(\u_cpu.ALU.u_wallace._4657_ ),
    .X(\u_cpu.ALU.u_wallace._0174_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._5999_  (.A(\u_cpu.ALU.u_wallace._0775_ ),
    .B(\u_cpu.ALU.u_wallace._0534_ ),
    .C(\u_cpu.ALU.SrcA[12] ),
    .D(\u_cpu.ALU.u_wallace._4920_ ),
    .Y(\u_cpu.ALU.u_wallace._0175_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6000_  (.A(\u_cpu.ALU.u_wallace._0174_ ),
    .B(\u_cpu.ALU.u_wallace._0175_ ),
    .C(\u_cpu.ALU.u_wallace._4662_ ),
    .D(\u_cpu.ALU.u_wallace._4798_ ),
    .Y(\u_cpu.ALU.u_wallace._0176_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6001_  (.A(\u_cpu.ALU.SrcA[14] ),
    .X(\u_cpu.ALU.u_wallace._0177_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6002_  (.A1(\u_cpu.ALU.u_wallace._2856_ ),
    .A2(\u_cpu.ALU.u_wallace._3689_ ),
    .B1(\u_cpu.ALU.u_wallace._0177_ ),
    .B2(\u_cpu.ALU.u_wallace._2747_ ),
    .Y(\u_cpu.ALU.u_wallace._0178_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6003_  (.A(\u_cpu.ALU.SrcA[14] ),
    .X(\u_cpu.ALU.u_wallace._0179_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6004_  (.A(\u_cpu.ALU.u_wallace._1859_ ),
    .B(\u_cpu.ALU.u_wallace._1826_ ),
    .C(\u_cpu.ALU.u_wallace._4449_ ),
    .D(\u_cpu.ALU.u_wallace._0179_ ),
    .Y(\u_cpu.ALU.u_wallace._0180_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._6005_  (.A_N(\u_cpu.ALU.u_wallace._0178_ ),
    .B(\u_cpu.ALU.u_wallace._0180_ ),
    .C(\u_cpu.ALU.u_wallace._4910_ ),
    .Y(\u_cpu.ALU.u_wallace._0181_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6006_  (.A(\u_cpu.ALU.SrcA[14] ),
    .X(\u_cpu.ALU.u_wallace._0182_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6007_  (.A(\u_cpu.ALU.u_wallace._0862_ ),
    .B(\u_cpu.ALU.u_wallace._2768_ ),
    .C(\u_cpu.ALU.u_wallace._3645_ ),
    .D(\u_cpu.ALU.u_wallace._0182_ ),
    .X(\u_cpu.ALU.u_wallace._0183_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6008_  (.A1(\u_cpu.ALU.u_wallace._0178_ ),
    .A2(\u_cpu.ALU.u_wallace._0183_ ),
    .B1(\u_cpu.ALU.u_wallace._4922_ ),
    .Y(\u_cpu.ALU.u_wallace._0185_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6009_  (.A1(\u_cpu.ALU.u_wallace._0172_ ),
    .A2(\u_cpu.ALU.u_wallace._0176_ ),
    .B1(\u_cpu.ALU.u_wallace._0181_ ),
    .B2(\u_cpu.ALU.u_wallace._0185_ ),
    .X(\u_cpu.ALU.u_wallace._0186_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6010_  (.A(\u_cpu.ALU.u_wallace._1903_ ),
    .X(\u_cpu.ALU.u_wallace._0187_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6011_  (.A(\u_cpu.ALU.u_wallace._4920_ ),
    .X(\u_cpu.ALU.u_wallace._0188_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6012_  (.A(\u_cpu.ALU.u_wallace._0742_ ),
    .B(\u_cpu.ALU.u_wallace._4650_ ),
    .Y(\u_cpu.ALU.u_wallace._0189_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._6013_  (.A1(\u_cpu.ALU.u_wallace._0187_ ),
    .A2(\u_cpu.ALU.u_wallace._0304_ ),
    .A3(\u_cpu.ALU.u_wallace._4917_ ),
    .A4(\u_cpu.ALU.u_wallace._0188_ ),
    .B1(\u_cpu.ALU.u_wallace._0189_ ),
    .X(\u_cpu.ALU.u_wallace._0190_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._6014_  (.A1(\u_cpu.ALU.u_wallace._0190_ ),
    .A2(\u_cpu.ALU.u_wallace._0170_ ),
    .B1(\u_cpu.ALU.u_wallace._0172_ ),
    .C1(\u_cpu.ALU.u_wallace._0181_ ),
    .D1(\u_cpu.ALU.u_wallace._0185_ ),
    .Y(\u_cpu.ALU.u_wallace._0191_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6015_  (.A(\u_cpu.ALU.u_wallace._0168_ ),
    .B(\u_cpu.ALU.u_wallace._0186_ ),
    .C(\u_cpu.ALU.u_wallace._0191_ ),
    .Y(\u_cpu.ALU.u_wallace._0192_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6016_  (.A1(\u_cpu.ALU.u_wallace._0172_ ),
    .A2(\u_cpu.ALU.u_wallace._0176_ ),
    .B1(\u_cpu.ALU.u_wallace._0181_ ),
    .B2(\u_cpu.ALU.u_wallace._0185_ ),
    .Y(\u_cpu.ALU.u_wallace._0193_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._6017_  (.A1(\u_cpu.ALU.u_wallace._0190_ ),
    .A2(\u_cpu.ALU.u_wallace._0170_ ),
    .B1(\u_cpu.ALU.u_wallace._0172_ ),
    .C1(\u_cpu.ALU.u_wallace._0181_ ),
    .D1(\u_cpu.ALU.u_wallace._0185_ ),
    .X(\u_cpu.ALU.u_wallace._0194_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._6018_  (.A1(\u_cpu.ALU.u_wallace._4903_ ),
    .A2(\u_cpu.ALU.u_wallace._4906_ ),
    .A3(\u_cpu.ALU.u_wallace._4926_ ),
    .B1(\u_cpu.ALU.u_wallace._4911_ ),
    .Y(\u_cpu.ALU.u_wallace._0196_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6019_  (.A1(\u_cpu.ALU.u_wallace._0193_ ),
    .A2(\u_cpu.ALU.u_wallace._0194_ ),
    .B1(\u_cpu.ALU.u_wallace._0196_ ),
    .Y(\u_cpu.ALU.u_wallace._0197_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6020_  (.A(\u_cpu.ALU.u_wallace._1848_ ),
    .X(\u_cpu.ALU.u_wallace._0198_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6021_  (.A(\u_cpu.ALU.u_wallace._0002_ ),
    .B(\u_cpu.ALU.u_wallace._0015_ ),
    .C(\u_cpu.ALU.u_wallace._0198_ ),
    .Y(\u_cpu.ALU.u_wallace._0199_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6022_  (.A1(\u_cpu.ALU.u_wallace._2538_ ),
    .A2(\u_cpu.ALU.u_wallace._4444_ ),
    .B1(\u_cpu.ALU.u_wallace._4557_ ),
    .B2(\u_cpu.ALU.u_wallace._1465_ ),
    .X(\u_cpu.ALU.u_wallace._0200_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6023_  (.A(\u_cpu.ALU.u_wallace._2045_ ),
    .B(\u_cpu.ALU.u_wallace._2582_ ),
    .C(\u_cpu.ALU.u_wallace._4439_ ),
    .D(\u_cpu.ALU.u_wallace._4642_ ),
    .Y(\u_cpu.ALU.u_wallace._0201_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6024_  (.A(\u_cpu.ALU.u_wallace._0200_ ),
    .B(\u_cpu.ALU.u_wallace._0201_ ),
    .C(\u_cpu.ALU.u_wallace._2801_ ),
    .D(\u_cpu.ALU.u_wallace._2626_ ),
    .Y(\u_cpu.ALU.u_wallace._0202_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._6025_  (.A(\u_cpu.ALU.u_wallace._4447_ ),
    .Y(\u_cpu.ALU.u_wallace._0203_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6026_  (.A1(\u_cpu.ALU.u_wallace._2582_ ),
    .A2(\u_cpu.ALU.u_wallace._4439_ ),
    .B1(\u_cpu.ALU.u_wallace._4551_ ),
    .B2(\u_cpu.ALU.u_wallace._2571_ ),
    .Y(\u_cpu.ALU.u_wallace._0204_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6027_  (.A(\u_cpu.ALU.u_wallace._2144_ ),
    .B(\u_cpu.ALU.u_wallace._2538_ ),
    .C(\u_cpu.ALU.u_wallace._4444_ ),
    .D(\u_cpu.ALU.u_wallace._4553_ ),
    .X(\u_cpu.ALU.u_wallace._0205_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6028_  (.A1(\u_cpu.ALU.u_wallace._0203_ ),
    .A2(\u_cpu.ALU.u_wallace._4471_ ),
    .B1(\u_cpu.ALU.u_wallace._0204_ ),
    .B2(\u_cpu.ALU.u_wallace._0205_ ),
    .Y(\u_cpu.ALU.u_wallace._0207_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6029_  (.A(\u_cpu.ALU.u_wallace._0202_ ),
    .B(\u_cpu.ALU.u_wallace._0207_ ),
    .Y(\u_cpu.ALU.u_wallace._0208_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._6030_  (.A1(\u_cpu.ALU.u_wallace._4678_ ),
    .A2(\u_cpu.ALU.u_wallace._4904_ ),
    .A3(\u_cpu.ALU.u_wallace._4901_ ),
    .B1(\u_cpu.ALU.u_wallace._4902_ ),
    .X(\u_cpu.ALU.u_wallace._0209_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6031_  (.A(\u_cpu.ALU.u_wallace._4796_ ),
    .B(\u_cpu.ALU.u_wallace._4794_ ),
    .Y(\u_cpu.ALU.u_wallace._0210_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6032_  (.A(\u_cpu.ALU.u_wallace._0187_ ),
    .B(\u_cpu.ALU.u_wallace._4917_ ),
    .Y(\u_cpu.ALU.u_wallace._0211_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6033_  (.A1(\u_cpu.ALU.u_wallace._0210_ ),
    .A2(\u_cpu.ALU.u_wallace._0211_ ),
    .B1(\u_cpu.ALU.u_wallace._4918_ ),
    .Y(\u_cpu.ALU.u_wallace._0212_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6034_  (.A1(\u_cpu.ALU.u_wallace._4905_ ),
    .A2(\u_cpu.ALU.u_wallace._0212_ ),
    .B1(\u_cpu.ALU.u_wallace._0202_ ),
    .C1(\u_cpu.ALU.u_wallace._0207_ ),
    .X(\u_cpu.ALU.u_wallace._0213_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.ALU.u_wallace._6035_  (.A1(\u_cpu.ALU.u_wallace._0003_ ),
    .A2(\u_cpu.ALU.u_wallace._0199_ ),
    .B1(\u_cpu.ALU.u_wallace._0208_ ),
    .B2(\u_cpu.ALU.u_wallace._0209_ ),
    .C1(\u_cpu.ALU.u_wallace._0213_ ),
    .Y(\u_cpu.ALU.u_wallace._0214_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6036_  (.A1(\u_cpu.ALU.u_wallace._4918_ ),
    .A2(\u_cpu.ALU.u_wallace._4901_ ),
    .B1(\u_cpu.ALU.u_wallace._4902_ ),
    .Y(\u_cpu.ALU.u_wallace._0215_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6037_  (.A1(\u_cpu.ALU.u_wallace._0202_ ),
    .A2(\u_cpu.ALU.u_wallace._0207_ ),
    .B1(\u_cpu.ALU.u_wallace._0215_ ),
    .Y(\u_cpu.ALU.u_wallace._0216_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._6038_  (.A1(\u_cpu.ALU.u_wallace._4454_ ),
    .A2(\u_cpu.ALU.u_wallace._4539_ ),
    .A3(\u_cpu.ALU.u_wallace._0005_ ),
    .B1(\u_cpu.ALU.u_wallace._0003_ ),
    .X(\u_cpu.ALU.u_wallace._0218_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._6039_  (.A1(\u_cpu.ALU.u_wallace._0213_ ),
    .A2(\u_cpu.ALU.u_wallace._0216_ ),
    .B1(\u_cpu.ALU.u_wallace._0218_ ),
    .X(\u_cpu.ALU.u_wallace._0219_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6040_  (.A1_N(\u_cpu.ALU.u_wallace._0192_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0197_ ),
    .B1(\u_cpu.ALU.u_wallace._0214_ ),
    .B2(\u_cpu.ALU.u_wallace._0219_ ),
    .Y(\u_cpu.ALU.u_wallace._0220_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6041_  (.A1(\u_cpu.ALU.u_wallace._4905_ ),
    .A2(\u_cpu.ALU.u_wallace._0212_ ),
    .B1(\u_cpu.ALU.u_wallace._0202_ ),
    .C1(\u_cpu.ALU.u_wallace._0207_ ),
    .Y(\u_cpu.ALU.u_wallace._0221_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6042_  (.A1(\u_cpu.ALU.u_wallace._0202_ ),
    .A2(\u_cpu.ALU.u_wallace._0207_ ),
    .B1(\u_cpu.ALU.u_wallace._0215_ ),
    .X(\u_cpu.ALU.u_wallace._0222_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._6043_  (.A_N(\u_cpu.ALU.u_wallace._0218_ ),
    .B(\u_cpu.ALU.u_wallace._0221_ ),
    .C(\u_cpu.ALU.u_wallace._0222_ ),
    .Y(\u_cpu.ALU.u_wallace._0223_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6044_  (.A1(\u_cpu.ALU.u_wallace._0213_ ),
    .A2(\u_cpu.ALU.u_wallace._0216_ ),
    .B1(\u_cpu.ALU.u_wallace._0218_ ),
    .Y(\u_cpu.ALU.u_wallace._0224_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6045_  (.A(\u_cpu.ALU.u_wallace._0192_ ),
    .B(\u_cpu.ALU.u_wallace._0197_ ),
    .C(\u_cpu.ALU.u_wallace._0223_ ),
    .D(\u_cpu.ALU.u_wallace._0224_ ),
    .Y(\u_cpu.ALU.u_wallace._0225_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6046_  (.A1(\u_cpu.ALU.u_wallace._0072_ ),
    .A2(\u_cpu.ALU.u_wallace._0167_ ),
    .B1(\u_cpu.ALU.u_wallace._0220_ ),
    .C1(\u_cpu.ALU.u_wallace._0225_ ),
    .X(\u_cpu.ALU.u_wallace._0226_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU.u_wallace._6047_  (.A1(\u_cpu.ALU.u_wallace._0220_ ),
    .A2(\u_cpu.ALU.u_wallace._0225_ ),
    .B1(\u_cpu.ALU.u_wallace._0072_ ),
    .C1(\u_cpu.ALU.u_wallace._0167_ ),
    .Y(\u_cpu.ALU.u_wallace._0227_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6048_  (.A1(\u_cpu.ALU.u_wallace._0161_ ),
    .A2(\u_cpu.ALU.u_wallace._0163_ ),
    .B1(\u_cpu.ALU.u_wallace._0226_ ),
    .B2(\u_cpu.ALU.u_wallace._0227_ ),
    .Y(\u_cpu.ALU.u_wallace._0229_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6049_  (.A1(\u_cpu.ALU.u_wallace._0155_ ),
    .A2(\u_cpu.ALU.u_wallace._0159_ ),
    .B1(\u_cpu.ALU.u_wallace._0160_ ),
    .X(\u_cpu.ALU.u_wallace._0230_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6050_  (.A(\u_cpu.ALU.u_wallace._0160_ ),
    .B(\u_cpu.ALU.u_wallace._0155_ ),
    .C(\u_cpu.ALU.u_wallace._0159_ ),
    .Y(\u_cpu.ALU.u_wallace._0231_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6051_  (.A1(\u_cpu.ALU.u_wallace._0072_ ),
    .A2(\u_cpu.ALU.u_wallace._0167_ ),
    .B1(\u_cpu.ALU.u_wallace._0220_ ),
    .C1(\u_cpu.ALU.u_wallace._0225_ ),
    .Y(\u_cpu.ALU.u_wallace._0232_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6052_  (.A(\u_cpu.ALU.u_wallace._0220_ ),
    .B(\u_cpu.ALU.u_wallace._0225_ ),
    .Y(\u_cpu.ALU.u_wallace._0233_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._6053_  (.A1(\u_cpu.ALU.u_wallace._4932_ ),
    .A2(\u_cpu.ALU.u_wallace._0019_ ),
    .A3(\u_cpu.ALU.u_wallace._0020_ ),
    .B1(\u_cpu.ALU.u_wallace._0072_ ),
    .Y(\u_cpu.ALU.u_wallace._0234_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6054_  (.A(\u_cpu.ALU.u_wallace._0233_ ),
    .B(\u_cpu.ALU.u_wallace._0234_ ),
    .Y(\u_cpu.ALU.u_wallace._0235_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6055_  (.A(\u_cpu.ALU.u_wallace._0230_ ),
    .B(\u_cpu.ALU.u_wallace._0231_ ),
    .C(\u_cpu.ALU.u_wallace._0232_ ),
    .D(\u_cpu.ALU.u_wallace._0235_ ),
    .Y(\u_cpu.ALU.u_wallace._0236_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6056_  (.A(\u_cpu.ALU.u_wallace._0069_ ),
    .B(\u_cpu.ALU.u_wallace._0070_ ),
    .Y(\u_cpu.ALU.u_wallace._0237_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6057_  (.A1(\u_cpu.ALU.u_wallace._0025_ ),
    .A2(\u_cpu.ALU.u_wallace._0237_ ),
    .B1(\u_cpu.ALU.u_wallace._0079_ ),
    .Y(\u_cpu.ALU.u_wallace._0238_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6058_  (.A1(\u_cpu.ALU.u_wallace._0229_ ),
    .A2(\u_cpu.ALU.u_wallace._0236_ ),
    .B1(\u_cpu.ALU.u_wallace._0238_ ),
    .X(\u_cpu.ALU.u_wallace._0240_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6059_  (.A1(\u_cpu.ALU.u_wallace._0234_ ),
    .A2(\u_cpu.ALU.u_wallace._0233_ ),
    .B1(\u_cpu.ALU.u_wallace._0230_ ),
    .C1(\u_cpu.ALU.u_wallace._0231_ ),
    .Y(\u_cpu.ALU.u_wallace._0241_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6060_  (.A1(\u_cpu.ALU.u_wallace._0227_ ),
    .A2(\u_cpu.ALU.u_wallace._0241_ ),
    .B1(\u_cpu.ALU.u_wallace._0229_ ),
    .C1(\u_cpu.ALU.u_wallace._0238_ ),
    .Y(\u_cpu.ALU.u_wallace._0242_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._6061_  (.A_N(\u_cpu.ALU.u_wallace._0131_ ),
    .B(\u_cpu.ALU.u_wallace._0240_ ),
    .C(\u_cpu.ALU.u_wallace._0242_ ),
    .Y(\u_cpu.ALU.u_wallace._0243_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._6062_  (.A(\u_cpu.ALU.u_wallace._0130_ ),
    .Y(\u_cpu.ALU.u_wallace._0244_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6063_  (.A1(\u_cpu.ALU.u_wallace._0229_ ),
    .A2(\u_cpu.ALU.u_wallace._0236_ ),
    .B1(\u_cpu.ALU.u_wallace._0238_ ),
    .Y(\u_cpu.ALU.u_wallace._0245_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6064_  (.A1(\u_cpu.ALU.u_wallace._0227_ ),
    .A2(\u_cpu.ALU.u_wallace._0241_ ),
    .B1(\u_cpu.ALU.u_wallace._0229_ ),
    .C1(\u_cpu.ALU.u_wallace._0238_ ),
    .X(\u_cpu.ALU.u_wallace._0246_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6065_  (.A1(\u_cpu.ALU.u_wallace._0128_ ),
    .A2(\u_cpu.ALU.u_wallace._0244_ ),
    .B1(\u_cpu.ALU.u_wallace._0245_ ),
    .B2(\u_cpu.ALU.u_wallace._0246_ ),
    .Y(\u_cpu.ALU.u_wallace._0247_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6066_  (.A(\u_cpu.ALU.u_wallace._0116_ ),
    .B(\u_cpu.ALU.u_wallace._0243_ ),
    .C(\u_cpu.ALU.u_wallace._0247_ ),
    .Y(\u_cpu.ALU.u_wallace._0248_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6067_  (.A(\u_cpu.ALU.u_wallace._0243_ ),
    .B(\u_cpu.ALU.u_wallace._0247_ ),
    .Y(\u_cpu.ALU.u_wallace._0249_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._6068_  (.A1(\u_cpu.ALU.u_wallace._4896_ ),
    .A2(\u_cpu.ALU.u_wallace._4897_ ),
    .A3(\u_cpu.ALU.u_wallace._0091_ ),
    .B1(\u_cpu.ALU.u_wallace._0094_ ),
    .X(\u_cpu.ALU.u_wallace._0251_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6069_  (.A1(\u_cpu.ALU.u_wallace._4868_ ),
    .A2(\u_cpu.ALU.u_wallace._4867_ ),
    .B1(\u_cpu.ALU.u_wallace._4895_ ),
    .X(\u_cpu.ALU.u_wallace._0252_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6070_  (.A1(\u_cpu.ALU.u_wallace._0249_ ),
    .A2(\u_cpu.ALU.u_wallace._0251_ ),
    .B1(\u_cpu.ALU.u_wallace._0252_ ),
    .Y(\u_cpu.ALU.u_wallace._0253_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6071_  (.A1(\u_cpu.ALU.u_wallace._0243_ ),
    .A2(\u_cpu.ALU.u_wallace._0247_ ),
    .B1(\u_cpu.ALU.u_wallace._0116_ ),
    .X(\u_cpu.ALU.u_wallace._0254_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6072_  (.A(\u_cpu.ALU.u_wallace._0248_ ),
    .B(\u_cpu.ALU.u_wallace._0254_ ),
    .Y(\u_cpu.ALU.u_wallace._0255_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6073_  (.A1(\u_cpu.ALU.u_wallace._0248_ ),
    .A2(\u_cpu.ALU.u_wallace._0253_ ),
    .B1(\u_cpu.ALU.u_wallace._0255_ ),
    .B2(\u_cpu.ALU.u_wallace._0252_ ),
    .Y(\u_cpu.ALU.u_wallace._0256_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6074_  (.A1(\u_cpu.ALU.u_wallace._4882_ ),
    .A2(\u_cpu.ALU.u_wallace._0115_ ),
    .B1(\u_cpu.ALU.u_wallace._0100_ ),
    .C1(\u_cpu.ALU.u_wallace._0256_ ),
    .X(\u_cpu.ALU.u_wallace._0257_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6075_  (.A(\u_cpu.ALU.u_wallace._0116_ ),
    .B(\u_cpu.ALU.u_wallace._0243_ ),
    .C(\u_cpu.ALU.u_wallace._0247_ ),
    .X(\u_cpu.ALU.u_wallace._0258_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._6076_  (.A1(\u_cpu.ALU.u_wallace._0094_ ),
    .A2(\u_cpu.ALU.u_wallace._0249_ ),
    .B1(\u_cpu.ALU.u_wallace._0252_ ),
    .C1(\u_cpu.ALU.u_wallace._0258_ ),
    .X(\u_cpu.ALU.u_wallace._0259_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6077_  (.A1(\u_cpu.ALU.u_wallace._0243_ ),
    .A2(\u_cpu.ALU.u_wallace._0247_ ),
    .B1(\u_cpu.ALU.u_wallace._0116_ ),
    .Y(\u_cpu.ALU.u_wallace._0260_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6078_  (.A1(\u_cpu.ALU.u_wallace._0258_ ),
    .A2(\u_cpu.ALU.u_wallace._0260_ ),
    .B1(\u_cpu.ALU.u_wallace._0252_ ),
    .Y(\u_cpu.ALU.u_wallace._0262_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6079_  (.A(\u_cpu.ALU.u_wallace._4769_ ),
    .B(\u_cpu.ALU.u_wallace._4878_ ),
    .C(\u_cpu.ALU.u_wallace._4881_ ),
    .D(\u_cpu.ALU.u_wallace._0099_ ),
    .X(\u_cpu.ALU.u_wallace._0263_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._6080_  (.A(\u_cpu.ALU.u_wallace._0100_ ),
    .Y(\u_cpu.ALU.u_wallace._0264_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU.u_wallace._6081_  (.A1_N(\u_cpu.ALU.u_wallace._0259_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0262_ ),
    .B1(\u_cpu.ALU.u_wallace._0263_ ),
    .B2(\u_cpu.ALU.u_wallace._0264_ ),
    .X(\u_cpu.ALU.u_wallace._0265_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._6082_  (.A(\u_cpu.ALU.u_wallace._0257_ ),
    .B(\u_cpu.ALU.u_wallace._0265_ ),
    .Y(\u_cpu.ALU.u_wallace._0266_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6083_  (.A1(\u_cpu.ALU.u_wallace._0107_ ),
    .A2(\u_cpu.ALU.u_wallace._0114_ ),
    .B1(\u_cpu.ALU.u_wallace._0266_ ),
    .Y(\u_cpu.ALU.u_wallace._0267_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.ALU.u_wallace._6084_  (.A_N(\u_cpu.ALU.u_wallace._0102_ ),
    .B(\u_cpu.ALU.u_wallace._0100_ ),
    .C(\u_cpu.ALU.u_wallace._0099_ ),
    .D(\u_cpu.ALU.u_wallace._4882_ ),
    .X(\u_cpu.ALU.u_wallace._0268_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6085_  (.A1(\u_cpu.ALU.u_wallace._0257_ ),
    .A2(\u_cpu.ALU.u_wallace._0265_ ),
    .B1(\u_cpu.ALU.u_wallace._0268_ ),
    .Y(\u_cpu.ALU.u_wallace._0269_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6086_  (.A(\u_cpu.ALU.u_wallace._0267_ ),
    .B(\u_cpu.ALU.u_wallace._0269_ ),
    .Y(\u_cpu.ALU.u_wallace._0270_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6087_  (.A1(\u_cpu.ALU.u_wallace._4884_ ),
    .A2(\u_cpu.ALU.u_wallace._4888_ ),
    .B1(\u_cpu.ALU.u_wallace._4889_ ),
    .X(\u_cpu.ALU.u_wallace._0271_ ));
 sky130_fd_sc_hd__a32oi_2 \u_cpu.ALU.u_wallace._6088_  (.A1(\u_cpu.ALU.u_wallace._0109_ ),
    .A2(\u_cpu.ALU.u_wallace._0110_ ),
    .A3(\u_cpu.ALU.u_wallace._0105_ ),
    .B1(\u_cpu.ALU.u_wallace._0106_ ),
    .B2(\u_cpu.ALU.u_wallace._0271_ ),
    .Y(\u_cpu.ALU.u_wallace._0273_ ));
 sky130_fd_sc_hd__a41oi_2 \u_cpu.ALU.u_wallace._6089_  (.A1(\u_cpu.ALU.u_wallace._4766_ ),
    .A2(\u_cpu.ALU.u_wallace._4893_ ),
    .A3(\u_cpu.ALU.u_wallace._0106_ ),
    .A4(\u_cpu.ALU.u_wallace._0111_ ),
    .B1(\u_cpu.ALU.u_wallace._0273_ ),
    .Y(\u_cpu.ALU.u_wallace._0274_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._6090_  (.A(\u_cpu.ALU.u_wallace._0270_ ),
    .B(\u_cpu.ALU.u_wallace._0274_ ),
    .X(\u_cpu.ALU.Product_Wallace[14] ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6091_  (.A(\u_cpu.ALU.u_wallace._0256_ ),
    .B(\u_cpu.ALU.u_wallace._0263_ ),
    .C(\u_cpu.ALU.u_wallace._0100_ ),
    .X(\u_cpu.ALU.u_wallace._0275_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._6092_  (.A1(\u_cpu.ALU.u_wallace._0131_ ),
    .A2(\u_cpu.ALU.u_wallace._0245_ ),
    .B1(\u_cpu.ALU.u_wallace._0242_ ),
    .X(\u_cpu.ALU.u_wallace._0276_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6093_  (.A(\u_cpu.ALU.u_wallace._0159_ ),
    .B(\u_cpu.ALU.u_wallace._0231_ ),
    .Y(\u_cpu.ALU.u_wallace._0277_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6094_  (.A(\u_cpu.ALU.SrcB[15] ),
    .X(\u_cpu.ALU.u_wallace._0278_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6095_  (.A(\u_cpu.ALU.u_wallace._0278_ ),
    .X(\u_cpu.ALU.u_wallace._0279_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6096_  (.A(\u_cpu.ALU.u_wallace._0279_ ),
    .X(\u_cpu.ALU.u_wallace._0280_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6097_  (.A1(\u_cpu.ALU.u_wallace._4463_ ),
    .A2(\u_cpu.ALU.u_wallace._0121_ ),
    .B1(\u_cpu.ALU.u_wallace._0280_ ),
    .B2(\u_cpu.ALU.u_wallace._0108_ ),
    .X(\u_cpu.ALU.u_wallace._0281_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6098_  (.A(\u_cpu.ALU.u_wallace._0108_ ),
    .B(\u_cpu.ALU.u_wallace._0162_ ),
    .C(\u_cpu.ALU.u_wallace._0122_ ),
    .D(\u_cpu.ALU.u_wallace._0280_ ),
    .Y(\u_cpu.ALU.u_wallace._0283_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6099_  (.A(\u_cpu.ALU.u_wallace._1410_ ),
    .B(\u_cpu.ALU.u_wallace._1191_ ),
    .C(\u_cpu.ALU.u_wallace._4837_ ),
    .D(\u_cpu.ALU.u_wallace._0029_ ),
    .X(\u_cpu.ALU.u_wallace._0284_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._6100_  (.A1(\u_cpu.ALU.u_wallace._0145_ ),
    .A2(\u_cpu.ALU.u_wallace._0057_ ),
    .A3(\u_cpu.ALU.u_wallace._4463_ ),
    .B1(\u_cpu.ALU.u_wallace._0284_ ),
    .X(\u_cpu.ALU.u_wallace._0285_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6101_  (.A1(\u_cpu.ALU.u_wallace._0281_ ),
    .A2(\u_cpu.ALU.u_wallace._0283_ ),
    .B1(\u_cpu.ALU.u_wallace._0285_ ),
    .X(\u_cpu.ALU.u_wallace._0286_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6102_  (.A(\u_cpu.ALU.u_wallace._0285_ ),
    .B(\u_cpu.ALU.u_wallace._0281_ ),
    .C(\u_cpu.ALU.u_wallace._0283_ ),
    .Y(\u_cpu.ALU.u_wallace._0287_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6103_  (.A(\u_cpu.ALU.u_wallace._0286_ ),
    .B(\u_cpu.ALU.u_wallace._0287_ ),
    .Y(\u_cpu.ALU.u_wallace._0288_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._6104_  (.A(\u_cpu.ALU.u_wallace._0123_ ),
    .B(\u_cpu.ALU.u_wallace._0288_ ),
    .X(\u_cpu.ALU.u_wallace._0289_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._6105_  (.A(\u_cpu.ALU.u_wallace._0277_ ),
    .B(\u_cpu.ALU.u_wallace._0289_ ),
    .X(\u_cpu.ALU.u_wallace._0290_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._6106_  (.A(\u_cpu.ALU.u_wallace._0277_ ),
    .B(\u_cpu.ALU.u_wallace._0289_ ),
    .Y(\u_cpu.ALU.u_wallace._0291_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6107_  (.A1(\u_cpu.ALU.u_wallace._1486_ ),
    .A2(\u_cpu.ALU.SrcA[10] ),
    .B1(\u_cpu.ALU.u_wallace._4646_ ),
    .B2(\u_cpu.ALU.SrcB[4] ),
    .Y(\u_cpu.ALU.u_wallace._0292_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6108_  (.A(\u_cpu.ALU.u_wallace._1026_ ),
    .B(\u_cpu.ALU.u_wallace._1486_ ),
    .C(\u_cpu.ALU.u_wallace._4550_ ),
    .D(\u_cpu.ALU.u_wallace._4646_ ),
    .Y(\u_cpu.ALU.u_wallace._0294_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._6109_  (.A_N(\u_cpu.ALU.u_wallace._0292_ ),
    .B(\u_cpu.ALU.u_wallace._0294_ ),
    .C(\u_cpu.ALU.u_wallace._4449_ ),
    .D(\u_cpu.ALU.SrcB[7] ),
    .Y(\u_cpu.ALU.u_wallace._0295_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6110_  (.A(\u_cpu.ALU.SrcB[4] ),
    .B(\u_cpu.ALU.SrcB[5] ),
    .C(\u_cpu.ALU.SrcA[10] ),
    .D(\u_cpu.ALU.SrcA[11] ),
    .X(\u_cpu.ALU.u_wallace._0296_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6111_  (.A1(\u_cpu.ALU.u_wallace._4676_ ),
    .A2(\u_cpu.ALU.u_wallace._4470_ ),
    .B1(\u_cpu.ALU.u_wallace._0292_ ),
    .B2(\u_cpu.ALU.u_wallace._0296_ ),
    .Y(\u_cpu.ALU.u_wallace._0297_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6112_  (.A1(\u_cpu.ALU.u_wallace._0189_ ),
    .A2(\u_cpu.ALU.u_wallace._0170_ ),
    .B1(\u_cpu.ALU.u_wallace._0175_ ),
    .Y(\u_cpu.ALU.u_wallace._0298_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6113_  (.A1(\u_cpu.ALU.u_wallace._0295_ ),
    .A2(\u_cpu.ALU.u_wallace._0297_ ),
    .B1(\u_cpu.ALU.u_wallace._0298_ ),
    .Y(\u_cpu.ALU.u_wallace._0299_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6114_  (.A(\u_cpu.ALU.u_wallace._0295_ ),
    .B(\u_cpu.ALU.u_wallace._0297_ ),
    .C(\u_cpu.ALU.u_wallace._0298_ ),
    .X(\u_cpu.ALU.u_wallace._0300_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6115_  (.A(\u_cpu.ALU.u_wallace._0300_ ),
    .X(\u_cpu.ALU.u_wallace._0301_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._6116_  (.A1(\u_cpu.ALU.u_wallace._0200_ ),
    .A2(\u_cpu.ALU.u_wallace._3481_ ),
    .A3(\u_cpu.ALU.u_wallace._4698_ ),
    .B1(\u_cpu.ALU.u_wallace._0205_ ),
    .X(\u_cpu.ALU.u_wallace._0302_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._6117_  (.A1(\u_cpu.ALU.u_wallace._0299_ ),
    .A2(\u_cpu.ALU.u_wallace._0301_ ),
    .B1_N(\u_cpu.ALU.u_wallace._0302_ ),
    .Y(\u_cpu.ALU.u_wallace._0303_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6118_  (.A(\u_cpu.ALU.u_wallace._0200_ ),
    .B(\u_cpu.ALU.u_wallace._4542_ ),
    .C(\u_cpu.ALU.u_wallace._4698_ ),
    .X(\u_cpu.ALU.u_wallace._0305_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6119_  (.A1(\u_cpu.ALU.u_wallace._0295_ ),
    .A2(\u_cpu.ALU.u_wallace._0297_ ),
    .B1(\u_cpu.ALU.u_wallace._0298_ ),
    .X(\u_cpu.ALU.u_wallace._0306_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6120_  (.A(\u_cpu.ALU.u_wallace._4660_ ),
    .B(\u_cpu.ALU.u_wallace._3404_ ),
    .Y(\u_cpu.ALU.u_wallace._0307_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._6121_  (.A1(\u_cpu.ALU.u_wallace._1476_ ),
    .A2(\u_cpu.ALU.u_wallace._1508_ ),
    .A3(\u_cpu.ALU.u_wallace._4643_ ),
    .A4(\u_cpu.ALU.u_wallace._4798_ ),
    .B1(\u_cpu.ALU.u_wallace._0307_ ),
    .X(\u_cpu.ALU.u_wallace._0308_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6122_  (.A1(\u_cpu.ALU.u_wallace._0308_ ),
    .A2(\u_cpu.ALU.u_wallace._0292_ ),
    .B1(\u_cpu.ALU.u_wallace._0298_ ),
    .C1(\u_cpu.ALU.u_wallace._0297_ ),
    .Y(\u_cpu.ALU.u_wallace._0309_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6123_  (.A1(\u_cpu.ALU.u_wallace._0205_ ),
    .A2(\u_cpu.ALU.u_wallace._0305_ ),
    .B1(\u_cpu.ALU.u_wallace._0306_ ),
    .C1(\u_cpu.ALU.u_wallace._0309_ ),
    .Y(\u_cpu.ALU.u_wallace._0310_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._6124_  (.A(\u_cpu.ALU.u_wallace._4922_ ),
    .B(\u_cpu.ALU.u_wallace._0178_ ),
    .C(\u_cpu.ALU.u_wallace._0183_ ),
    .Y(\u_cpu.ALU.u_wallace._0311_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._6125_  (.A1(\u_cpu.ALU.u_wallace._0172_ ),
    .A2(\u_cpu.ALU.u_wallace._0176_ ),
    .A3(\u_cpu.ALU.u_wallace._0185_ ),
    .B1(\u_cpu.ALU.u_wallace._0311_ ),
    .X(\u_cpu.ALU.u_wallace._0312_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6126_  (.A(\u_cpu.ALU.SrcA[14] ),
    .X(\u_cpu.ALU.u_wallace._0313_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6127_  (.A1(\u_cpu.ALU.u_wallace._4658_ ),
    .A2(\u_cpu.ALU.u_wallace._4907_ ),
    .B1(\u_cpu.ALU.u_wallace._0313_ ),
    .B2(\u_cpu.ALU.u_wallace._4657_ ),
    .Y(\u_cpu.ALU.u_wallace._0314_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6128_  (.A(\u_cpu.ALU.u_wallace._0479_ ),
    .B(\u_cpu.ALU.u_wallace._1914_ ),
    .C(\u_cpu.ALU.u_wallace._4909_ ),
    .D(\u_cpu.ALU.u_wallace._0182_ ),
    .X(\u_cpu.ALU.u_wallace._0316_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6129_  (.A(\u_cpu.ALU.u_wallace._0457_ ),
    .B(\u_cpu.ALU.u_wallace._4785_ ),
    .Y(\u_cpu.ALU.u_wallace._0317_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6130_  (.A1(\u_cpu.ALU.u_wallace._0314_ ),
    .A2(\u_cpu.ALU.u_wallace._0316_ ),
    .B1(\u_cpu.ALU.u_wallace._0317_ ),
    .Y(\u_cpu.ALU.u_wallace._0318_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6131_  (.A(\u_cpu.ALU.u_wallace._4909_ ),
    .X(\u_cpu.ALU.u_wallace._0319_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6132_  (.A(\u_cpu.ALU.u_wallace._0182_ ),
    .X(\u_cpu.ALU.u_wallace._0320_ ));
 sky130_fd_sc_hd__a41oi_2 \u_cpu.ALU.u_wallace._6133_  (.A1(\u_cpu.ALU.u_wallace._0187_ ),
    .A2(\u_cpu.ALU.u_wallace._0304_ ),
    .A3(\u_cpu.ALU.u_wallace._0319_ ),
    .A4(\u_cpu.ALU.u_wallace._0320_ ),
    .B1(\u_cpu.ALU.u_wallace._0317_ ),
    .Y(\u_cpu.ALU.u_wallace._0321_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6134_  (.A1(\u_cpu.ALU.u_wallace._0545_ ),
    .A2(\u_cpu.ALU.u_wallace._4921_ ),
    .B1(\u_cpu.ALU.u_wallace._0179_ ),
    .B2(\u_cpu.ALU.u_wallace._0523_ ),
    .X(\u_cpu.ALU.u_wallace._0322_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6135_  (.A(\u_cpu.ALU.u_wallace._0321_ ),
    .B(\u_cpu.ALU.u_wallace._0322_ ),
    .Y(\u_cpu.ALU.u_wallace._0323_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6136_  (.A(\u_cpu.ALU.SrcA[15] ),
    .X(\u_cpu.ALU.u_wallace._0324_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6137_  (.A(\u_cpu.ALU.u_wallace._0324_ ),
    .X(\u_cpu.ALU.u_wallace._0325_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6138_  (.A1(\u_cpu.ALU.u_wallace._4431_ ),
    .A2(\u_cpu.ALU.u_wallace._4439_ ),
    .B1(\u_cpu.ALU.u_wallace._0325_ ),
    .B2(\u_cpu.ALU.u_wallace._1749_ ),
    .Y(\u_cpu.ALU.u_wallace._0327_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6139_  (.A(\u_cpu.ALU.u_wallace._0862_ ),
    .B(\u_cpu.ALU.u_wallace._2768_ ),
    .C(\u_cpu.ALU.u_wallace._4401_ ),
    .D(\u_cpu.ALU.u_wallace._0324_ ),
    .X(\u_cpu.ALU.u_wallace._0328_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6140_  (.A1(\u_cpu.ALU.u_wallace._0327_ ),
    .A2(\u_cpu.ALU.u_wallace._0328_ ),
    .B1(\u_cpu.ALU.u_wallace._0180_ ),
    .Y(\u_cpu.ALU.u_wallace._0329_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6141_  (.A(\u_cpu.ALU.SrcA[15] ),
    .X(\u_cpu.ALU.u_wallace._0330_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6142_  (.A1(\u_cpu.ALU.u_wallace._4645_ ),
    .A2(\u_cpu.ALU.u_wallace._4412_ ),
    .B1(\u_cpu.ALU.u_wallace._0330_ ),
    .B2(\u_cpu.ALU.u_wallace._0075_ ),
    .X(\u_cpu.ALU.u_wallace._0331_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6143_  (.A(\u_cpu.ALU.SrcA[15] ),
    .X(\u_cpu.ALU.u_wallace._0332_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6144_  (.A(\u_cpu.ALU.u_wallace._0075_ ),
    .B(\u_cpu.ALU.u_wallace._2856_ ),
    .C(\u_cpu.ALU.u_wallace._4562_ ),
    .D(\u_cpu.ALU.u_wallace._0332_ ),
    .Y(\u_cpu.ALU.u_wallace._0333_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6145_  (.A(\u_cpu.ALU.u_wallace._0183_ ),
    .B(\u_cpu.ALU.u_wallace._0331_ ),
    .C(\u_cpu.ALU.u_wallace._0333_ ),
    .Y(\u_cpu.ALU.u_wallace._0334_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6146_  (.A1(\u_cpu.ALU.u_wallace._0318_ ),
    .A2(\u_cpu.ALU.u_wallace._0323_ ),
    .B1(\u_cpu.ALU.u_wallace._0329_ ),
    .B2(\u_cpu.ALU.u_wallace._0334_ ),
    .X(\u_cpu.ALU.u_wallace._0335_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._6147_  (.A1(\u_cpu.ALU.u_wallace._0217_ ),
    .A2(\u_cpu.ALU.u_wallace._4796_ ),
    .A3(\u_cpu.ALU.u_wallace._0319_ ),
    .A4(\u_cpu.ALU.u_wallace._0320_ ),
    .B1(\u_cpu.ALU.u_wallace._0317_ ),
    .X(\u_cpu.ALU.u_wallace._0336_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._6148_  (.A1(\u_cpu.ALU.u_wallace._0314_ ),
    .A2(\u_cpu.ALU.u_wallace._0336_ ),
    .B1(\u_cpu.ALU.u_wallace._0329_ ),
    .C1(\u_cpu.ALU.u_wallace._0334_ ),
    .D1(\u_cpu.ALU.u_wallace._0318_ ),
    .Y(\u_cpu.ALU.u_wallace._0338_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6149_  (.A(\u_cpu.ALU.u_wallace._0312_ ),
    .B(\u_cpu.ALU.u_wallace._0335_ ),
    .C(\u_cpu.ALU.u_wallace._0338_ ),
    .Y(\u_cpu.ALU.u_wallace._0339_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6150_  (.A1(\u_cpu.ALU.u_wallace._0318_ ),
    .A2(\u_cpu.ALU.u_wallace._0323_ ),
    .B1(\u_cpu.ALU.u_wallace._0329_ ),
    .B2(\u_cpu.ALU.u_wallace._0334_ ),
    .Y(\u_cpu.ALU.u_wallace._0340_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._6151_  (.A1(\u_cpu.ALU.u_wallace._0314_ ),
    .A2(\u_cpu.ALU.u_wallace._0336_ ),
    .B1(\u_cpu.ALU.u_wallace._0329_ ),
    .C1(\u_cpu.ALU.u_wallace._0334_ ),
    .D1(\u_cpu.ALU.u_wallace._0318_ ),
    .X(\u_cpu.ALU.u_wallace._0341_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._6152_  (.A1(\u_cpu.ALU.u_wallace._0172_ ),
    .A2(\u_cpu.ALU.u_wallace._0176_ ),
    .A3(\u_cpu.ALU.u_wallace._0185_ ),
    .B1(\u_cpu.ALU.u_wallace._0311_ ),
    .Y(\u_cpu.ALU.u_wallace._0342_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6153_  (.A1(\u_cpu.ALU.u_wallace._0340_ ),
    .A2(\u_cpu.ALU.u_wallace._0341_ ),
    .B1(\u_cpu.ALU.u_wallace._0342_ ),
    .Y(\u_cpu.ALU.u_wallace._0343_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6154_  (.A1(\u_cpu.ALU.u_wallace._0303_ ),
    .A2(\u_cpu.ALU.u_wallace._0310_ ),
    .B1(\u_cpu.ALU.u_wallace._0339_ ),
    .B2(\u_cpu.ALU.u_wallace._0343_ ),
    .X(\u_cpu.ALU.u_wallace._0344_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._6155_  (.A1(\u_cpu.ALU.u_wallace._4678_ ),
    .A2(\u_cpu.ALU.u_wallace._0169_ ),
    .A3(\u_cpu.ALU.u_wallace._0170_ ),
    .B1(\u_cpu.ALU.u_wallace._0175_ ),
    .X(\u_cpu.ALU.u_wallace._0345_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6156_  (.A1(\u_cpu.ALU.u_wallace._0292_ ),
    .A2(\u_cpu.ALU.u_wallace._0308_ ),
    .B1(\u_cpu.ALU.u_wallace._0297_ ),
    .Y(\u_cpu.ALU.u_wallace._0346_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6157_  (.A1_N(\u_cpu.ALU.u_wallace._0345_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0346_ ),
    .B1(\u_cpu.ALU.u_wallace._0305_ ),
    .B2(\u_cpu.ALU.u_wallace._0205_ ),
    .Y(\u_cpu.ALU.u_wallace._0347_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._6158_  (.A1(\u_cpu.ALU.u_wallace._0347_ ),
    .A2(\u_cpu.ALU.u_wallace._0301_ ),
    .B1(\u_cpu.ALU.u_wallace._0303_ ),
    .C1(\u_cpu.ALU.u_wallace._0339_ ),
    .D1(\u_cpu.ALU.u_wallace._0343_ ),
    .Y(\u_cpu.ALU.u_wallace._0349_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6159_  (.A(\u_cpu.ALU.u_wallace._0197_ ),
    .B(\u_cpu.ALU.u_wallace._0223_ ),
    .C(\u_cpu.ALU.u_wallace._0224_ ),
    .Y(\u_cpu.ALU.u_wallace._0350_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6160_  (.A(\u_cpu.ALU.u_wallace._0192_ ),
    .B(\u_cpu.ALU.u_wallace._0350_ ),
    .Y(\u_cpu.ALU.u_wallace._0351_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6161_  (.A1(\u_cpu.ALU.u_wallace._0344_ ),
    .A2(\u_cpu.ALU.u_wallace._0349_ ),
    .B1(\u_cpu.ALU.u_wallace._0351_ ),
    .Y(\u_cpu.ALU.u_wallace._0352_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6162_  (.A1(\u_cpu.ALU.u_wallace._0218_ ),
    .A2(\u_cpu.ALU.u_wallace._0216_ ),
    .B1(\u_cpu.ALU.u_wallace._0221_ ),
    .Y(\u_cpu.ALU.u_wallace._0353_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6163_  (.A1(\u_cpu.ALU.u_wallace._2878_ ),
    .A2(\u_cpu.ALU.u_wallace._4007_ ),
    .B1(\u_cpu.ALU.u_wallace._4291_ ),
    .B2(\u_cpu.ALU.u_wallace._1837_ ),
    .Y(\u_cpu.ALU.u_wallace._0354_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6164_  (.A(\u_cpu.ALU.u_wallace._2790_ ),
    .B(\u_cpu.ALU.u_wallace._1837_ ),
    .C(\u_cpu.ALU.u_wallace._4007_ ),
    .D(\u_cpu.ALU.u_wallace._4291_ ),
    .X(\u_cpu.ALU.u_wallace._0355_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6165_  (.A(\u_cpu.ALU.u_wallace._4529_ ),
    .B(\u_cpu.ALU.u_wallace._4609_ ),
    .Y(\u_cpu.ALU.u_wallace._0356_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6166_  (.A1(\u_cpu.ALU.u_wallace._0354_ ),
    .A2(\u_cpu.ALU.u_wallace._0355_ ),
    .B1(\u_cpu.ALU.u_wallace._0356_ ),
    .Y(\u_cpu.ALU.u_wallace._0357_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6167_  (.A(\u_cpu.ALU.u_wallace._4447_ ),
    .B(\u_cpu.ALU.u_wallace._2834_ ),
    .C(\u_cpu.ALU.u_wallace._4847_ ),
    .D(\u_cpu.ALU.u_wallace._0045_ ),
    .Y(\u_cpu.ALU.u_wallace._0358_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._6168_  (.A_N(\u_cpu.ALU.u_wallace._0354_ ),
    .B(\u_cpu.ALU.u_wallace._0358_ ),
    .C(\u_cpu.ALU.u_wallace._1322_ ),
    .D(\u_cpu.ALU.u_wallace._4604_ ),
    .Y(\u_cpu.ALU.u_wallace._0360_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6169_  (.A1(\u_cpu.ALU.u_wallace._0133_ ),
    .A2(\u_cpu.ALU.u_wallace._0135_ ),
    .B1(\u_cpu.ALU.u_wallace._0141_ ),
    .Y(\u_cpu.ALU.u_wallace._0361_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6170_  (.A1(\u_cpu.ALU.u_wallace._0357_ ),
    .A2(\u_cpu.ALU.u_wallace._0360_ ),
    .B1(\u_cpu.ALU.u_wallace._0361_ ),
    .X(\u_cpu.ALU.u_wallace._0362_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6171_  (.A(\u_cpu.ALU.SrcB[13] ),
    .X(\u_cpu.ALU.u_wallace._0363_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6172_  (.A(\u_cpu.ALU.SrcB[11] ),
    .X(\u_cpu.ALU.u_wallace._0364_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6173_  (.A(\u_cpu.ALU.SrcB[12] ),
    .X(\u_cpu.ALU.u_wallace._0365_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6174_  (.A1(\u_cpu.ALU.u_wallace._2922_ ),
    .A2(\u_cpu.ALU.u_wallace._0364_ ),
    .B1(\u_cpu.ALU.u_wallace._0365_ ),
    .B2(\u_cpu.ALU.u_wallace._0600_ ),
    .X(\u_cpu.ALU.u_wallace._0366_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6175_  (.A(\u_cpu.ALU.u_wallace._1267_ ),
    .B(\u_cpu.ALU.u_wallace._1278_ ),
    .C(\u_cpu.ALU.u_wallace._4731_ ),
    .D(\u_cpu.ALU.u_wallace._0144_ ),
    .Y(\u_cpu.ALU.u_wallace._0367_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6176_  (.A1(\u_cpu.ALU.u_wallace._0359_ ),
    .A2(\u_cpu.ALU.u_wallace._0363_ ),
    .B1(\u_cpu.ALU.u_wallace._0366_ ),
    .B2(\u_cpu.ALU.u_wallace._0367_ ),
    .Y(\u_cpu.ALU.u_wallace._0368_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6177_  (.A(\u_cpu.ALU.u_wallace._0366_ ),
    .B(\u_cpu.ALU.u_wallace._0367_ ),
    .C(\u_cpu.ALU.u_wallace._4597_ ),
    .D(\u_cpu.ALU.u_wallace._0363_ ),
    .X(\u_cpu.ALU.u_wallace._0369_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._6178_  (.A(\u_cpu.ALU.u_wallace._0368_ ),
    .B(\u_cpu.ALU.u_wallace._0369_ ),
    .Y(\u_cpu.ALU.u_wallace._0371_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._6179_  (.A(\u_cpu.ALU.u_wallace._0133_ ),
    .B(\u_cpu.ALU.u_wallace._0135_ ),
    .Y(\u_cpu.ALU.u_wallace._0372_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6180_  (.A1(\u_cpu.ALU.u_wallace._0137_ ),
    .A2(\u_cpu.ALU.u_wallace._0372_ ),
    .B1(\u_cpu.ALU.u_wallace._0360_ ),
    .C1(\u_cpu.ALU.u_wallace._0357_ ),
    .Y(\u_cpu.ALU.u_wallace._0373_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6181_  (.A(\u_cpu.ALU.u_wallace._0362_ ),
    .B(\u_cpu.ALU.u_wallace._0371_ ),
    .C(\u_cpu.ALU.u_wallace._0373_ ),
    .Y(\u_cpu.ALU.u_wallace._0374_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6182_  (.A1(\u_cpu.ALU.u_wallace._0137_ ),
    .A2(\u_cpu.ALU.u_wallace._0372_ ),
    .B1(\u_cpu.ALU.u_wallace._0360_ ),
    .C1(\u_cpu.ALU.u_wallace._0357_ ),
    .X(\u_cpu.ALU.u_wallace._0375_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6183_  (.A1(\u_cpu.ALU.u_wallace._0357_ ),
    .A2(\u_cpu.ALU.u_wallace._0360_ ),
    .B1(\u_cpu.ALU.u_wallace._0361_ ),
    .Y(\u_cpu.ALU.u_wallace._0376_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6184_  (.A1(\u_cpu.ALU.u_wallace._0368_ ),
    .A2(\u_cpu.ALU.u_wallace._0369_ ),
    .B1(\u_cpu.ALU.u_wallace._0375_ ),
    .B2(\u_cpu.ALU.u_wallace._0376_ ),
    .Y(\u_cpu.ALU.u_wallace._0377_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6185_  (.A(\u_cpu.ALU.u_wallace._0353_ ),
    .B(\u_cpu.ALU.u_wallace._0374_ ),
    .C(\u_cpu.ALU.u_wallace._0377_ ),
    .X(\u_cpu.ALU.u_wallace._0378_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._6186_  (.A1(\u_cpu.ALU.u_wallace._0218_ ),
    .A2(\u_cpu.ALU.u_wallace._0216_ ),
    .B1(\u_cpu.ALU.u_wallace._0221_ ),
    .X(\u_cpu.ALU.u_wallace._0379_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6187_  (.A1(\u_cpu.ALU.u_wallace._0375_ ),
    .A2(\u_cpu.ALU.u_wallace._0376_ ),
    .B1(\u_cpu.ALU.u_wallace._0371_ ),
    .Y(\u_cpu.ALU.u_wallace._0380_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6188_  (.A1(\u_cpu.ALU.u_wallace._0368_ ),
    .A2(\u_cpu.ALU.u_wallace._0369_ ),
    .B1(\u_cpu.ALU.u_wallace._0373_ ),
    .C1(\u_cpu.ALU.u_wallace._0362_ ),
    .Y(\u_cpu.ALU.u_wallace._0382_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._6189_  (.A1(\u_cpu.ALU.u_wallace._0147_ ),
    .A2(\u_cpu.ALU.u_wallace._0148_ ),
    .A3(\u_cpu.ALU.u_wallace._0143_ ),
    .B1(\u_cpu.ALU.u_wallace._0152_ ),
    .X(\u_cpu.ALU.u_wallace._0383_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._6190_  (.A1(\u_cpu.ALU.u_wallace._0379_ ),
    .A2(\u_cpu.ALU.u_wallace._0380_ ),
    .A3(\u_cpu.ALU.u_wallace._0382_ ),
    .B1(\u_cpu.ALU.u_wallace._0383_ ),
    .X(\u_cpu.ALU.u_wallace._0384_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6191_  (.A(\u_cpu.ALU.u_wallace._0379_ ),
    .B(\u_cpu.ALU.u_wallace._0380_ ),
    .C(\u_cpu.ALU.u_wallace._0382_ ),
    .Y(\u_cpu.ALU.u_wallace._0385_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6192_  (.A(\u_cpu.ALU.u_wallace._0353_ ),
    .B(\u_cpu.ALU.u_wallace._0374_ ),
    .C(\u_cpu.ALU.u_wallace._0377_ ),
    .Y(\u_cpu.ALU.u_wallace._0386_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._6193_  (.A1(\u_cpu.ALU.u_wallace._0136_ ),
    .A2(\u_cpu.ALU.u_wallace._0138_ ),
    .A3(\u_cpu.ALU.u_wallace._0142_ ),
    .B1(\u_cpu.ALU.u_wallace._0153_ ),
    .B2(\u_cpu.ALU.u_wallace._0149_ ),
    .X(\u_cpu.ALU.u_wallace._0387_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6194_  (.A1(\u_cpu.ALU.u_wallace._0385_ ),
    .A2(\u_cpu.ALU.u_wallace._0386_ ),
    .B1(\u_cpu.ALU.u_wallace._0387_ ),
    .X(\u_cpu.ALU.u_wallace._0388_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6195_  (.A(\u_cpu.ALU.u_wallace._0351_ ),
    .B(\u_cpu.ALU.u_wallace._0344_ ),
    .C(\u_cpu.ALU.u_wallace._0349_ ),
    .Y(\u_cpu.ALU.u_wallace._0389_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6196_  (.A1(\u_cpu.ALU.u_wallace._0378_ ),
    .A2(\u_cpu.ALU.u_wallace._0384_ ),
    .B1(\u_cpu.ALU.u_wallace._0388_ ),
    .C1(\u_cpu.ALU.u_wallace._0389_ ),
    .Y(\u_cpu.ALU.u_wallace._0390_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6197_  (.A1(\u_cpu.ALU.u_wallace._0303_ ),
    .A2(\u_cpu.ALU.u_wallace._0310_ ),
    .B1(\u_cpu.ALU.u_wallace._0339_ ),
    .B2(\u_cpu.ALU.u_wallace._0343_ ),
    .Y(\u_cpu.ALU.u_wallace._0391_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._6198_  (.A1(\u_cpu.ALU.u_wallace._0347_ ),
    .A2(\u_cpu.ALU.u_wallace._0301_ ),
    .B1(\u_cpu.ALU.u_wallace._0303_ ),
    .C1(\u_cpu.ALU.u_wallace._0339_ ),
    .D1(\u_cpu.ALU.u_wallace._0343_ ),
    .X(\u_cpu.ALU.u_wallace._0393_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._6199_  (.A1(\u_cpu.ALU.u_wallace._0196_ ),
    .A2(\u_cpu.ALU.u_wallace._0193_ ),
    .A3(\u_cpu.ALU.u_wallace._0194_ ),
    .B1(\u_cpu.ALU.u_wallace._0350_ ),
    .X(\u_cpu.ALU.u_wallace._0394_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6200_  (.A1(\u_cpu.ALU.u_wallace._0391_ ),
    .A2(\u_cpu.ALU.u_wallace._0393_ ),
    .B1(\u_cpu.ALU.u_wallace._0394_ ),
    .Y(\u_cpu.ALU.u_wallace._0395_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6201_  (.A1(\u_cpu.ALU.u_wallace._0385_ ),
    .A2(\u_cpu.ALU.u_wallace._0386_ ),
    .B1(\u_cpu.ALU.u_wallace._0387_ ),
    .Y(\u_cpu.ALU.u_wallace._0396_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6202_  (.A(\u_cpu.ALU.u_wallace._0387_ ),
    .B(\u_cpu.ALU.u_wallace._0385_ ),
    .C(\u_cpu.ALU.u_wallace._0386_ ),
    .Y(\u_cpu.ALU.u_wallace._0397_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._6203_  (.A(\u_cpu.ALU.u_wallace._0397_ ),
    .Y(\u_cpu.ALU.u_wallace._0398_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6204_  (.A1_N(\u_cpu.ALU.u_wallace._0395_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0389_ ),
    .B1(\u_cpu.ALU.u_wallace._0396_ ),
    .B2(\u_cpu.ALU.u_wallace._0398_ ),
    .Y(\u_cpu.ALU.u_wallace._0399_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._6205_  (.A1(\u_cpu.ALU.u_wallace._0072_ ),
    .A2(\u_cpu.ALU.u_wallace._0167_ ),
    .B1(\u_cpu.ALU.u_wallace._0225_ ),
    .X(\u_cpu.ALU.u_wallace._0400_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6206_  (.A(\u_cpu.ALU.u_wallace._0230_ ),
    .B(\u_cpu.ALU.u_wallace._0231_ ),
    .Y(\u_cpu.ALU.u_wallace._0401_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6207_  (.A1_N(\u_cpu.ALU.u_wallace._0220_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0400_ ),
    .B1(\u_cpu.ALU.u_wallace._0227_ ),
    .B2(\u_cpu.ALU.u_wallace._0401_ ),
    .Y(\u_cpu.ALU.u_wallace._0402_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6208_  (.A1(\u_cpu.ALU.u_wallace._0352_ ),
    .A2(\u_cpu.ALU.u_wallace._0390_ ),
    .B1(\u_cpu.ALU.u_wallace._0399_ ),
    .C1(\u_cpu.ALU.u_wallace._0402_ ),
    .X(\u_cpu.ALU.u_wallace._0404_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._6209_  (.A1(\u_cpu.ALU.u_wallace._0378_ ),
    .A2(\u_cpu.ALU.u_wallace._0384_ ),
    .B1(\u_cpu.ALU.u_wallace._0388_ ),
    .C1(\u_cpu.ALU.u_wallace._0395_ ),
    .D1(\u_cpu.ALU.u_wallace._0389_ ),
    .Y(\u_cpu.ALU.u_wallace._0405_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6210_  (.A1(\u_cpu.ALU.u_wallace._0399_ ),
    .A2(\u_cpu.ALU.u_wallace._0405_ ),
    .B1(\u_cpu.ALU.u_wallace._0402_ ),
    .Y(\u_cpu.ALU.u_wallace._0406_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6211_  (.A1(\u_cpu.ALU.u_wallace._0290_ ),
    .A2(\u_cpu.ALU.u_wallace._0291_ ),
    .B1(\u_cpu.ALU.u_wallace._0404_ ),
    .B2(\u_cpu.ALU.u_wallace._0406_ ),
    .Y(\u_cpu.ALU.u_wallace._0407_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6212_  (.A1(\u_cpu.ALU.u_wallace._0159_ ),
    .A2(\u_cpu.ALU.u_wallace._0231_ ),
    .B1(\u_cpu.ALU.u_wallace._0289_ ),
    .X(\u_cpu.ALU.u_wallace._0408_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6213_  (.A(\u_cpu.ALU.u_wallace._0159_ ),
    .B(\u_cpu.ALU.u_wallace._0231_ ),
    .C(\u_cpu.ALU.u_wallace._0289_ ),
    .Y(\u_cpu.ALU.u_wallace._0409_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6214_  (.A(\u_cpu.ALU.u_wallace._0408_ ),
    .B(\u_cpu.ALU.u_wallace._0409_ ),
    .Y(\u_cpu.ALU.u_wallace._0410_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6215_  (.A1(\u_cpu.ALU.u_wallace._0352_ ),
    .A2(\u_cpu.ALU.u_wallace._0390_ ),
    .B1(\u_cpu.ALU.u_wallace._0399_ ),
    .C1(\u_cpu.ALU.u_wallace._0402_ ),
    .Y(\u_cpu.ALU.u_wallace._0411_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6216_  (.A1(\u_cpu.ALU.u_wallace._0399_ ),
    .A2(\u_cpu.ALU.u_wallace._0405_ ),
    .B1(\u_cpu.ALU.u_wallace._0402_ ),
    .X(\u_cpu.ALU.u_wallace._0412_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6217_  (.A(\u_cpu.ALU.u_wallace._0410_ ),
    .B(\u_cpu.ALU.u_wallace._0411_ ),
    .C(\u_cpu.ALU.u_wallace._0412_ ),
    .Y(\u_cpu.ALU.u_wallace._0413_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6218_  (.A(\u_cpu.ALU.u_wallace._0276_ ),
    .B(\u_cpu.ALU.u_wallace._0407_ ),
    .C(\u_cpu.ALU.u_wallace._0413_ ),
    .Y(\u_cpu.ALU.u_wallace._0415_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6219_  (.A1(\u_cpu.ALU.u_wallace._0131_ ),
    .A2(\u_cpu.ALU.u_wallace._0245_ ),
    .B1(\u_cpu.ALU.u_wallace._0242_ ),
    .Y(\u_cpu.ALU.u_wallace._0416_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6220_  (.A1(\u_cpu.ALU.u_wallace._0290_ ),
    .A2(\u_cpu.ALU.u_wallace._0291_ ),
    .B1(\u_cpu.ALU.u_wallace._0411_ ),
    .C1(\u_cpu.ALU.u_wallace._0412_ ),
    .Y(\u_cpu.ALU.u_wallace._0417_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6221_  (.A1_N(\u_cpu.ALU.u_wallace._0408_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0409_ ),
    .B1(\u_cpu.ALU.u_wallace._0404_ ),
    .B2(\u_cpu.ALU.u_wallace._0406_ ),
    .Y(\u_cpu.ALU.u_wallace._0418_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6222_  (.A(\u_cpu.ALU.u_wallace._0416_ ),
    .B(\u_cpu.ALU.u_wallace._0417_ ),
    .C(\u_cpu.ALU.u_wallace._0418_ ),
    .Y(\u_cpu.ALU.u_wallace._0419_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._6223_  (.A(\u_cpu.ALU.u_wallace._0066_ ),
    .B(\u_cpu.ALU.u_wallace._0070_ ),
    .X(\u_cpu.ALU.u_wallace._0420_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6224_  (.A1_N(\u_cpu.ALU.u_wallace._0415_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0419_ ),
    .B1(\u_cpu.ALU.u_wallace._0420_ ),
    .B2(\u_cpu.ALU.u_wallace._0127_ ),
    .Y(\u_cpu.ALU.u_wallace._0421_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6225_  (.A(\u_cpu.ALU.u_wallace._0419_ ),
    .B(\u_cpu.ALU.u_wallace._0128_ ),
    .C(\u_cpu.ALU.u_wallace._0415_ ),
    .Y(\u_cpu.ALU.u_wallace._0422_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6226_  (.A1(\u_cpu.ALU.u_wallace._0252_ ),
    .A2(\u_cpu.ALU.u_wallace._0260_ ),
    .B1(\u_cpu.ALU.u_wallace._0248_ ),
    .Y(\u_cpu.ALU.u_wallace._0423_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6227_  (.A1(\u_cpu.ALU.u_wallace._0421_ ),
    .A2(\u_cpu.ALU.u_wallace._0422_ ),
    .B1(\u_cpu.ALU.u_wallace._0423_ ),
    .Y(\u_cpu.ALU.u_wallace._0424_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6228_  (.A1(\u_cpu.ALU.u_wallace._0258_ ),
    .A2(\u_cpu.ALU.u_wallace._0253_ ),
    .B1(\u_cpu.ALU.u_wallace._0421_ ),
    .C1(\u_cpu.ALU.u_wallace._0422_ ),
    .X(\u_cpu.ALU.u_wallace._0426_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6229_  (.A(\u_cpu.ALU.u_wallace._0262_ ),
    .B(\u_cpu.ALU.u_wallace._0264_ ),
    .C(\u_cpu.ALU.u_wallace._0259_ ),
    .Y(\u_cpu.ALU.u_wallace._0427_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6230_  (.A1(\u_cpu.ALU.u_wallace._0424_ ),
    .A2(\u_cpu.ALU.u_wallace._0426_ ),
    .B1(\u_cpu.ALU.u_wallace._0427_ ),
    .Y(\u_cpu.ALU.u_wallace._0428_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6231_  (.A1(\u_cpu.ALU.u_wallace._0421_ ),
    .A2(\u_cpu.ALU.u_wallace._0422_ ),
    .B1(\u_cpu.ALU.u_wallace._0423_ ),
    .X(\u_cpu.ALU.u_wallace._0429_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6232_  (.A(\u_cpu.ALU.u_wallace._0259_ ),
    .B(\u_cpu.ALU.u_wallace._0262_ ),
    .C(\u_cpu.ALU.u_wallace._0429_ ),
    .D(\u_cpu.ALU.u_wallace._0264_ ),
    .Y(\u_cpu.ALU.u_wallace._0430_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6233_  (.A1(\u_cpu.ALU.u_wallace._0428_ ),
    .A2(\u_cpu.ALU.u_wallace._0430_ ),
    .B1(\u_cpu.ALU.u_wallace._0275_ ),
    .Y(\u_cpu.ALU.u_wallace._0431_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6234_  (.A1(\u_cpu.ALU.u_wallace._0275_ ),
    .A2(\u_cpu.ALU.u_wallace._0428_ ),
    .B1(\u_cpu.ALU.u_wallace._0431_ ),
    .Y(\u_cpu.ALU.u_wallace._0432_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.ALU.u_wallace._6235_  (.A1(\u_cpu.ALU.u_wallace._0107_ ),
    .A2(\u_cpu.ALU.u_wallace._0266_ ),
    .A3(\u_cpu.ALU.u_wallace._0114_ ),
    .B1(\u_cpu.ALU.u_wallace._0274_ ),
    .B2(\u_cpu.ALU.u_wallace._0270_ ),
    .X(\u_cpu.ALU.u_wallace._0433_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu.ALU.u_wallace._6236_  (.A(\u_cpu.ALU.u_wallace._0432_ ),
    .B(\u_cpu.ALU.u_wallace._0433_ ),
    .Y(\u_cpu.ALU.Product_Wallace[15] ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6237_  (.A1(\u_cpu.ALU.u_wallace._0258_ ),
    .A2(\u_cpu.ALU.u_wallace._0253_ ),
    .B1(\u_cpu.ALU.u_wallace._0421_ ),
    .C1(\u_cpu.ALU.u_wallace._0422_ ),
    .Y(\u_cpu.ALU.u_wallace._0434_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._6238_  (.A1(\u_cpu.ALU.u_wallace._0427_ ),
    .A2(\u_cpu.ALU.u_wallace._0424_ ),
    .B1(\u_cpu.ALU.u_wallace._0434_ ),
    .X(\u_cpu.ALU.u_wallace._0436_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6239_  (.A1(\u_cpu.ALU.u_wallace._0410_ ),
    .A2(\u_cpu.ALU.u_wallace._0406_ ),
    .B1(\u_cpu.ALU.u_wallace._0411_ ),
    .Y(\u_cpu.ALU.u_wallace._0437_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6240_  (.A(\u_cpu.ALU.u_wallace._0742_ ),
    .B(\u_cpu.ALU.u_wallace._4909_ ),
    .Y(\u_cpu.ALU.u_wallace._0438_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._6241_  (.A1(\u_cpu.ALU.u_wallace._0523_ ),
    .A2(\u_cpu.ALU.u_wallace._0545_ ),
    .A3(\u_cpu.ALU.u_wallace._0313_ ),
    .A4(\u_cpu.ALU.u_wallace._0325_ ),
    .B1(\u_cpu.ALU.u_wallace._0438_ ),
    .X(\u_cpu.ALU.u_wallace._0439_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6242_  (.A1(\u_cpu.ALU.u_wallace._1968_ ),
    .A2(\u_cpu.ALU.u_wallace._0313_ ),
    .B1(\u_cpu.ALU.u_wallace._0325_ ),
    .B2(\u_cpu.ALU.u_wallace._1957_ ),
    .Y(\u_cpu.ALU.u_wallace._0440_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6243_  (.A(\u_cpu.ALU.SrcA[16] ),
    .X(\u_cpu.ALU.u_wallace._0441_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._6244_  (.A(\u_cpu.ALU.u_wallace._0441_ ),
    .Y(\u_cpu.ALU.u_wallace._0442_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6245_  (.A(\u_cpu.ALU.u_wallace._1749_ ),
    .B(\u_cpu.ALU.u_wallace._1771_ ),
    .C(\u_cpu.ALU.u_wallace._4557_ ),
    .Y(\u_cpu.ALU.u_wallace._0443_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6246_  (.A1(\u_cpu.ALU.u_wallace._3678_ ),
    .A2(\u_cpu.ALU.u_wallace._4553_ ),
    .B1(\u_cpu.ALU.u_wallace._0441_ ),
    .B2(\u_cpu.ALU.u_wallace._0862_ ),
    .X(\u_cpu.ALU.u_wallace._0444_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6247_  (.A1(\u_cpu.ALU.u_wallace._0442_ ),
    .A2(\u_cpu.ALU.u_wallace._0443_ ),
    .B1(\u_cpu.ALU.u_wallace._0444_ ),
    .C1(\u_cpu.ALU.u_wallace._0328_ ),
    .Y(\u_cpu.ALU.u_wallace._0445_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6248_  (.A(\u_cpu.ALU.SrcA[16] ),
    .X(\u_cpu.ALU.u_wallace._0447_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6249_  (.A(\u_cpu.ALU.u_wallace._0447_ ),
    .X(\u_cpu.ALU.u_wallace._0448_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6250_  (.A1(\u_cpu.ALU.u_wallace._3678_ ),
    .A2(\u_cpu.ALU.u_wallace._4553_ ),
    .B1(\u_cpu.ALU.u_wallace._0448_ ),
    .B2(\u_cpu.ALU.u_wallace._0862_ ),
    .Y(\u_cpu.ALU.u_wallace._0449_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6251_  (.A(\u_cpu.ALU.SrcB[0] ),
    .B(\u_cpu.ALU.SrcB[6] ),
    .C(\u_cpu.ALU.SrcA[10] ),
    .D(\u_cpu.ALU.SrcA[16] ),
    .X(\u_cpu.ALU.u_wallace._0450_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6252_  (.A(\u_cpu.ALU.u_wallace._0450_ ),
    .X(\u_cpu.ALU.u_wallace._0451_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6253_  (.A1(\u_cpu.ALU.u_wallace._0449_ ),
    .A2(\u_cpu.ALU.u_wallace._0451_ ),
    .B1(\u_cpu.ALU.u_wallace._0333_ ),
    .Y(\u_cpu.ALU.u_wallace._0452_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6254_  (.A1(\u_cpu.ALU.u_wallace._0293_ ),
    .A2(\u_cpu.ALU.SrcA[14] ),
    .B1(\u_cpu.ALU.u_wallace._0324_ ),
    .B2(\u_cpu.ALU.u_wallace._0797_ ),
    .X(\u_cpu.ALU.u_wallace._0453_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6255_  (.A(\u_cpu.ALU.u_wallace._0479_ ),
    .B(\u_cpu.ALU.u_wallace._0807_ ),
    .C(\u_cpu.ALU.u_wallace._0182_ ),
    .D(\u_cpu.ALU.u_wallace._0332_ ),
    .Y(\u_cpu.ALU.u_wallace._0454_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6256_  (.A1(\u_cpu.ALU.u_wallace._0753_ ),
    .A2(\u_cpu.ALU.u_wallace._0188_ ),
    .B1(\u_cpu.ALU.u_wallace._0453_ ),
    .B2(\u_cpu.ALU.u_wallace._0454_ ),
    .X(\u_cpu.ALU.u_wallace._0455_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._6257_  (.A1(\u_cpu.ALU.u_wallace._0439_ ),
    .A2(\u_cpu.ALU.u_wallace._0440_ ),
    .B1(\u_cpu.ALU.u_wallace._0445_ ),
    .C1(\u_cpu.ALU.u_wallace._0452_ ),
    .D1(\u_cpu.ALU.u_wallace._0455_ ),
    .Y(\u_cpu.ALU.u_wallace._0456_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._6258_  (.A(\u_cpu.ALU.u_wallace._4920_ ),
    .Y(\u_cpu.ALU.u_wallace._0458_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6259_  (.A(\u_cpu.ALU.u_wallace._4657_ ),
    .B(\u_cpu.ALU.u_wallace._4658_ ),
    .C(\u_cpu.ALU.u_wallace._0177_ ),
    .D(\u_cpu.ALU.u_wallace._0330_ ),
    .X(\u_cpu.ALU.u_wallace._0459_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._6260_  (.A1(\u_cpu.ALU.u_wallace._1892_ ),
    .A2(\u_cpu.ALU.u_wallace._0458_ ),
    .B1(\u_cpu.ALU.u_wallace._0440_ ),
    .B2(\u_cpu.ALU.u_wallace._0459_ ),
    .X(\u_cpu.ALU.u_wallace._0460_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6261_  (.A(\u_cpu.ALU.u_wallace._0453_ ),
    .B(\u_cpu.ALU.u_wallace._0454_ ),
    .C(\u_cpu.ALU.u_wallace._4662_ ),
    .D(\u_cpu.ALU.u_wallace._0319_ ),
    .X(\u_cpu.ALU.u_wallace._0461_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6262_  (.A1_N(\u_cpu.ALU.u_wallace._0452_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0445_ ),
    .B1(\u_cpu.ALU.u_wallace._0460_ ),
    .B2(\u_cpu.ALU.u_wallace._0461_ ),
    .Y(\u_cpu.ALU.u_wallace._0462_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6263_  (.A(\u_cpu.ALU.u_wallace._0183_ ),
    .B(\u_cpu.ALU.u_wallace._0331_ ),
    .C(\u_cpu.ALU.u_wallace._0333_ ),
    .X(\u_cpu.ALU.u_wallace._0463_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._6264_  (.A1(\u_cpu.ALU.u_wallace._0318_ ),
    .A2(\u_cpu.ALU.u_wallace._0323_ ),
    .A3(\u_cpu.ALU.u_wallace._0329_ ),
    .B1(\u_cpu.ALU.u_wallace._0463_ ),
    .X(\u_cpu.ALU.u_wallace._0464_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6265_  (.A1(\u_cpu.ALU.u_wallace._0456_ ),
    .A2(\u_cpu.ALU.u_wallace._0462_ ),
    .B1(\u_cpu.ALU.u_wallace._0464_ ),
    .Y(\u_cpu.ALU.u_wallace._0465_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6266_  (.A(\u_cpu.ALU.u_wallace._0464_ ),
    .B(\u_cpu.ALU.u_wallace._0456_ ),
    .C(\u_cpu.ALU.u_wallace._0462_ ),
    .Y(\u_cpu.ALU.u_wallace._0466_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._6267_  (.A1(\u_cpu.ALU.u_wallace._4677_ ),
    .A2(\u_cpu.ALU.u_wallace._4539_ ),
    .A3(\u_cpu.ALU.u_wallace._0292_ ),
    .B1(\u_cpu.ALU.u_wallace._0294_ ),
    .X(\u_cpu.ALU.u_wallace._0467_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._6268_  (.A(\u_cpu.ALU.u_wallace._0317_ ),
    .B(\u_cpu.ALU.u_wallace._0314_ ),
    .Y(\u_cpu.ALU.u_wallace._0469_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6269_  (.A1(\u_cpu.ALU.u_wallace._2582_ ),
    .A2(\u_cpu.ALU.u_wallace._4647_ ),
    .B1(\u_cpu.ALU.u_wallace._4785_ ),
    .B2(\u_cpu.ALU.u_wallace._2571_ ),
    .X(\u_cpu.ALU.u_wallace._0470_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6270_  (.A(\u_cpu.ALU.u_wallace._1530_ ),
    .B(\u_cpu.ALU.u_wallace._1552_ ),
    .C(\u_cpu.ALU.u_wallace._4794_ ),
    .D(\u_cpu.ALU.u_wallace._4917_ ),
    .Y(\u_cpu.ALU.u_wallace._0471_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6271_  (.A(\u_cpu.ALU.u_wallace._0470_ ),
    .B(\u_cpu.ALU.u_wallace._0471_ ),
    .C(\u_cpu.ALU.u_wallace._2604_ ),
    .D(\u_cpu.ALU.u_wallace._4783_ ),
    .Y(\u_cpu.ALU.u_wallace._0472_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6272_  (.A1_N(\u_cpu.ALU.u_wallace._0470_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0471_ ),
    .B1(\u_cpu.ALU.u_wallace._4471_ ),
    .B2(\u_cpu.ALU.u_wallace._4573_ ),
    .Y(\u_cpu.ALU.u_wallace._0473_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6273_  (.A1(\u_cpu.ALU.u_wallace._0316_ ),
    .A2(\u_cpu.ALU.u_wallace._0469_ ),
    .B1(\u_cpu.ALU.u_wallace._0472_ ),
    .C1(\u_cpu.ALU.u_wallace._0473_ ),
    .Y(\u_cpu.ALU.u_wallace._0474_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6274_  (.A(\u_cpu.ALU.u_wallace._4900_ ),
    .X(\u_cpu.ALU.u_wallace._0475_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._6275_  (.A1(\u_cpu.ALU.u_wallace._0322_ ),
    .A2(\u_cpu.ALU.u_wallace._0475_ ),
    .A3(\u_cpu.ALU.u_wallace._0578_ ),
    .B1(\u_cpu.ALU.u_wallace._0316_ ),
    .X(\u_cpu.ALU.u_wallace._0476_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6276_  (.A1(\u_cpu.ALU.u_wallace._0472_ ),
    .A2(\u_cpu.ALU.u_wallace._0473_ ),
    .B1(\u_cpu.ALU.u_wallace._0476_ ),
    .X(\u_cpu.ALU.u_wallace._0477_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._6277_  (.A_N(\u_cpu.ALU.u_wallace._0467_ ),
    .B(\u_cpu.ALU.u_wallace._0474_ ),
    .C(\u_cpu.ALU.u_wallace._0477_ ),
    .Y(\u_cpu.ALU.u_wallace._0478_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6278_  (.A1(\u_cpu.ALU.u_wallace._0316_ ),
    .A2(\u_cpu.ALU.u_wallace._0469_ ),
    .B1(\u_cpu.ALU.u_wallace._0472_ ),
    .C1(\u_cpu.ALU.u_wallace._0473_ ),
    .X(\u_cpu.ALU.u_wallace._0480_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6279_  (.A1(\u_cpu.ALU.u_wallace._0472_ ),
    .A2(\u_cpu.ALU.u_wallace._0473_ ),
    .B1(\u_cpu.ALU.u_wallace._0476_ ),
    .Y(\u_cpu.ALU.u_wallace._0481_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6280_  (.A1(\u_cpu.ALU.u_wallace._0480_ ),
    .A2(\u_cpu.ALU.u_wallace._0481_ ),
    .B1(\u_cpu.ALU.u_wallace._0467_ ),
    .Y(\u_cpu.ALU.u_wallace._0482_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6281_  (.A(\u_cpu.ALU.u_wallace._0466_ ),
    .B(\u_cpu.ALU.u_wallace._0478_ ),
    .C(\u_cpu.ALU.u_wallace._0482_ ),
    .Y(\u_cpu.ALU.u_wallace._0483_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6282_  (.A1(\u_cpu.ALU.u_wallace._0456_ ),
    .A2(\u_cpu.ALU.u_wallace._0462_ ),
    .B1(\u_cpu.ALU.u_wallace._0464_ ),
    .X(\u_cpu.ALU.u_wallace._0484_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._6283_  (.A(\u_cpu.ALU.u_wallace._0467_ ),
    .B(\u_cpu.ALU.u_wallace._0480_ ),
    .C(\u_cpu.ALU.u_wallace._0481_ ),
    .Y(\u_cpu.ALU.u_wallace._0485_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._6284_  (.A1(\u_cpu.ALU.u_wallace._0307_ ),
    .A2(\u_cpu.ALU.u_wallace._0292_ ),
    .B1(\u_cpu.ALU.u_wallace._0480_ ),
    .B2(\u_cpu.ALU.u_wallace._0481_ ),
    .C1(\u_cpu.ALU.u_wallace._0294_ ),
    .X(\u_cpu.ALU.u_wallace._0486_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6285_  (.A1_N(\u_cpu.ALU.u_wallace._0466_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0484_ ),
    .B1(\u_cpu.ALU.u_wallace._0485_ ),
    .B2(\u_cpu.ALU.u_wallace._0486_ ),
    .Y(\u_cpu.ALU.u_wallace._0487_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6286_  (.A1(\u_cpu.ALU.u_wallace._0347_ ),
    .A2(\u_cpu.ALU.u_wallace._0301_ ),
    .B1(\u_cpu.ALU.u_wallace._0303_ ),
    .C1(\u_cpu.ALU.u_wallace._0343_ ),
    .Y(\u_cpu.ALU.u_wallace._0488_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.ALU.u_wallace._6287_  (.A1(\u_cpu.ALU.u_wallace._0342_ ),
    .A2(\u_cpu.ALU.u_wallace._0340_ ),
    .A3(\u_cpu.ALU.u_wallace._0341_ ),
    .B1(\u_cpu.ALU.u_wallace._0488_ ),
    .Y(\u_cpu.ALU.u_wallace._0489_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6288_  (.A1(\u_cpu.ALU.u_wallace._0465_ ),
    .A2(\u_cpu.ALU.u_wallace._0483_ ),
    .B1(\u_cpu.ALU.u_wallace._0487_ ),
    .C1(\u_cpu.ALU.u_wallace._0489_ ),
    .X(\u_cpu.ALU.u_wallace._0491_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6289_  (.A(\u_cpu.ALU.u_wallace._0466_ ),
    .B(\u_cpu.ALU.u_wallace._0484_ ),
    .C(\u_cpu.ALU.u_wallace._0478_ ),
    .D(\u_cpu.ALU.u_wallace._0482_ ),
    .Y(\u_cpu.ALU.u_wallace._0492_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6290_  (.A1(\u_cpu.ALU.u_wallace._0487_ ),
    .A2(\u_cpu.ALU.u_wallace._0492_ ),
    .B1(\u_cpu.ALU.u_wallace._0489_ ),
    .Y(\u_cpu.ALU.u_wallace._0493_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._6291_  (.A1(\u_cpu.ALU.u_wallace._0346_ ),
    .A2(\u_cpu.ALU.u_wallace._0345_ ),
    .B1_N(\u_cpu.ALU.u_wallace._0302_ ),
    .Y(\u_cpu.ALU.u_wallace._0494_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6292_  (.A1(\u_cpu.ALU.u_wallace._1979_ ),
    .A2(\u_cpu.ALU.u_wallace._0364_ ),
    .B1(\u_cpu.ALU.u_wallace._0365_ ),
    .B2(\u_cpu.ALU.u_wallace._2922_ ),
    .X(\u_cpu.ALU.u_wallace._0495_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6293_  (.A(\u_cpu.ALU.u_wallace._4529_ ),
    .B(\u_cpu.ALU.u_wallace._1180_ ),
    .C(\u_cpu.ALU.u_wallace._0028_ ),
    .D(\u_cpu.ALU.u_wallace._0029_ ),
    .Y(\u_cpu.ALU.u_wallace._0496_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6294_  (.A(\u_cpu.ALU.u_wallace._1421_ ),
    .B(\u_cpu.ALU.u_wallace._0033_ ),
    .Y(\u_cpu.ALU.u_wallace._0497_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6295_  (.A1(\u_cpu.ALU.u_wallace._0495_ ),
    .A2(\u_cpu.ALU.u_wallace._0496_ ),
    .B1(\u_cpu.ALU.u_wallace._0497_ ),
    .X(\u_cpu.ALU.u_wallace._0498_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6296_  (.A1(\u_cpu.ALU.u_wallace._0610_ ),
    .A2(\u_cpu.ALU.u_wallace._0037_ ),
    .B1(\u_cpu.ALU.u_wallace._0495_ ),
    .C1(\u_cpu.ALU.u_wallace._0496_ ),
    .Y(\u_cpu.ALU.u_wallace._0499_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6297_  (.A(\u_cpu.ALU.u_wallace._0498_ ),
    .B(\u_cpu.ALU.u_wallace._0499_ ),
    .Y(\u_cpu.ALU.u_wallace._0500_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6298_  (.A(\u_cpu.ALU.u_wallace._3777_ ),
    .B(\u_cpu.ALU.u_wallace._0041_ ),
    .Y(\u_cpu.ALU.u_wallace._0502_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._6299_  (.A1(\u_cpu.ALU.u_wallace._4660_ ),
    .A2(\u_cpu.ALU.u_wallace._3821_ ),
    .A3(\u_cpu.ALU.u_wallace._4018_ ),
    .A4(\u_cpu.ALU.u_wallace._4302_ ),
    .B1(\u_cpu.ALU.u_wallace._0502_ ),
    .X(\u_cpu.ALU.u_wallace._0503_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6300_  (.A1(\u_cpu.ALU.u_wallace._4561_ ),
    .A2(\u_cpu.ALU.u_wallace._4847_ ),
    .B1(\u_cpu.ALU.u_wallace._4848_ ),
    .B2(\u_cpu.ALU.u_wallace._4447_ ),
    .Y(\u_cpu.ALU.u_wallace._0504_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6301_  (.A1(\u_cpu.ALU.u_wallace._0356_ ),
    .A2(\u_cpu.ALU.u_wallace._0354_ ),
    .B1(\u_cpu.ALU.u_wallace._0358_ ),
    .Y(\u_cpu.ALU.u_wallace._0505_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6302_  (.A(\u_cpu.ALU.u_wallace._4561_ ),
    .B(\u_cpu.ALU.u_wallace._4447_ ),
    .C(\u_cpu.ALU.u_wallace._4847_ ),
    .D(\u_cpu.ALU.u_wallace._0045_ ),
    .X(\u_cpu.ALU.u_wallace._0506_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6303_  (.A1(\u_cpu.ALU.u_wallace._0504_ ),
    .A2(\u_cpu.ALU.u_wallace._0506_ ),
    .B1(\u_cpu.ALU.u_wallace._0502_ ),
    .Y(\u_cpu.ALU.u_wallace._0507_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6304_  (.A1(\u_cpu.ALU.u_wallace._0503_ ),
    .A2(\u_cpu.ALU.u_wallace._0504_ ),
    .B1(\u_cpu.ALU.u_wallace._0505_ ),
    .C1(\u_cpu.ALU.u_wallace._0507_ ),
    .Y(\u_cpu.ALU.u_wallace._0508_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6305_  (.A(\u_cpu.ALU.u_wallace._4660_ ),
    .B(\u_cpu.ALU.u_wallace._2725_ ),
    .C(\u_cpu.ALU.u_wallace._4018_ ),
    .D(\u_cpu.ALU.u_wallace._4302_ ),
    .Y(\u_cpu.ALU.u_wallace._0509_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._6306_  (.A_N(\u_cpu.ALU.u_wallace._0504_ ),
    .B(\u_cpu.ALU.u_wallace._0509_ ),
    .C(\u_cpu.ALU.u_wallace._0198_ ),
    .D(\u_cpu.ALU.u_wallace._4610_ ),
    .Y(\u_cpu.ALU.u_wallace._0510_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6307_  (.A1(\u_cpu.ALU.u_wallace._0510_ ),
    .A2(\u_cpu.ALU.u_wallace._0507_ ),
    .B1(\u_cpu.ALU.u_wallace._0505_ ),
    .X(\u_cpu.ALU.u_wallace._0511_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6308_  (.A(\u_cpu.ALU.u_wallace._0500_ ),
    .B(\u_cpu.ALU.u_wallace._0508_ ),
    .C(\u_cpu.ALU.u_wallace._0511_ ),
    .Y(\u_cpu.ALU.u_wallace._0513_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6309_  (.A1(\u_cpu.ALU.u_wallace._0503_ ),
    .A2(\u_cpu.ALU.u_wallace._0504_ ),
    .B1(\u_cpu.ALU.u_wallace._0505_ ),
    .C1(\u_cpu.ALU.u_wallace._0507_ ),
    .X(\u_cpu.ALU.u_wallace._0514_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6310_  (.A1(\u_cpu.ALU.u_wallace._0510_ ),
    .A2(\u_cpu.ALU.u_wallace._0507_ ),
    .B1(\u_cpu.ALU.u_wallace._0505_ ),
    .Y(\u_cpu.ALU.u_wallace._0515_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._6311_  (.A1(\u_cpu.ALU.u_wallace._0514_ ),
    .A2(\u_cpu.ALU.u_wallace._0515_ ),
    .B1_N(\u_cpu.ALU.u_wallace._0500_ ),
    .Y(\u_cpu.ALU.u_wallace._0516_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6312_  (.A1(\u_cpu.ALU.u_wallace._0301_ ),
    .A2(\u_cpu.ALU.u_wallace._0494_ ),
    .B1(\u_cpu.ALU.u_wallace._0513_ ),
    .C1(\u_cpu.ALU.u_wallace._0516_ ),
    .X(\u_cpu.ALU.u_wallace._0517_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6313_  (.A1(\u_cpu.ALU.u_wallace._0302_ ),
    .A2(\u_cpu.ALU.u_wallace._0306_ ),
    .B1(\u_cpu.ALU.u_wallace._0301_ ),
    .Y(\u_cpu.ALU.u_wallace._0518_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6314_  (.A1(\u_cpu.ALU.u_wallace._0514_ ),
    .A2(\u_cpu.ALU.u_wallace._0515_ ),
    .B1(\u_cpu.ALU.u_wallace._0500_ ),
    .Y(\u_cpu.ALU.u_wallace._0519_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._6315_  (.A_N(\u_cpu.ALU.u_wallace._0500_ ),
    .B(\u_cpu.ALU.u_wallace._0508_ ),
    .C(\u_cpu.ALU.u_wallace._0511_ ),
    .Y(\u_cpu.ALU.u_wallace._0520_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._6316_  (.A1(\u_cpu.ALU.u_wallace._0368_ ),
    .A2(\u_cpu.ALU.u_wallace._0369_ ),
    .A3(\u_cpu.ALU.u_wallace._0376_ ),
    .B1(\u_cpu.ALU.u_wallace._0373_ ),
    .X(\u_cpu.ALU.u_wallace._0521_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._6317_  (.A1(\u_cpu.ALU.u_wallace._0518_ ),
    .A2(\u_cpu.ALU.u_wallace._0519_ ),
    .A3(\u_cpu.ALU.u_wallace._0520_ ),
    .B1(\u_cpu.ALU.u_wallace._0521_ ),
    .X(\u_cpu.ALU.u_wallace._0522_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6318_  (.A(\u_cpu.ALU.u_wallace._0518_ ),
    .B(\u_cpu.ALU.u_wallace._0519_ ),
    .C(\u_cpu.ALU.u_wallace._0520_ ),
    .Y(\u_cpu.ALU.u_wallace._0524_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6319_  (.A1(\u_cpu.ALU.u_wallace._0301_ ),
    .A2(\u_cpu.ALU.u_wallace._0494_ ),
    .B1(\u_cpu.ALU.u_wallace._0513_ ),
    .C1(\u_cpu.ALU.u_wallace._0516_ ),
    .Y(\u_cpu.ALU.u_wallace._0525_ ));
 sky130_fd_sc_hd__a21bo_2 \u_cpu.ALU.u_wallace._6320_  (.A1(\u_cpu.ALU.u_wallace._0524_ ),
    .A2(\u_cpu.ALU.u_wallace._0525_ ),
    .B1_N(\u_cpu.ALU.u_wallace._0521_ ),
    .X(\u_cpu.ALU.u_wallace._0526_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._6321_  (.A1(\u_cpu.ALU.u_wallace._0517_ ),
    .A2(\u_cpu.ALU.u_wallace._0522_ ),
    .B1(\u_cpu.ALU.u_wallace._0526_ ),
    .X(\u_cpu.ALU.u_wallace._0527_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6322_  (.A1(\u_cpu.ALU.u_wallace._0491_ ),
    .A2(\u_cpu.ALU.u_wallace._0493_ ),
    .B1(\u_cpu.ALU.u_wallace._0527_ ),
    .Y(\u_cpu.ALU.u_wallace._0528_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6323_  (.A1(\u_cpu.ALU.u_wallace._0517_ ),
    .A2(\u_cpu.ALU.u_wallace._0522_ ),
    .B1(\u_cpu.ALU.u_wallace._0526_ ),
    .Y(\u_cpu.ALU.u_wallace._0529_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6324_  (.A1(\u_cpu.ALU.u_wallace._0465_ ),
    .A2(\u_cpu.ALU.u_wallace._0483_ ),
    .B1(\u_cpu.ALU.u_wallace._0487_ ),
    .C1(\u_cpu.ALU.u_wallace._0489_ ),
    .Y(\u_cpu.ALU.u_wallace._0530_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6325_  (.A1(\u_cpu.ALU.u_wallace._0487_ ),
    .A2(\u_cpu.ALU.u_wallace._0492_ ),
    .B1(\u_cpu.ALU.u_wallace._0489_ ),
    .X(\u_cpu.ALU.u_wallace._0531_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6326_  (.A(\u_cpu.ALU.u_wallace._0529_ ),
    .B(\u_cpu.ALU.u_wallace._0530_ ),
    .C(\u_cpu.ALU.u_wallace._0531_ ),
    .Y(\u_cpu.ALU.u_wallace._0532_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6327_  (.A1(\u_cpu.ALU.u_wallace._0192_ ),
    .A2(\u_cpu.ALU.u_wallace._0350_ ),
    .B1(\u_cpu.ALU.u_wallace._0393_ ),
    .Y(\u_cpu.ALU.u_wallace._0533_ ));
 sky130_fd_sc_hd__a32oi_2 \u_cpu.ALU.u_wallace._6328_  (.A1(\u_cpu.ALU.u_wallace._0395_ ),
    .A2(\u_cpu.ALU.u_wallace._0388_ ),
    .A3(\u_cpu.ALU.u_wallace._0397_ ),
    .B1(\u_cpu.ALU.u_wallace._0533_ ),
    .B2(\u_cpu.ALU.u_wallace._0344_ ),
    .Y(\u_cpu.ALU.u_wallace._0535_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6329_  (.A(\u_cpu.ALU.u_wallace._0528_ ),
    .B(\u_cpu.ALU.u_wallace._0532_ ),
    .C(\u_cpu.ALU.u_wallace._0535_ ),
    .Y(\u_cpu.ALU.u_wallace._0536_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6330_  (.A1(\u_cpu.ALU.u_wallace._0522_ ),
    .A2(\u_cpu.ALU.u_wallace._0517_ ),
    .B1(\u_cpu.ALU.u_wallace._0526_ ),
    .C1(\u_cpu.ALU.u_wallace._0530_ ),
    .Y(\u_cpu.ALU.u_wallace._0537_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6331_  (.A1(\u_cpu.ALU.u_wallace._0192_ ),
    .A2(\u_cpu.ALU.u_wallace._0350_ ),
    .B1(\u_cpu.ALU.u_wallace._0393_ ),
    .X(\u_cpu.ALU.u_wallace._0538_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6332_  (.A1(\u_cpu.ALU.u_wallace._0378_ ),
    .A2(\u_cpu.ALU.u_wallace._0384_ ),
    .B1(\u_cpu.ALU.u_wallace._0388_ ),
    .Y(\u_cpu.ALU.u_wallace._0539_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6333_  (.A1(\u_cpu.ALU.u_wallace._0391_ ),
    .A2(\u_cpu.ALU.u_wallace._0538_ ),
    .B1(\u_cpu.ALU.u_wallace._0352_ ),
    .B2(\u_cpu.ALU.u_wallace._0539_ ),
    .Y(\u_cpu.ALU.u_wallace._0540_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._6334_  (.A1(\u_cpu.ALU.u_wallace._0518_ ),
    .A2(\u_cpu.ALU.u_wallace._0519_ ),
    .A3(\u_cpu.ALU.u_wallace._0520_ ),
    .B1(\u_cpu.ALU.u_wallace._0521_ ),
    .Y(\u_cpu.ALU.u_wallace._0541_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6335_  (.A(\u_cpu.ALU.u_wallace._0541_ ),
    .B(\u_cpu.ALU.u_wallace._0525_ ),
    .Y(\u_cpu.ALU.u_wallace._0542_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6336_  (.A1_N(\u_cpu.ALU.u_wallace._0526_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0542_ ),
    .B1(\u_cpu.ALU.u_wallace._0491_ ),
    .B2(\u_cpu.ALU.u_wallace._0493_ ),
    .Y(\u_cpu.ALU.u_wallace._0543_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6337_  (.A1(\u_cpu.ALU.u_wallace._0537_ ),
    .A2(\u_cpu.ALU.u_wallace._0493_ ),
    .B1(\u_cpu.ALU.u_wallace._0540_ ),
    .C1(\u_cpu.ALU.u_wallace._0543_ ),
    .Y(\u_cpu.ALU.u_wallace._0544_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6338_  (.A(\u_cpu.ALU.SrcB[14] ),
    .X(\u_cpu.ALU.u_wallace._0546_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6339_  (.A(\u_cpu.ALU.SrcB[15] ),
    .X(\u_cpu.ALU.u_wallace._0547_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6340_  (.A1(\u_cpu.ALU.u_wallace._0512_ ),
    .A2(\u_cpu.ALU.u_wallace._0546_ ),
    .B1(\u_cpu.ALU.u_wallace._0547_ ),
    .B2(\u_cpu.ALU.u_wallace._0250_ ),
    .X(\u_cpu.ALU.u_wallace._0548_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6341_  (.A(\u_cpu.ALU.u_wallace._4597_ ),
    .B(\u_cpu.ALU.u_wallace._0151_ ),
    .C(\u_cpu.ALU.u_wallace._0546_ ),
    .D(\u_cpu.ALU.u_wallace._0279_ ),
    .Y(\u_cpu.ALU.u_wallace._0549_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6342_  (.A(\u_cpu.ALU.SrcB[16] ),
    .X(\u_cpu.ALU.u_wallace._0550_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6343_  (.A(\u_cpu.ALU.u_wallace._0550_ ),
    .X(\u_cpu.ALU.u_wallace._0551_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6344_  (.A(\u_cpu.ALU.u_wallace._0548_ ),
    .B(\u_cpu.ALU.u_wallace._0549_ ),
    .C(\u_cpu.ALU.u_wallace._0994_ ),
    .D(\u_cpu.ALU.u_wallace._0551_ ),
    .Y(\u_cpu.ALU.u_wallace._0552_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._6345_  (.A(\u_cpu.ALU.SrcB[16] ),
    .Y(\u_cpu.ALU.u_wallace._0553_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6346_  (.A(\u_cpu.ALU.u_wallace._0553_ ),
    .X(\u_cpu.ALU.u_wallace._0554_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6347_  (.A(\u_cpu.ALU.u_wallace._1410_ ),
    .B(\u_cpu.ALU.u_wallace._0546_ ),
    .Y(\u_cpu.ALU.u_wallace._0555_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6348_  (.A(\u_cpu.ALU.u_wallace._0555_ ),
    .B(\u_cpu.ALU.u_wallace._0279_ ),
    .C(\u_cpu.ALU.u_wallace._1454_ ),
    .Y(\u_cpu.ALU.u_wallace._0557_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6349_  (.A(\u_cpu.ALU.u_wallace._0731_ ),
    .B(\u_cpu.ALU.u_wallace._0279_ ),
    .Y(\u_cpu.ALU.u_wallace._0558_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6350_  (.A(\u_cpu.ALU.u_wallace._0558_ ),
    .B(\u_cpu.ALU.u_wallace._0121_ ),
    .C(\u_cpu.ALU.u_wallace._0359_ ),
    .Y(\u_cpu.ALU.u_wallace._0559_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6351_  (.A1(\u_cpu.ALU.u_wallace._0032_ ),
    .A2(\u_cpu.ALU.u_wallace._0554_ ),
    .B1(\u_cpu.ALU.u_wallace._0557_ ),
    .C1(\u_cpu.ALU.u_wallace._0559_ ),
    .Y(\u_cpu.ALU.u_wallace._0560_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6352_  (.A(\u_cpu.ALU.u_wallace._0359_ ),
    .B(\u_cpu.ALU.u_wallace._0363_ ),
    .Y(\u_cpu.ALU.u_wallace._0561_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6353_  (.A1(\u_cpu.ALU.u_wallace._2933_ ),
    .A2(\u_cpu.ALU.u_wallace._4840_ ),
    .B1(\u_cpu.ALU.u_wallace._4842_ ),
    .B2(\u_cpu.ALU.u_wallace._4527_ ),
    .Y(\u_cpu.ALU.u_wallace._0562_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6354_  (.A1(\u_cpu.ALU.u_wallace._0561_ ),
    .A2(\u_cpu.ALU.u_wallace._0562_ ),
    .B1(\u_cpu.ALU.u_wallace._0367_ ),
    .Y(\u_cpu.ALU.u_wallace._0563_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6355_  (.A1(\u_cpu.ALU.u_wallace._0552_ ),
    .A2(\u_cpu.ALU.u_wallace._0560_ ),
    .B1(\u_cpu.ALU.u_wallace._0563_ ),
    .Y(\u_cpu.ALU.u_wallace._0564_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6356_  (.A(\u_cpu.ALU.u_wallace._0563_ ),
    .B(\u_cpu.ALU.u_wallace._0552_ ),
    .C(\u_cpu.ALU.u_wallace._0560_ ),
    .X(\u_cpu.ALU.u_wallace._0565_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._6357_  (.A1(\u_cpu.ALU.u_wallace._0283_ ),
    .A2(\u_cpu.ALU.u_wallace._0287_ ),
    .B1(\u_cpu.ALU.u_wallace._0564_ ),
    .C1(\u_cpu.ALU.u_wallace._0565_ ),
    .X(\u_cpu.ALU.u_wallace._0566_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6358_  (.A1(\u_cpu.ALU.u_wallace._0564_ ),
    .A2(\u_cpu.ALU.u_wallace._0565_ ),
    .B1(\u_cpu.ALU.u_wallace._0283_ ),
    .C1(\u_cpu.ALU.u_wallace._0287_ ),
    .Y(\u_cpu.ALU.u_wallace._0568_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6359_  (.A(\u_cpu.ALU.u_wallace._0566_ ),
    .B(\u_cpu.ALU.u_wallace._0568_ ),
    .Y(\u_cpu.ALU.u_wallace._0569_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6360_  (.A1(\u_cpu.ALU.u_wallace._0386_ ),
    .A2(\u_cpu.ALU.u_wallace._0384_ ),
    .B1(\u_cpu.ALU.u_wallace._0569_ ),
    .Y(\u_cpu.ALU.u_wallace._0570_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6361_  (.A1(\u_cpu.ALU.u_wallace._0374_ ),
    .A2(\u_cpu.ALU.u_wallace._0377_ ),
    .B1(\u_cpu.ALU.u_wallace._0353_ ),
    .Y(\u_cpu.ALU.u_wallace._0571_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6362_  (.A1(\u_cpu.ALU.u_wallace._0383_ ),
    .A2(\u_cpu.ALU.u_wallace._0571_ ),
    .B1(\u_cpu.ALU.u_wallace._0386_ ),
    .C1(\u_cpu.ALU.u_wallace._0569_ ),
    .Y(\u_cpu.ALU.u_wallace._0572_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6363_  (.A(\u_cpu.ALU.u_wallace._0286_ ),
    .B(\u_cpu.ALU.u_wallace._0287_ ),
    .C(\u_cpu.ALU.u_wallace._0572_ ),
    .D(\u_cpu.ALU.u_wallace._0123_ ),
    .Y(\u_cpu.ALU.u_wallace._0573_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._6364_  (.A(\u_cpu.ALU.u_wallace._0119_ ),
    .Y(\u_cpu.ALU.u_wallace._0574_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6365_  (.A1(\u_cpu.ALU.u_wallace._0383_ ),
    .A2(\u_cpu.ALU.u_wallace._0571_ ),
    .B1(\u_cpu.ALU.u_wallace._0386_ ),
    .C1(\u_cpu.ALU.u_wallace._0569_ ),
    .X(\u_cpu.ALU.u_wallace._0575_ ));
 sky130_fd_sc_hd__o32ai_2 \u_cpu.ALU.u_wallace._6366_  (.A1(\u_cpu.ALU.u_wallace._0125_ ),
    .A2(\u_cpu.ALU.u_wallace._0288_ ),
    .A3(\u_cpu.ALU.u_wallace._0574_ ),
    .B1(\u_cpu.ALU.u_wallace._0575_ ),
    .B2(\u_cpu.ALU.u_wallace._0570_ ),
    .Y(\u_cpu.ALU.u_wallace._0576_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._6367_  (.A1(\u_cpu.ALU.u_wallace._0570_ ),
    .A2(\u_cpu.ALU.u_wallace._0573_ ),
    .B1(\u_cpu.ALU.u_wallace._0576_ ),
    .X(\u_cpu.ALU.u_wallace._0577_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6368_  (.A1(\u_cpu.ALU.u_wallace._0536_ ),
    .A2(\u_cpu.ALU.u_wallace._0544_ ),
    .B1(\u_cpu.ALU.u_wallace._0577_ ),
    .X(\u_cpu.ALU.u_wallace._0579_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._6369_  (.A1(\u_cpu.ALU.u_wallace._0570_ ),
    .A2(\u_cpu.ALU.u_wallace._0573_ ),
    .B1(\u_cpu.ALU.u_wallace._0576_ ),
    .C1(\u_cpu.ALU.u_wallace._0536_ ),
    .D1(\u_cpu.ALU.u_wallace._0544_ ),
    .Y(\u_cpu.ALU.u_wallace._0580_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6370_  (.A(\u_cpu.ALU.u_wallace._0437_ ),
    .B(\u_cpu.ALU.u_wallace._0579_ ),
    .C(\u_cpu.ALU.u_wallace._0580_ ),
    .Y(\u_cpu.ALU.u_wallace._0581_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6371_  (.A1(\u_cpu.ALU.u_wallace._0536_ ),
    .A2(\u_cpu.ALU.u_wallace._0544_ ),
    .B1(\u_cpu.ALU.u_wallace._0577_ ),
    .Y(\u_cpu.ALU.u_wallace._0582_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._6372_  (.A1(\u_cpu.ALU.u_wallace._0570_ ),
    .A2(\u_cpu.ALU.u_wallace._0573_ ),
    .B1(\u_cpu.ALU.u_wallace._0576_ ),
    .C1(\u_cpu.ALU.u_wallace._0536_ ),
    .D1(\u_cpu.ALU.u_wallace._0544_ ),
    .X(\u_cpu.ALU.u_wallace._0583_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._6373_  (.A1(\u_cpu.ALU.u_wallace._0582_ ),
    .A2(\u_cpu.ALU.u_wallace._0583_ ),
    .B1_N(\u_cpu.ALU.u_wallace._0437_ ),
    .Y(\u_cpu.ALU.u_wallace._0584_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._6374_  (.A(\u_cpu.ALU.u_wallace._0277_ ),
    .Y(\u_cpu.ALU.u_wallace._0585_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6375_  (.A1_N(\u_cpu.ALU.u_wallace._0581_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0584_ ),
    .B1(\u_cpu.ALU.u_wallace._0585_ ),
    .B2(\u_cpu.ALU.u_wallace._0289_ ),
    .Y(\u_cpu.ALU.u_wallace._0586_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6376_  (.A1(\u_cpu.ALU.u_wallace._0159_ ),
    .A2(\u_cpu.ALU.u_wallace._0231_ ),
    .B1(\u_cpu.ALU.u_wallace._0289_ ),
    .Y(\u_cpu.ALU.u_wallace._0587_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6377_  (.A(\u_cpu.ALU.u_wallace._0584_ ),
    .B(\u_cpu.ALU.u_wallace._0587_ ),
    .C(\u_cpu.ALU.u_wallace._0581_ ),
    .Y(\u_cpu.ALU.u_wallace._0588_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6378_  (.A(\u_cpu.ALU.u_wallace._0416_ ),
    .B(\u_cpu.ALU.u_wallace._0417_ ),
    .C(\u_cpu.ALU.u_wallace._0418_ ),
    .X(\u_cpu.ALU.u_wallace._0590_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU.u_wallace._6379_  (.A1(\u_cpu.ALU.u_wallace._0415_ ),
    .A2(\u_cpu.ALU.u_wallace._0128_ ),
    .B1(\u_cpu.ALU.u_wallace._0586_ ),
    .B2(\u_cpu.ALU.u_wallace._0588_ ),
    .C1(\u_cpu.ALU.u_wallace._0590_ ),
    .X(\u_cpu.ALU.u_wallace._0591_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._6380_  (.A1(\u_cpu.ALU.u_wallace._0416_ ),
    .A2(\u_cpu.ALU.u_wallace._0417_ ),
    .A3(\u_cpu.ALU.u_wallace._0418_ ),
    .B1(\u_cpu.ALU.u_wallace._0415_ ),
    .B2(\u_cpu.ALU.u_wallace._0128_ ),
    .X(\u_cpu.ALU.u_wallace._0592_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6381_  (.A(\u_cpu.ALU.u_wallace._0592_ ),
    .B(\u_cpu.ALU.u_wallace._0588_ ),
    .C(\u_cpu.ALU.u_wallace._0586_ ),
    .Y(\u_cpu.ALU.u_wallace._0593_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6382_  (.A(\u_cpu.ALU.u_wallace._0591_ ),
    .B(\u_cpu.ALU.u_wallace._0593_ ),
    .Y(\u_cpu.ALU.u_wallace._0594_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._6383_  (.A(\u_cpu.ALU.u_wallace._0436_ ),
    .B(\u_cpu.ALU.u_wallace._0594_ ),
    .X(\u_cpu.ALU.u_wallace._0595_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._6384_  (.A1(\u_cpu.ALU.u_wallace._0100_ ),
    .A2(\u_cpu.ALU.u_wallace._0256_ ),
    .A3(\u_cpu.ALU.u_wallace._0263_ ),
    .B1(\u_cpu.ALU.u_wallace._0428_ ),
    .B2(\u_cpu.ALU.u_wallace._0430_ ),
    .X(\u_cpu.ALU.u_wallace._0596_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6385_  (.A(\u_cpu.ALU.u_wallace._0275_ ),
    .B(\u_cpu.ALU.u_wallace._0428_ ),
    .Y(\u_cpu.ALU.u_wallace._0597_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6386_  (.A(\u_cpu.ALU.u_wallace._0267_ ),
    .B(\u_cpu.ALU.u_wallace._0269_ ),
    .C(\u_cpu.ALU.u_wallace._0596_ ),
    .D(\u_cpu.ALU.u_wallace._0597_ ),
    .Y(\u_cpu.ALU.u_wallace._0598_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6387_  (.A1(\u_cpu.ALU.u_wallace._0269_ ),
    .A2(\u_cpu.ALU.u_wallace._0597_ ),
    .B1(\u_cpu.ALU.u_wallace._0431_ ),
    .X(\u_cpu.ALU.u_wallace._0599_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6388_  (.A1(\u_cpu.ALU.u_wallace._0274_ ),
    .A2(\u_cpu.ALU.u_wallace._0598_ ),
    .B1(\u_cpu.ALU.u_wallace._0599_ ),
    .Y(\u_cpu.ALU.u_wallace._0601_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._6389_  (.A(\u_cpu.ALU.u_wallace._0595_ ),
    .B(\u_cpu.ALU.u_wallace._0601_ ),
    .X(\u_cpu.ALU.Product_Wallace[16] ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6390_  (.A(\u_cpu.ALU.u_wallace._0592_ ),
    .B(\u_cpu.ALU.u_wallace._0588_ ),
    .C(\u_cpu.ALU.u_wallace._0586_ ),
    .X(\u_cpu.ALU.u_wallace._0602_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6391_  (.A1(\u_cpu.ALU.u_wallace._0588_ ),
    .A2(\u_cpu.ALU.u_wallace._0586_ ),
    .B1(\u_cpu.ALU.u_wallace._0592_ ),
    .Y(\u_cpu.ALU.u_wallace._0603_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6392_  (.A1(\u_cpu.ALU.u_wallace._0537_ ),
    .A2(\u_cpu.ALU.u_wallace._0493_ ),
    .B1(\u_cpu.ALU.u_wallace._0540_ ),
    .C1(\u_cpu.ALU.u_wallace._0543_ ),
    .X(\u_cpu.ALU.u_wallace._0604_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6393_  (.A1(\u_cpu.ALU.u_wallace._0570_ ),
    .A2(\u_cpu.ALU.u_wallace._0573_ ),
    .B1(\u_cpu.ALU.u_wallace._0576_ ),
    .C1(\u_cpu.ALU.u_wallace._0536_ ),
    .X(\u_cpu.ALU.u_wallace._0605_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6394_  (.A(\u_cpu.ALU.u_wallace._2045_ ),
    .B(\u_cpu.ALU.u_wallace._2056_ ),
    .C(\u_cpu.ALU.u_wallace._4653_ ),
    .D(\u_cpu.ALU.u_wallace._4787_ ),
    .X(\u_cpu.ALU.u_wallace._0606_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6395_  (.A(\u_cpu.ALU.u_wallace._4567_ ),
    .X(\u_cpu.ALU.u_wallace._0607_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6396_  (.A(\u_cpu.ALU.u_wallace._0470_ ),
    .B(\u_cpu.ALU.u_wallace._0607_ ),
    .C(\u_cpu.ALU.u_wallace._0015_ ),
    .X(\u_cpu.ALU.u_wallace._0608_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._6397_  (.A(\u_cpu.ALU.u_wallace._0438_ ),
    .B(\u_cpu.ALU.u_wallace._0440_ ),
    .Y(\u_cpu.ALU.u_wallace._0609_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6398_  (.A1(\u_cpu.ALU.u_wallace._2078_ ),
    .A2(\u_cpu.ALU.u_wallace._4785_ ),
    .B1(\u_cpu.ALU.u_wallace._4907_ ),
    .B2(\u_cpu.ALU.u_wallace._4467_ ),
    .X(\u_cpu.ALU.u_wallace._0611_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6399_  (.A(\u_cpu.ALU.u_wallace._1530_ ),
    .B(\u_cpu.ALU.u_wallace._2056_ ),
    .C(\u_cpu.ALU.u_wallace._4787_ ),
    .D(\u_cpu.ALU.u_wallace._4921_ ),
    .Y(\u_cpu.ALU.u_wallace._0612_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6400_  (.A(\u_cpu.ALU.u_wallace._0611_ ),
    .B(\u_cpu.ALU.u_wallace._0612_ ),
    .C(\u_cpu.ALU.u_wallace._2626_ ),
    .D(\u_cpu.ALU.u_wallace._4643_ ),
    .Y(\u_cpu.ALU.u_wallace._0613_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6401_  (.A1(\u_cpu.ALU.u_wallace._2056_ ),
    .A2(\u_cpu.ALU.u_wallace._4787_ ),
    .B1(\u_cpu.ALU.u_wallace._0188_ ),
    .B2(\u_cpu.ALU.u_wallace._1530_ ),
    .Y(\u_cpu.ALU.u_wallace._0614_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6402_  (.A(\u_cpu.ALU.u_wallace._4467_ ),
    .B(\u_cpu.ALU.u_wallace._1497_ ),
    .C(\u_cpu.ALU.u_wallace._4785_ ),
    .D(\u_cpu.ALU.u_wallace._4907_ ),
    .X(\u_cpu.ALU.u_wallace._0615_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6403_  (.A1(\u_cpu.ALU.u_wallace._4471_ ),
    .A2(\u_cpu.ALU.u_wallace._4904_ ),
    .B1(\u_cpu.ALU.u_wallace._0614_ ),
    .B2(\u_cpu.ALU.u_wallace._0615_ ),
    .Y(\u_cpu.ALU.u_wallace._0616_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6404_  (.A1(\u_cpu.ALU.u_wallace._0459_ ),
    .A2(\u_cpu.ALU.u_wallace._0609_ ),
    .B1(\u_cpu.ALU.u_wallace._0613_ ),
    .C1(\u_cpu.ALU.u_wallace._0616_ ),
    .Y(\u_cpu.ALU.u_wallace._0617_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6405_  (.A1(\u_cpu.ALU.u_wallace._0438_ ),
    .A2(\u_cpu.ALU.u_wallace._0440_ ),
    .B1(\u_cpu.ALU.u_wallace._0454_ ),
    .Y(\u_cpu.ALU.u_wallace._0618_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6406_  (.A1(\u_cpu.ALU.u_wallace._0613_ ),
    .A2(\u_cpu.ALU.u_wallace._0616_ ),
    .B1(\u_cpu.ALU.u_wallace._0618_ ),
    .X(\u_cpu.ALU.u_wallace._0619_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._6407_  (.A1_N(\u_cpu.ALU.u_wallace._0606_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0608_ ),
    .B1(\u_cpu.ALU.u_wallace._0617_ ),
    .B2(\u_cpu.ALU.u_wallace._0619_ ),
    .Y(\u_cpu.ALU.u_wallace._0620_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._6408_  (.A1(\u_cpu.ALU.u_wallace._0459_ ),
    .A2(\u_cpu.ALU.u_wallace._0609_ ),
    .B1(\u_cpu.ALU.u_wallace._0616_ ),
    .X(\u_cpu.ALU.u_wallace._0622_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._6409_  (.A1(\u_cpu.ALU.u_wallace._0470_ ),
    .A2(\u_cpu.ALU.u_wallace._0607_ ),
    .A3(\u_cpu.ALU.u_wallace._3481_ ),
    .B1(\u_cpu.ALU.u_wallace._0606_ ),
    .X(\u_cpu.ALU.u_wallace._0623_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6410_  (.A1(\u_cpu.ALU.u_wallace._0613_ ),
    .A2(\u_cpu.ALU.u_wallace._0616_ ),
    .B1(\u_cpu.ALU.u_wallace._0618_ ),
    .Y(\u_cpu.ALU.u_wallace._0624_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU.u_wallace._6411_  (.A1(\u_cpu.ALU.u_wallace._0622_ ),
    .A2(\u_cpu.ALU.u_wallace._0613_ ),
    .B1(\u_cpu.ALU.u_wallace._0623_ ),
    .C1(\u_cpu.ALU.u_wallace._0624_ ),
    .Y(\u_cpu.ALU.u_wallace._0625_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6412_  (.A(\u_cpu.ALU.SrcB[17] ),
    .X(\u_cpu.ALU.u_wallace._0626_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6413_  (.A1(\u_cpu.ALU.u_wallace._1815_ ),
    .A2(\u_cpu.ALU.u_wallace._4646_ ),
    .B1(\u_cpu.ALU.u_wallace._0626_ ),
    .B2(\u_cpu.ALU.u_wallace._0010_ ),
    .Y(\u_cpu.ALU.u_wallace._0627_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6414_  (.A(\u_cpu.ALU.SrcB[17] ),
    .X(\u_cpu.ALU.u_wallace._0628_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6415_  (.A(\u_cpu.ALU.u_wallace._0628_ ),
    .X(\u_cpu.ALU.u_wallace._0629_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6416_  (.A(\u_cpu.ALU.SrcA[17] ),
    .X(\u_cpu.ALU.u_wallace._0630_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6417_  (.A(\u_cpu.ALU.u_wallace._0862_ ),
    .B(\u_cpu.ALU.u_wallace._0630_ ),
    .Y(\u_cpu.ALU.u_wallace._0631_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._6418_  (.A1(\u_cpu.ALU.u_wallace._0010_ ),
    .A2(\u_cpu.ALU.u_wallace._4431_ ),
    .A3(\u_cpu.ALU.u_wallace._4653_ ),
    .A4(\u_cpu.ALU.u_wallace._0629_ ),
    .B1(\u_cpu.ALU.u_wallace._0631_ ),
    .X(\u_cpu.ALU.u_wallace._0633_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6419_  (.A(\u_cpu.ALU.u_wallace._4912_ ),
    .X(\u_cpu.ALU.u_wallace._0634_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._6420_  (.A(\u_cpu.ALU.u_wallace._0630_ ),
    .Y(\u_cpu.ALU.u_wallace._0635_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6421_  (.A(\u_cpu.ALU.SrcA[0] ),
    .B(\u_cpu.ALU.u_wallace._1760_ ),
    .C(\u_cpu.ALU.u_wallace._4646_ ),
    .D(\u_cpu.ALU.SrcB[17] ),
    .X(\u_cpu.ALU.u_wallace._0636_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6422_  (.A1(\u_cpu.ALU.u_wallace._0634_ ),
    .A2(\u_cpu.ALU.u_wallace._0635_ ),
    .B1(\u_cpu.ALU.u_wallace._0627_ ),
    .B2(\u_cpu.ALU.u_wallace._0636_ ),
    .Y(\u_cpu.ALU.u_wallace._0637_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6423_  (.A1(\u_cpu.ALU.u_wallace._0627_ ),
    .A2(\u_cpu.ALU.u_wallace._0633_ ),
    .B1(\u_cpu.ALU.u_wallace._0451_ ),
    .C1(\u_cpu.ALU.u_wallace._0637_ ),
    .X(\u_cpu.ALU.u_wallace._0638_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6424_  (.A(\u_cpu.ALU.SrcB[17] ),
    .X(\u_cpu.ALU.u_wallace._0639_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6425_  (.A1(\u_cpu.ALU.u_wallace._2856_ ),
    .A2(\u_cpu.ALU.u_wallace._4797_ ),
    .B1(\u_cpu.ALU.u_wallace._0639_ ),
    .B2(\u_cpu.ALU.u_wallace._0010_ ),
    .X(\u_cpu.ALU.u_wallace._0640_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6426_  (.A(\u_cpu.ALU.u_wallace._0010_ ),
    .B(\u_cpu.ALU.u_wallace._2856_ ),
    .C(\u_cpu.ALU.u_wallace._4797_ ),
    .D(\u_cpu.ALU.u_wallace._0639_ ),
    .Y(\u_cpu.ALU.u_wallace._0641_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6427_  (.A(\u_cpu.ALU.SrcA[17] ),
    .X(\u_cpu.ALU.u_wallace._0642_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6428_  (.A(\u_cpu.ALU.u_wallace._0640_ ),
    .B(\u_cpu.ALU.u_wallace._0641_ ),
    .C(\u_cpu.ALU.u_wallace._2757_ ),
    .D(\u_cpu.ALU.u_wallace._0642_ ),
    .Y(\u_cpu.ALU.u_wallace._0644_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6429_  (.A1(\u_cpu.ALU.u_wallace._0644_ ),
    .A2(\u_cpu.ALU.u_wallace._0637_ ),
    .B1(\u_cpu.ALU.u_wallace._0451_ ),
    .Y(\u_cpu.ALU.u_wallace._0645_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6430_  (.A(\u_cpu.ALU.u_wallace._0797_ ),
    .B(\u_cpu.ALU.u_wallace._0293_ ),
    .C(\u_cpu.ALU.u_wallace._0324_ ),
    .D(\u_cpu.ALU.u_wallace._0447_ ),
    .Y(\u_cpu.ALU.u_wallace._0646_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6431_  (.A(\u_cpu.ALU.u_wallace._0646_ ),
    .B(\u_cpu.ALU.u_wallace._0179_ ),
    .C(\u_cpu.ALU.u_wallace._0753_ ),
    .X(\u_cpu.ALU.u_wallace._0647_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6432_  (.A1(\u_cpu.ALU.u_wallace._0293_ ),
    .A2(\u_cpu.ALU.u_wallace._0324_ ),
    .B1(\u_cpu.ALU.u_wallace._0441_ ),
    .B2(\u_cpu.ALU.u_wallace._0797_ ),
    .X(\u_cpu.ALU.u_wallace._0648_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6433_  (.A1(\u_cpu.ALU.u_wallace._0840_ ),
    .A2(\u_cpu.ALU.u_wallace._0320_ ),
    .B1(\u_cpu.ALU.u_wallace._0648_ ),
    .B2(\u_cpu.ALU.u_wallace._0646_ ),
    .Y(\u_cpu.ALU.u_wallace._0649_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6434_  (.A1(\u_cpu.ALU.u_wallace._0647_ ),
    .A2(\u_cpu.ALU.u_wallace._0648_ ),
    .B1(\u_cpu.ALU.u_wallace._0649_ ),
    .Y(\u_cpu.ALU.u_wallace._0650_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6435_  (.A1(\u_cpu.ALU.u_wallace._0638_ ),
    .A2(\u_cpu.ALU.u_wallace._0645_ ),
    .B1(\u_cpu.ALU.u_wallace._0650_ ),
    .Y(\u_cpu.ALU.u_wallace._0651_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6436_  (.A(\u_cpu.ALU.u_wallace._0313_ ),
    .X(\u_cpu.ALU.u_wallace._0652_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6437_  (.A(\u_cpu.ALU.u_wallace._0648_ ),
    .B(\u_cpu.ALU.u_wallace._0646_ ),
    .C(\u_cpu.ALU.u_wallace._0578_ ),
    .D(\u_cpu.ALU.u_wallace._0652_ ),
    .X(\u_cpu.ALU.u_wallace._0653_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6438_  (.A1(\u_cpu.ALU.u_wallace._0627_ ),
    .A2(\u_cpu.ALU.u_wallace._0633_ ),
    .B1(\u_cpu.ALU.u_wallace._0451_ ),
    .C1(\u_cpu.ALU.u_wallace._0637_ ),
    .Y(\u_cpu.ALU.u_wallace._0655_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6439_  (.A1_N(\u_cpu.ALU.u_wallace._0644_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0637_ ),
    .B1(\u_cpu.ALU.u_wallace._0442_ ),
    .B2(\u_cpu.ALU.u_wallace._0443_ ),
    .Y(\u_cpu.ALU.u_wallace._0656_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6440_  (.A1(\u_cpu.ALU.u_wallace._0653_ ),
    .A2(\u_cpu.ALU.u_wallace._0649_ ),
    .B1(\u_cpu.ALU.u_wallace._0655_ ),
    .C1(\u_cpu.ALU.u_wallace._0656_ ),
    .Y(\u_cpu.ALU.u_wallace._0657_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._6441_  (.A1(\u_cpu.ALU.u_wallace._0333_ ),
    .A2(\u_cpu.ALU.u_wallace._0449_ ),
    .A3(\u_cpu.ALU.u_wallace._0451_ ),
    .B1(\u_cpu.ALU.u_wallace._0456_ ),
    .X(\u_cpu.ALU.u_wallace._0658_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6442_  (.A(\u_cpu.ALU.u_wallace._0651_ ),
    .B(\u_cpu.ALU.u_wallace._0657_ ),
    .C(\u_cpu.ALU.u_wallace._0658_ ),
    .Y(\u_cpu.ALU.u_wallace._0659_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6443_  (.A1(\u_cpu.ALU.u_wallace._0620_ ),
    .A2(\u_cpu.ALU.u_wallace._0625_ ),
    .B1(\u_cpu.ALU.u_wallace._0659_ ),
    .Y(\u_cpu.ALU.u_wallace._0660_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._6444_  (.A(\u_cpu.ALU.u_wallace._0333_ ),
    .B(\u_cpu.ALU.u_wallace._0449_ ),
    .C(\u_cpu.ALU.u_wallace._0451_ ),
    .Y(\u_cpu.ALU.u_wallace._0661_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._6445_  (.A1(\u_cpu.ALU.u_wallace._0439_ ),
    .A2(\u_cpu.ALU.u_wallace._0440_ ),
    .B1(\u_cpu.ALU.u_wallace._0445_ ),
    .C1(\u_cpu.ALU.u_wallace._0452_ ),
    .D1(\u_cpu.ALU.u_wallace._0455_ ),
    .X(\u_cpu.ALU.u_wallace._0662_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6446_  (.A(\u_cpu.ALU.u_wallace._0656_ ),
    .B(\u_cpu.ALU.u_wallace._0650_ ),
    .Y(\u_cpu.ALU.u_wallace._0663_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6447_  (.A1(\u_cpu.ALU.u_wallace._0653_ ),
    .A2(\u_cpu.ALU.u_wallace._0649_ ),
    .B1(\u_cpu.ALU.u_wallace._0638_ ),
    .B2(\u_cpu.ALU.u_wallace._0645_ ),
    .Y(\u_cpu.ALU.u_wallace._0664_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._6448_  (.A1(\u_cpu.ALU.u_wallace._0661_ ),
    .A2(\u_cpu.ALU.u_wallace._0662_ ),
    .B1(\u_cpu.ALU.u_wallace._0638_ ),
    .B2(\u_cpu.ALU.u_wallace._0663_ ),
    .C1(\u_cpu.ALU.u_wallace._0664_ ),
    .X(\u_cpu.ALU.u_wallace._0666_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6449_  (.A(\u_cpu.ALU.u_wallace._0464_ ),
    .B(\u_cpu.ALU.u_wallace._0456_ ),
    .C(\u_cpu.ALU.u_wallace._0462_ ),
    .X(\u_cpu.ALU.u_wallace._0667_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._6450_  (.A1(\u_cpu.ALU.u_wallace._0484_ ),
    .A2(\u_cpu.ALU.u_wallace._0478_ ),
    .A3(\u_cpu.ALU.u_wallace._0482_ ),
    .B1(\u_cpu.ALU.u_wallace._0667_ ),
    .X(\u_cpu.ALU.u_wallace._0668_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6451_  (.A1(\u_cpu.ALU.u_wallace._0606_ ),
    .A2(\u_cpu.ALU.u_wallace._0608_ ),
    .B1(\u_cpu.ALU.u_wallace._0617_ ),
    .C1(\u_cpu.ALU.u_wallace._0619_ ),
    .X(\u_cpu.ALU.u_wallace._0669_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6452_  (.A1(\u_cpu.ALU.u_wallace._0617_ ),
    .A2(\u_cpu.ALU.u_wallace._0619_ ),
    .B1(\u_cpu.ALU.u_wallace._0623_ ),
    .Y(\u_cpu.ALU.u_wallace._0670_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._6453_  (.A1(\u_cpu.ALU.u_wallace._0661_ ),
    .A2(\u_cpu.ALU.u_wallace._0662_ ),
    .B1(\u_cpu.ALU.u_wallace._0638_ ),
    .B2(\u_cpu.ALU.u_wallace._0663_ ),
    .C1(\u_cpu.ALU.u_wallace._0664_ ),
    .Y(\u_cpu.ALU.u_wallace._0671_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.ALU.u_wallace._6454_  (.A1_N(\u_cpu.ALU.u_wallace._0669_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0670_ ),
    .B1(\u_cpu.ALU.u_wallace._0671_ ),
    .B2(\u_cpu.ALU.u_wallace._0659_ ),
    .X(\u_cpu.ALU.u_wallace._0672_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6455_  (.A1(\u_cpu.ALU.u_wallace._0660_ ),
    .A2(\u_cpu.ALU.u_wallace._0666_ ),
    .B1(\u_cpu.ALU.u_wallace._0668_ ),
    .C1(\u_cpu.ALU.u_wallace._0672_ ),
    .X(\u_cpu.ALU.u_wallace._0673_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6456_  (.A(\u_cpu.ALU.u_wallace._0656_ ),
    .B(\u_cpu.ALU.u_wallace._0650_ ),
    .C(\u_cpu.ALU.u_wallace._0655_ ),
    .Y(\u_cpu.ALU.u_wallace._0674_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._6457_  (.A1(\u_cpu.ALU.u_wallace._0674_ ),
    .A2(\u_cpu.ALU.u_wallace._0664_ ),
    .B1_N(\u_cpu.ALU.u_wallace._0658_ ),
    .Y(\u_cpu.ALU.u_wallace._0675_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6458_  (.A1(\u_cpu.ALU.u_wallace._0620_ ),
    .A2(\u_cpu.ALU.u_wallace._0625_ ),
    .B1(\u_cpu.ALU.u_wallace._0666_ ),
    .B2(\u_cpu.ALU.u_wallace._0675_ ),
    .Y(\u_cpu.ALU.u_wallace._0677_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6459_  (.A1(\u_cpu.ALU.u_wallace._0669_ ),
    .A2(\u_cpu.ALU.u_wallace._0670_ ),
    .B1(\u_cpu.ALU.u_wallace._0671_ ),
    .C1(\u_cpu.ALU.u_wallace._0659_ ),
    .Y(\u_cpu.ALU.u_wallace._0678_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._6460_  (.A1(\u_cpu.ALU.u_wallace._0484_ ),
    .A2(\u_cpu.ALU.u_wallace._0478_ ),
    .A3(\u_cpu.ALU.u_wallace._0482_ ),
    .B1(\u_cpu.ALU.u_wallace._0667_ ),
    .Y(\u_cpu.ALU.u_wallace._0679_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6461_  (.A(\u_cpu.ALU.u_wallace._0677_ ),
    .B(\u_cpu.ALU.u_wallace._0678_ ),
    .C(\u_cpu.ALU.u_wallace._0679_ ),
    .Y(\u_cpu.ALU.u_wallace._0680_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._6462_  (.A1(\u_cpu.ALU.u_wallace._0502_ ),
    .A2(\u_cpu.ALU.u_wallace._0504_ ),
    .B1(\u_cpu.ALU.u_wallace._0509_ ),
    .X(\u_cpu.ALU.u_wallace._0681_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6463_  (.A1(\u_cpu.ALU.u_wallace._4594_ ),
    .A2(\u_cpu.ALU.u_wallace._4439_ ),
    .B1(\u_cpu.ALU.u_wallace._4595_ ),
    .B2(\u_cpu.ALU.u_wallace._3623_ ),
    .X(\u_cpu.ALU.u_wallace._0682_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6464_  (.A(\u_cpu.ALU.u_wallace._3689_ ),
    .B(\u_cpu.ALU.u_wallace._4716_ ),
    .C(\u_cpu.ALU.u_wallace._4562_ ),
    .D(\u_cpu.ALU.u_wallace._0045_ ),
    .Y(\u_cpu.ALU.u_wallace._0683_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6465_  (.A1(\u_cpu.ALU.u_wallace._2801_ ),
    .A2(\u_cpu.ALU.u_wallace._0052_ ),
    .B1(\u_cpu.ALU.u_wallace._0682_ ),
    .B2(\u_cpu.ALU.u_wallace._0683_ ),
    .Y(\u_cpu.ALU.u_wallace._0684_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6466_  (.A1(\u_cpu.ALU.u_wallace._4720_ ),
    .A2(\u_cpu.ALU.u_wallace._4439_ ),
    .B1(\u_cpu.ALU.u_wallace._4595_ ),
    .B2(\u_cpu.ALU.u_wallace._3623_ ),
    .Y(\u_cpu.ALU.u_wallace._0685_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6467_  (.A(\u_cpu.ALU.u_wallace._0683_ ),
    .B(\u_cpu.ALU.u_wallace._4604_ ),
    .C(\u_cpu.ALU.u_wallace._2801_ ),
    .Y(\u_cpu.ALU.u_wallace._0686_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._6468_  (.A(\u_cpu.ALU.u_wallace._0685_ ),
    .B(\u_cpu.ALU.u_wallace._0686_ ),
    .Y(\u_cpu.ALU.u_wallace._0688_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6469_  (.A1(\u_cpu.ALU.u_wallace._1793_ ),
    .A2(\u_cpu.ALU.u_wallace._0364_ ),
    .B1(\u_cpu.ALU.u_wallace._0365_ ),
    .B2(\u_cpu.ALU.u_wallace._2955_ ),
    .X(\u_cpu.ALU.u_wallace._0689_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6470_  (.A(\u_cpu.ALU.u_wallace._3832_ ),
    .B(\u_cpu.ALU.u_wallace._1125_ ),
    .C(\u_cpu.ALU.u_wallace._0028_ ),
    .D(\u_cpu.ALU.u_wallace._0144_ ),
    .Y(\u_cpu.ALU.u_wallace._0690_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6471_  (.A1(\u_cpu.ALU.u_wallace._2933_ ),
    .A2(\u_cpu.ALU.u_wallace._0057_ ),
    .B1(\u_cpu.ALU.u_wallace._0689_ ),
    .B2(\u_cpu.ALU.u_wallace._0690_ ),
    .Y(\u_cpu.ALU.u_wallace._0691_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6472_  (.A(\u_cpu.ALU.u_wallace._0689_ ),
    .B(\u_cpu.ALU.u_wallace._0690_ ),
    .C(\u_cpu.ALU.u_wallace._2933_ ),
    .D(\u_cpu.ALU.u_wallace._0363_ ),
    .X(\u_cpu.ALU.u_wallace._0692_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._6473_  (.A(\u_cpu.ALU.u_wallace._0691_ ),
    .B(\u_cpu.ALU.u_wallace._0692_ ),
    .Y(\u_cpu.ALU.u_wallace._0693_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6474_  (.A1(\u_cpu.ALU.u_wallace._0684_ ),
    .A2(\u_cpu.ALU.u_wallace._0688_ ),
    .B1(\u_cpu.ALU.u_wallace._0681_ ),
    .Y(\u_cpu.ALU.u_wallace._0694_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU.u_wallace._6475_  (.A1(\u_cpu.ALU.u_wallace._0681_ ),
    .A2(\u_cpu.ALU.u_wallace._0684_ ),
    .A3(\u_cpu.ALU.u_wallace._0688_ ),
    .B1(\u_cpu.ALU.u_wallace._0693_ ),
    .C1(\u_cpu.ALU.u_wallace._0694_ ),
    .X(\u_cpu.ALU.u_wallace._0695_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6476_  (.A1(\u_cpu.ALU.u_wallace._0467_ ),
    .A2(\u_cpu.ALU.u_wallace._0481_ ),
    .B1(\u_cpu.ALU.u_wallace._0474_ ),
    .Y(\u_cpu.ALU.u_wallace._0696_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6477_  (.A1(\u_cpu.ALU.u_wallace._0502_ ),
    .A2(\u_cpu.ALU.u_wallace._0504_ ),
    .B1(\u_cpu.ALU.u_wallace._0509_ ),
    .Y(\u_cpu.ALU.u_wallace._0697_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6478_  (.A1(\u_cpu.ALU.u_wallace._4698_ ),
    .A2(\u_cpu.ALU.u_wallace._4610_ ),
    .B1(\u_cpu.ALU.u_wallace._0682_ ),
    .B2(\u_cpu.ALU.u_wallace._0683_ ),
    .X(\u_cpu.ALU.u_wallace._0699_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6479_  (.A1(\u_cpu.ALU.u_wallace._0686_ ),
    .A2(\u_cpu.ALU.u_wallace._0685_ ),
    .B1(\u_cpu.ALU.u_wallace._0697_ ),
    .C1(\u_cpu.ALU.u_wallace._0699_ ),
    .Y(\u_cpu.ALU.u_wallace._0700_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6480_  (.A1_N(\u_cpu.ALU.u_wallace._0700_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0694_ ),
    .B1(\u_cpu.ALU.u_wallace._0691_ ),
    .B2(\u_cpu.ALU.u_wallace._0692_ ),
    .Y(\u_cpu.ALU.u_wallace._0701_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6481_  (.A(\u_cpu.ALU.u_wallace._0696_ ),
    .B(\u_cpu.ALU.u_wallace._0701_ ),
    .Y(\u_cpu.ALU.u_wallace._0702_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6482_  (.A1(\u_cpu.ALU.u_wallace._0700_ ),
    .A2(\u_cpu.ALU.u_wallace._0694_ ),
    .B1(\u_cpu.ALU.u_wallace._0693_ ),
    .Y(\u_cpu.ALU.u_wallace._0703_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._6483_  (.A1(\u_cpu.ALU.u_wallace._0695_ ),
    .A2(\u_cpu.ALU.u_wallace._0703_ ),
    .B1_N(\u_cpu.ALU.u_wallace._0696_ ),
    .Y(\u_cpu.ALU.u_wallace._0704_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6484_  (.A1(\u_cpu.ALU.u_wallace._0500_ ),
    .A2(\u_cpu.ALU.u_wallace._0511_ ),
    .B1(\u_cpu.ALU.u_wallace._0514_ ),
    .X(\u_cpu.ALU.u_wallace._0705_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6485_  (.A1(\u_cpu.ALU.u_wallace._0695_ ),
    .A2(\u_cpu.ALU.u_wallace._0702_ ),
    .B1(\u_cpu.ALU.u_wallace._0704_ ),
    .C1(\u_cpu.ALU.u_wallace._0705_ ),
    .Y(\u_cpu.ALU.u_wallace._0706_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6486_  (.A1(\u_cpu.ALU.u_wallace._0686_ ),
    .A2(\u_cpu.ALU.u_wallace._0685_ ),
    .B1(\u_cpu.ALU.u_wallace._0697_ ),
    .C1(\u_cpu.ALU.u_wallace._0699_ ),
    .X(\u_cpu.ALU.u_wallace._0707_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6487_  (.A(\u_cpu.ALU.u_wallace._0694_ ),
    .B(\u_cpu.ALU.u_wallace._0693_ ),
    .Y(\u_cpu.ALU.u_wallace._0708_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6488_  (.A1(\u_cpu.ALU.u_wallace._0707_ ),
    .A2(\u_cpu.ALU.u_wallace._0708_ ),
    .B1(\u_cpu.ALU.u_wallace._0701_ ),
    .C1(\u_cpu.ALU.u_wallace._0696_ ),
    .Y(\u_cpu.ALU.u_wallace._0710_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6489_  (.A1(\u_cpu.ALU.u_wallace._0710_ ),
    .A2(\u_cpu.ALU.u_wallace._0704_ ),
    .B1(\u_cpu.ALU.u_wallace._0705_ ),
    .X(\u_cpu.ALU.u_wallace._0711_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6490_  (.A(\u_cpu.ALU.u_wallace._0680_ ),
    .B(\u_cpu.ALU.u_wallace._0706_ ),
    .C(\u_cpu.ALU.u_wallace._0711_ ),
    .Y(\u_cpu.ALU.u_wallace._0712_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6491_  (.A1(\u_cpu.ALU.u_wallace._0660_ ),
    .A2(\u_cpu.ALU.u_wallace._0666_ ),
    .B1(\u_cpu.ALU.u_wallace._0668_ ),
    .C1(\u_cpu.ALU.u_wallace._0672_ ),
    .Y(\u_cpu.ALU.u_wallace._0713_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6492_  (.A(\u_cpu.ALU.u_wallace._0705_ ),
    .B(\u_cpu.ALU.u_wallace._0710_ ),
    .C(\u_cpu.ALU.u_wallace._0704_ ),
    .X(\u_cpu.ALU.u_wallace._0714_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6493_  (.A1(\u_cpu.ALU.u_wallace._0710_ ),
    .A2(\u_cpu.ALU.u_wallace._0704_ ),
    .B1(\u_cpu.ALU.u_wallace._0705_ ),
    .Y(\u_cpu.ALU.u_wallace._0715_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6494_  (.A1_N(\u_cpu.ALU.u_wallace._0713_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0680_ ),
    .B1(\u_cpu.ALU.u_wallace._0714_ ),
    .B2(\u_cpu.ALU.u_wallace._0715_ ),
    .Y(\u_cpu.ALU.u_wallace._0716_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6495_  (.A1(\u_cpu.ALU.u_wallace._0493_ ),
    .A2(\u_cpu.ALU.u_wallace._0529_ ),
    .B1(\u_cpu.ALU.u_wallace._0530_ ),
    .Y(\u_cpu.ALU.u_wallace._0717_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6496_  (.A1(\u_cpu.ALU.u_wallace._0673_ ),
    .A2(\u_cpu.ALU.u_wallace._0712_ ),
    .B1(\u_cpu.ALU.u_wallace._0716_ ),
    .C1(\u_cpu.ALU.u_wallace._0717_ ),
    .Y(\u_cpu.ALU.u_wallace._0718_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6497_  (.A(\u_cpu.ALU.u_wallace._0706_ ),
    .B(\u_cpu.ALU.u_wallace._0711_ ),
    .Y(\u_cpu.ALU.u_wallace._0719_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6498_  (.A(\u_cpu.ALU.u_wallace._0713_ ),
    .B(\u_cpu.ALU.u_wallace._0680_ ),
    .Y(\u_cpu.ALU.u_wallace._0721_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6499_  (.A1_N(\u_cpu.ALU.u_wallace._0719_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0721_ ),
    .B1(\u_cpu.ALU.u_wallace._0673_ ),
    .B2(\u_cpu.ALU.u_wallace._0712_ ),
    .Y(\u_cpu.ALU.u_wallace._0722_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._6500_  (.A1(\u_cpu.ALU.u_wallace._0493_ ),
    .A2(\u_cpu.ALU.u_wallace._0529_ ),
    .B1(\u_cpu.ALU.u_wallace._0530_ ),
    .X(\u_cpu.ALU.u_wallace._0723_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6501_  (.A(\u_cpu.ALU.u_wallace._4529_ ),
    .B(\u_cpu.ALU.u_wallace._1180_ ),
    .C(\u_cpu.ALU.u_wallace._0028_ ),
    .D(\u_cpu.ALU.u_wallace._0029_ ),
    .X(\u_cpu.ALU.u_wallace._0724_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6502_  (.A1(\u_cpu.ALU.u_wallace._4529_ ),
    .A2(\u_cpu.ALU.u_wallace._4837_ ),
    .B1(\u_cpu.ALU.u_wallace._4838_ ),
    .B2(\u_cpu.ALU.u_wallace._0906_ ),
    .Y(\u_cpu.ALU.u_wallace._0725_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._6503_  (.A(\u_cpu.ALU.u_wallace._0497_ ),
    .B(\u_cpu.ALU.u_wallace._0725_ ),
    .Y(\u_cpu.ALU.u_wallace._0726_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6504_  (.A(\u_cpu.ALU.SrcB[14] ),
    .X(\u_cpu.ALU.u_wallace._0727_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6505_  (.A(\u_cpu.ALU.SrcB[15] ),
    .X(\u_cpu.ALU.u_wallace._0728_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6506_  (.A1(\u_cpu.ALU.u_wallace._2549_ ),
    .A2(\u_cpu.ALU.u_wallace._0727_ ),
    .B1(\u_cpu.ALU.u_wallace._0728_ ),
    .B2(\u_cpu.ALU.u_wallace._0392_ ),
    .X(\u_cpu.ALU.u_wallace._0729_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6507_  (.A(\u_cpu.ALU.SrcB[14] ),
    .X(\u_cpu.ALU.u_wallace._0730_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6508_  (.A(\u_cpu.ALU.SrcB[15] ),
    .X(\u_cpu.ALU.u_wallace._0732_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6509_  (.A(\u_cpu.ALU.u_wallace._0512_ ),
    .B(\u_cpu.ALU.u_wallace._1278_ ),
    .C(\u_cpu.ALU.u_wallace._0730_ ),
    .D(\u_cpu.ALU.u_wallace._0732_ ),
    .Y(\u_cpu.ALU.u_wallace._0733_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6510_  (.A(\u_cpu.ALU.u_wallace._0729_ ),
    .B(\u_cpu.ALU.u_wallace._0733_ ),
    .C(\u_cpu.ALU.u_wallace._1454_ ),
    .D(\u_cpu.ALU.u_wallace._0550_ ),
    .Y(\u_cpu.ALU.u_wallace._0734_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6511_  (.A(\u_cpu.ALU.u_wallace._0550_ ),
    .X(\u_cpu.ALU.u_wallace._0735_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6512_  (.A1(\u_cpu.ALU.u_wallace._1278_ ),
    .A2(\u_cpu.ALU.u_wallace._0730_ ),
    .B1(\u_cpu.ALU.u_wallace._0547_ ),
    .B2(\u_cpu.ALU.u_wallace._0348_ ),
    .Y(\u_cpu.ALU.u_wallace._0736_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6513_  (.A(\u_cpu.ALU.u_wallace._0392_ ),
    .B(\u_cpu.ALU.u_wallace._2549_ ),
    .C(\u_cpu.ALU.u_wallace._0727_ ),
    .D(\u_cpu.ALU.u_wallace._0278_ ),
    .X(\u_cpu.ALU.u_wallace._0737_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6514_  (.A1_N(\u_cpu.ALU.u_wallace._0261_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0735_ ),
    .B1(\u_cpu.ALU.u_wallace._0736_ ),
    .B2(\u_cpu.ALU.u_wallace._0737_ ),
    .Y(\u_cpu.ALU.u_wallace._0738_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6515_  (.A1(\u_cpu.ALU.u_wallace._0724_ ),
    .A2(\u_cpu.ALU.u_wallace._0726_ ),
    .B1(\u_cpu.ALU.u_wallace._0734_ ),
    .C1(\u_cpu.ALU.u_wallace._0738_ ),
    .X(\u_cpu.ALU.u_wallace._0739_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6516_  (.A1(\u_cpu.ALU.u_wallace._0558_ ),
    .A2(\u_cpu.ALU.u_wallace._0555_ ),
    .B1(\u_cpu.ALU.u_wallace._0552_ ),
    .Y(\u_cpu.ALU.u_wallace._0740_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._6517_  (.A1(\u_cpu.ALU.u_wallace._0495_ ),
    .A2(\u_cpu.ALU.u_wallace._0057_ ),
    .A3(\u_cpu.ALU.u_wallace._4541_ ),
    .B1(\u_cpu.ALU.u_wallace._0724_ ),
    .X(\u_cpu.ALU.u_wallace._0741_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6518_  (.A1(\u_cpu.ALU.u_wallace._0734_ ),
    .A2(\u_cpu.ALU.u_wallace._0738_ ),
    .B1(\u_cpu.ALU.u_wallace._0741_ ),
    .X(\u_cpu.ALU.u_wallace._0743_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._6519_  (.A_N(\u_cpu.ALU.u_wallace._0739_ ),
    .B(\u_cpu.ALU.u_wallace._0740_ ),
    .C(\u_cpu.ALU.u_wallace._0743_ ),
    .Y(\u_cpu.ALU.u_wallace._0744_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6520_  (.A1(\u_cpu.ALU.u_wallace._0734_ ),
    .A2(\u_cpu.ALU.u_wallace._0738_ ),
    .B1(\u_cpu.ALU.u_wallace._0741_ ),
    .Y(\u_cpu.ALU.u_wallace._0745_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._6521_  (.A1(\u_cpu.ALU.u_wallace._0739_ ),
    .A2(\u_cpu.ALU.u_wallace._0745_ ),
    .B1_N(\u_cpu.ALU.u_wallace._0740_ ),
    .Y(\u_cpu.ALU.u_wallace._0746_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6522_  (.A(\u_cpu.ALU.u_wallace._1070_ ),
    .B(\u_cpu.ALU.u_wallace._0272_ ),
    .C(\u_cpu.ALU.u_wallace._0122_ ),
    .D(\u_cpu.ALU.u_wallace._0280_ ),
    .X(\u_cpu.ALU.u_wallace._0747_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6523_  (.A1(\u_cpu.ALU.u_wallace._0552_ ),
    .A2(\u_cpu.ALU.u_wallace._0560_ ),
    .B1(\u_cpu.ALU.u_wallace._0563_ ),
    .X(\u_cpu.ALU.u_wallace._0748_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._6524_  (.A1(\u_cpu.ALU.u_wallace._0747_ ),
    .A2(\u_cpu.ALU.u_wallace._0565_ ),
    .B1(\u_cpu.ALU.u_wallace._0748_ ),
    .X(\u_cpu.ALU.u_wallace._0749_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6525_  (.A1(\u_cpu.ALU.u_wallace._0744_ ),
    .A2(\u_cpu.ALU.u_wallace._0746_ ),
    .B1(\u_cpu.ALU.u_wallace._0749_ ),
    .X(\u_cpu.ALU.u_wallace._0750_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._6526_  (.A1(\u_cpu.ALU.u_wallace._0747_ ),
    .A2(\u_cpu.ALU.u_wallace._0565_ ),
    .B1(\u_cpu.ALU.u_wallace._0744_ ),
    .C1(\u_cpu.ALU.u_wallace._0746_ ),
    .D1(\u_cpu.ALU.u_wallace._0748_ ),
    .Y(\u_cpu.ALU.u_wallace._0751_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6527_  (.A1(\u_cpu.ALU.u_wallace._0517_ ),
    .A2(\u_cpu.ALU.u_wallace._0541_ ),
    .B1(\u_cpu.ALU.u_wallace._0750_ ),
    .C1(\u_cpu.ALU.u_wallace._0751_ ),
    .Y(\u_cpu.ALU.u_wallace._0752_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6528_  (.A1(\u_cpu.ALU.u_wallace._0744_ ),
    .A2(\u_cpu.ALU.u_wallace._0746_ ),
    .B1(\u_cpu.ALU.u_wallace._0749_ ),
    .Y(\u_cpu.ALU.u_wallace._0754_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._6529_  (.A1(\u_cpu.ALU.u_wallace._0747_ ),
    .A2(\u_cpu.ALU.u_wallace._0565_ ),
    .B1(\u_cpu.ALU.u_wallace._0744_ ),
    .C1(\u_cpu.ALU.u_wallace._0746_ ),
    .D1(\u_cpu.ALU.u_wallace._0748_ ),
    .X(\u_cpu.ALU.u_wallace._0755_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6530_  (.A1(\u_cpu.ALU.u_wallace._0754_ ),
    .A2(\u_cpu.ALU.u_wallace._0755_ ),
    .B1(\u_cpu.ALU.u_wallace._0525_ ),
    .C1(\u_cpu.ALU.u_wallace._0522_ ),
    .Y(\u_cpu.ALU.u_wallace._0756_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.ALU.u_wallace._6531_  (.A(\u_cpu.ALU.u_wallace._0287_ ),
    .B(\u_cpu.ALU.u_wallace._0564_ ),
    .C(\u_cpu.ALU.u_wallace._0565_ ),
    .X(\u_cpu.ALU.u_wallace._0757_ ));
 sky130_fd_sc_hd__a21bo_2 \u_cpu.ALU.u_wallace._6532_  (.A1(\u_cpu.ALU.u_wallace._0752_ ),
    .A2(\u_cpu.ALU.u_wallace._0756_ ),
    .B1_N(\u_cpu.ALU.u_wallace._0757_ ),
    .X(\u_cpu.ALU.u_wallace._0758_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._6533_  (.A_N(\u_cpu.ALU.u_wallace._0757_ ),
    .B(\u_cpu.ALU.u_wallace._0752_ ),
    .C(\u_cpu.ALU.u_wallace._0756_ ),
    .Y(\u_cpu.ALU.u_wallace._0759_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6534_  (.A(\u_cpu.ALU.u_wallace._0758_ ),
    .B(\u_cpu.ALU.u_wallace._0759_ ),
    .Y(\u_cpu.ALU.u_wallace._0760_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6535_  (.A1(\u_cpu.ALU.u_wallace._0722_ ),
    .A2(\u_cpu.ALU.u_wallace._0723_ ),
    .B1(\u_cpu.ALU.u_wallace._0760_ ),
    .Y(\u_cpu.ALU.u_wallace._0761_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6536_  (.A(\u_cpu.ALU.u_wallace._0713_ ),
    .B(\u_cpu.ALU.u_wallace._0680_ ),
    .C(\u_cpu.ALU.u_wallace._0706_ ),
    .D(\u_cpu.ALU.u_wallace._0711_ ),
    .Y(\u_cpu.ALU.u_wallace._0762_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6537_  (.A1(\u_cpu.ALU.u_wallace._0762_ ),
    .A2(\u_cpu.ALU.u_wallace._0716_ ),
    .B1(\u_cpu.ALU.u_wallace._0717_ ),
    .X(\u_cpu.ALU.u_wallace._0763_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6538_  (.A(\u_cpu.ALU.u_wallace._0718_ ),
    .B(\u_cpu.ALU.u_wallace._0763_ ),
    .Y(\u_cpu.ALU.u_wallace._0765_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6539_  (.A1(\u_cpu.ALU.u_wallace._0718_ ),
    .A2(\u_cpu.ALU.u_wallace._0761_ ),
    .B1(\u_cpu.ALU.u_wallace._0765_ ),
    .B2(\u_cpu.ALU.u_wallace._0760_ ),
    .Y(\u_cpu.ALU.u_wallace._0766_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6540_  (.A1(\u_cpu.ALU.u_wallace._0604_ ),
    .A2(\u_cpu.ALU.u_wallace._0583_ ),
    .B1(\u_cpu.ALU.u_wallace._0766_ ),
    .Y(\u_cpu.ALU.u_wallace._0767_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6541_  (.A(\u_cpu.ALU.u_wallace._0286_ ),
    .B(\u_cpu.ALU.u_wallace._0287_ ),
    .C(\u_cpu.ALU.u_wallace._0572_ ),
    .D(\u_cpu.ALU.u_wallace._0123_ ),
    .X(\u_cpu.ALU.u_wallace._0768_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6542_  (.A1(\u_cpu.ALU.u_wallace._0577_ ),
    .A2(\u_cpu.ALU.u_wallace._0536_ ),
    .B1(\u_cpu.ALU.u_wallace._0604_ ),
    .X(\u_cpu.ALU.u_wallace._0769_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6543_  (.A1(\u_cpu.ALU.u_wallace._0570_ ),
    .A2(\u_cpu.ALU.u_wallace._0768_ ),
    .B1(\u_cpu.ALU.u_wallace._0769_ ),
    .B2(\u_cpu.ALU.u_wallace._0766_ ),
    .Y(\u_cpu.ALU.u_wallace._0770_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.ALU.u_wallace._6544_  (.A1(\u_cpu.ALU.u_wallace._0604_ ),
    .A2(\u_cpu.ALU.u_wallace._0605_ ),
    .A3(\u_cpu.ALU.u_wallace._0766_ ),
    .B1(\u_cpu.ALU.u_wallace._0767_ ),
    .C1(\u_cpu.ALU.u_wallace._0770_ ),
    .Y(\u_cpu.ALU.u_wallace._0771_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6545_  (.A1(\u_cpu.ALU.u_wallace._0579_ ),
    .A2(\u_cpu.ALU.u_wallace._0580_ ),
    .B1(\u_cpu.ALU.u_wallace._0437_ ),
    .Y(\u_cpu.ALU.u_wallace._0772_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._6546_  (.A1(\u_cpu.ALU.u_wallace._0585_ ),
    .A2(\u_cpu.ALU.u_wallace._0289_ ),
    .A3(\u_cpu.ALU.u_wallace._0772_ ),
    .B1(\u_cpu.ALU.u_wallace._0581_ ),
    .X(\u_cpu.ALU.u_wallace._0773_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._6547_  (.A_N(\u_cpu.ALU.u_wallace._0760_ ),
    .B(\u_cpu.ALU.u_wallace._0763_ ),
    .C(\u_cpu.ALU.u_wallace._0718_ ),
    .Y(\u_cpu.ALU.u_wallace._0774_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6548_  (.A1(\u_cpu.ALU.u_wallace._0673_ ),
    .A2(\u_cpu.ALU.u_wallace._0712_ ),
    .B1(\u_cpu.ALU.u_wallace._0716_ ),
    .C1(\u_cpu.ALU.u_wallace._0717_ ),
    .X(\u_cpu.ALU.u_wallace._0776_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6549_  (.A1(\u_cpu.ALU.u_wallace._0762_ ),
    .A2(\u_cpu.ALU.u_wallace._0716_ ),
    .B1(\u_cpu.ALU.u_wallace._0717_ ),
    .Y(\u_cpu.ALU.u_wallace._0777_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6550_  (.A1(\u_cpu.ALU.u_wallace._0776_ ),
    .A2(\u_cpu.ALU.u_wallace._0777_ ),
    .B1(\u_cpu.ALU.u_wallace._0760_ ),
    .Y(\u_cpu.ALU.u_wallace._0778_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6551_  (.A1(\u_cpu.ALU.u_wallace._0604_ ),
    .A2(\u_cpu.ALU.u_wallace._0605_ ),
    .B1(\u_cpu.ALU.u_wallace._0774_ ),
    .C1(\u_cpu.ALU.u_wallace._0778_ ),
    .X(\u_cpu.ALU.u_wallace._0779_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6552_  (.A1(\u_cpu.ALU.u_wallace._0774_ ),
    .A2(\u_cpu.ALU.u_wallace._0778_ ),
    .B1(\u_cpu.ALU.u_wallace._0769_ ),
    .Y(\u_cpu.ALU.u_wallace._0780_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6553_  (.A1(\u_cpu.ALU.u_wallace._0570_ ),
    .A2(\u_cpu.ALU.u_wallace._0768_ ),
    .B1(\u_cpu.ALU.u_wallace._0779_ ),
    .B2(\u_cpu.ALU.u_wallace._0780_ ),
    .Y(\u_cpu.ALU.u_wallace._0781_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6554_  (.A(\u_cpu.ALU.u_wallace._0771_ ),
    .B(\u_cpu.ALU.u_wallace._0773_ ),
    .C(\u_cpu.ALU.u_wallace._0781_ ),
    .Y(\u_cpu.ALU.u_wallace._0782_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._6555_  (.A1(\u_cpu.ALU.u_wallace._0437_ ),
    .A2(\u_cpu.ALU.u_wallace._0579_ ),
    .A3(\u_cpu.ALU.u_wallace._0580_ ),
    .B1(\u_cpu.ALU.u_wallace._0584_ ),
    .B2(\u_cpu.ALU.u_wallace._0587_ ),
    .X(\u_cpu.ALU.u_wallace._0783_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._6556_  (.A(\u_cpu.ALU.u_wallace._0570_ ),
    .B(\u_cpu.ALU.u_wallace._0768_ ),
    .Y(\u_cpu.ALU.u_wallace._0784_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6557_  (.A1(\u_cpu.ALU.u_wallace._0779_ ),
    .A2(\u_cpu.ALU.u_wallace._0780_ ),
    .B1(\u_cpu.ALU.u_wallace._0784_ ),
    .Y(\u_cpu.ALU.u_wallace._0785_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6558_  (.A1(\u_cpu.ALU.u_wallace._0770_ ),
    .A2(\u_cpu.ALU.u_wallace._0779_ ),
    .B1(\u_cpu.ALU.u_wallace._0783_ ),
    .C1(\u_cpu.ALU.u_wallace._0785_ ),
    .Y(\u_cpu.ALU.u_wallace._0787_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6559_  (.A1(\u_cpu.ALU.u_wallace._0434_ ),
    .A2(\u_cpu.ALU.u_wallace._0603_ ),
    .B1(\u_cpu.ALU.u_wallace._0782_ ),
    .C1(\u_cpu.ALU.u_wallace._0787_ ),
    .Y(\u_cpu.ALU.u_wallace._0788_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6560_  (.A1(\u_cpu.ALU.u_wallace._0128_ ),
    .A2(\u_cpu.ALU.u_wallace._0415_ ),
    .B1(\u_cpu.ALU.u_wallace._0590_ ),
    .Y(\u_cpu.ALU.u_wallace._0789_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6561_  (.A1(\u_cpu.ALU.u_wallace._0581_ ),
    .A2(\u_cpu.ALU.u_wallace._0584_ ),
    .B1(\u_cpu.ALU.u_wallace._0408_ ),
    .X(\u_cpu.ALU.u_wallace._0790_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6562_  (.A1(\u_cpu.ALU.u_wallace._0585_ ),
    .A2(\u_cpu.ALU.u_wallace._0289_ ),
    .B1(\u_cpu.ALU.u_wallace._0581_ ),
    .C1(\u_cpu.ALU.u_wallace._0584_ ),
    .Y(\u_cpu.ALU.u_wallace._0791_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._6563_  (.A1(\u_cpu.ALU.u_wallace._0789_ ),
    .A2(\u_cpu.ALU.u_wallace._0790_ ),
    .A3(\u_cpu.ALU.u_wallace._0791_ ),
    .B1(\u_cpu.ALU.u_wallace._0434_ ),
    .Y(\u_cpu.ALU.u_wallace._0792_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6564_  (.A(\u_cpu.ALU.u_wallace._0782_ ),
    .B(\u_cpu.ALU.u_wallace._0787_ ),
    .Y(\u_cpu.ALU.u_wallace._0793_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6565_  (.A1(\u_cpu.ALU.u_wallace._0602_ ),
    .A2(\u_cpu.ALU.u_wallace._0792_ ),
    .B1(\u_cpu.ALU.u_wallace._0793_ ),
    .Y(\u_cpu.ALU.u_wallace._0794_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6566_  (.A1(\u_cpu.ALU.u_wallace._0602_ ),
    .A2(\u_cpu.ALU.u_wallace._0788_ ),
    .B1(\u_cpu.ALU.u_wallace._0794_ ),
    .Y(\u_cpu.ALU.u_wallace._0795_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.ALU.u_wallace._6567_  (.A1_N(\u_cpu.ALU.u_wallace._0430_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0594_ ),
    .B1(\u_cpu.ALU.u_wallace._0595_ ),
    .B2(\u_cpu.ALU.u_wallace._0601_ ),
    .X(\u_cpu.ALU.u_wallace._0796_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._6568_  (.A(\u_cpu.ALU.u_wallace._0795_ ),
    .B(\u_cpu.ALU.u_wallace._0796_ ),
    .X(\u_cpu.ALU.Product_Wallace[17] ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._6569_  (.A1(\u_cpu.ALU.u_wallace._0771_ ),
    .A2(\u_cpu.ALU.u_wallace._0773_ ),
    .A3(\u_cpu.ALU.u_wallace._0781_ ),
    .B1(\u_cpu.ALU.u_wallace._0593_ ),
    .X(\u_cpu.ALU.u_wallace._0798_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6570_  (.A1(\u_cpu.ALU.u_wallace._0784_ ),
    .A2(\u_cpu.ALU.u_wallace._0780_ ),
    .B1(\u_cpu.ALU.u_wallace._0767_ ),
    .Y(\u_cpu.ALU.u_wallace._0799_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6571_  (.A1(\u_cpu.ALU.u_wallace._1815_ ),
    .A2(\u_cpu.ALU.SrcA[12] ),
    .B1(\u_cpu.ALU.u_wallace._0626_ ),
    .B2(\u_cpu.ALU.u_wallace._0140_ ),
    .Y(\u_cpu.ALU.u_wallace._0800_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6572_  (.A(\u_cpu.ALU.u_wallace._4649_ ),
    .B(\u_cpu.ALU.u_wallace._0140_ ),
    .C(\u_cpu.ALU.u_wallace._4790_ ),
    .D(\u_cpu.ALU.u_wallace._0626_ ),
    .Y(\u_cpu.ALU.u_wallace._0801_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6573_  (.A(\u_cpu.ALU.SrcA[18] ),
    .X(\u_cpu.ALU.u_wallace._0802_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6574_  (.A(\u_cpu.ALU.u_wallace._0801_ ),
    .B(\u_cpu.ALU.u_wallace._0802_ ),
    .C(\u_cpu.ALU.u_wallace._1859_ ),
    .Y(\u_cpu.ALU.u_wallace._0803_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6575_  (.A(\u_cpu.ALU.u_wallace._1771_ ),
    .B(\u_cpu.ALU.u_wallace._4647_ ),
    .Y(\u_cpu.ALU.u_wallace._0804_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6576_  (.A(\u_cpu.ALU.u_wallace._0010_ ),
    .B(\u_cpu.ALU.u_wallace._0639_ ),
    .Y(\u_cpu.ALU.u_wallace._0805_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6577_  (.A1(\u_cpu.ALU.u_wallace._0804_ ),
    .A2(\u_cpu.ALU.u_wallace._0805_ ),
    .B1(\u_cpu.ALU.u_wallace._0631_ ),
    .Y(\u_cpu.ALU.u_wallace._0806_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6578_  (.A(\u_cpu.ALU.SrcA[18] ),
    .X(\u_cpu.ALU.u_wallace._0808_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._6579_  (.A(\u_cpu.ALU.u_wallace._0808_ ),
    .Y(\u_cpu.ALU.u_wallace._0809_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6580_  (.A(\u_cpu.ALU.u_wallace._1815_ ),
    .B(\u_cpu.ALU.u_wallace._0140_ ),
    .C(\u_cpu.ALU.SrcA[12] ),
    .D(\u_cpu.ALU.u_wallace._0628_ ),
    .X(\u_cpu.ALU.u_wallace._0810_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6581_  (.A1(\u_cpu.ALU.u_wallace._0634_ ),
    .A2(\u_cpu.ALU.u_wallace._0809_ ),
    .B1(\u_cpu.ALU.u_wallace._0800_ ),
    .B2(\u_cpu.ALU.u_wallace._0810_ ),
    .Y(\u_cpu.ALU.u_wallace._0811_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._6582_  (.A1(\u_cpu.ALU.u_wallace._0800_ ),
    .A2(\u_cpu.ALU.u_wallace._0803_ ),
    .B1(\u_cpu.ALU.u_wallace._0636_ ),
    .B2(\u_cpu.ALU.u_wallace._0806_ ),
    .C1(\u_cpu.ALU.u_wallace._0811_ ),
    .X(\u_cpu.ALU.u_wallace._0812_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6583_  (.A(\u_cpu.ALU.SrcB[17] ),
    .X(\u_cpu.ALU.u_wallace._0813_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6584_  (.A1(\u_cpu.ALU.u_wallace._4649_ ),
    .A2(\u_cpu.ALU.u_wallace._4790_ ),
    .B1(\u_cpu.ALU.u_wallace._0813_ ),
    .B2(\u_cpu.ALU.u_wallace._0140_ ),
    .X(\u_cpu.ALU.u_wallace._0814_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6585_  (.A(\u_cpu.ALU.u_wallace._0808_ ),
    .X(\u_cpu.ALU.u_wallace._0815_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6586_  (.A(\u_cpu.ALU.u_wallace._0814_ ),
    .B(\u_cpu.ALU.u_wallace._0801_ ),
    .C(\u_cpu.ALU.u_wallace._0873_ ),
    .D(\u_cpu.ALU.u_wallace._0815_ ),
    .Y(\u_cpu.ALU.u_wallace._0816_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6587_  (.A1(\u_cpu.ALU.u_wallace._0631_ ),
    .A2(\u_cpu.ALU.u_wallace._0627_ ),
    .B1(\u_cpu.ALU.u_wallace._0641_ ),
    .Y(\u_cpu.ALU.u_wallace._0817_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6588_  (.A1(\u_cpu.ALU.u_wallace._0811_ ),
    .A2(\u_cpu.ALU.u_wallace._0816_ ),
    .B1(\u_cpu.ALU.u_wallace._0817_ ),
    .Y(\u_cpu.ALU.u_wallace._0819_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6589_  (.A(\u_cpu.ALU.u_wallace._1903_ ),
    .B(\u_cpu.ALU.u_wallace._0293_ ),
    .C(\u_cpu.ALU.u_wallace._0447_ ),
    .D(\u_cpu.ALU.u_wallace._0630_ ),
    .Y(\u_cpu.ALU.u_wallace._0820_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6590_  (.A(\u_cpu.ALU.u_wallace._0820_ ),
    .B(\u_cpu.ALU.u_wallace._0325_ ),
    .C(\u_cpu.ALU.u_wallace._0753_ ),
    .X(\u_cpu.ALU.u_wallace._0821_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6591_  (.A1(\u_cpu.ALU.u_wallace._0807_ ),
    .A2(\u_cpu.ALU.u_wallace._0447_ ),
    .B1(\u_cpu.ALU.u_wallace._0630_ ),
    .B2(\u_cpu.ALU.u_wallace._0797_ ),
    .X(\u_cpu.ALU.u_wallace._0822_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6592_  (.A1(\u_cpu.ALU.u_wallace._0840_ ),
    .A2(\u_cpu.ALU.u_wallace._0325_ ),
    .B1(\u_cpu.ALU.u_wallace._0822_ ),
    .B2(\u_cpu.ALU.u_wallace._0820_ ),
    .Y(\u_cpu.ALU.u_wallace._0823_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6593_  (.A1(\u_cpu.ALU.u_wallace._0821_ ),
    .A2(\u_cpu.ALU.u_wallace._0822_ ),
    .B1(\u_cpu.ALU.u_wallace._0823_ ),
    .Y(\u_cpu.ALU.u_wallace._0824_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6594_  (.A1(\u_cpu.ALU.u_wallace._0812_ ),
    .A2(\u_cpu.ALU.u_wallace._0819_ ),
    .B1(\u_cpu.ALU.u_wallace._0824_ ),
    .Y(\u_cpu.ALU.u_wallace._0825_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6595_  (.A(\u_cpu.ALU.u_wallace._0332_ ),
    .X(\u_cpu.ALU.u_wallace._0826_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6596_  (.A(\u_cpu.ALU.u_wallace._0822_ ),
    .B(\u_cpu.ALU.u_wallace._0820_ ),
    .C(\u_cpu.ALU.u_wallace._4662_ ),
    .D(\u_cpu.ALU.u_wallace._0826_ ),
    .X(\u_cpu.ALU.u_wallace._0827_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6597_  (.A1(\u_cpu.ALU.u_wallace._1859_ ),
    .A2(\u_cpu.ALU.u_wallace._0815_ ),
    .B1(\u_cpu.ALU.u_wallace._0814_ ),
    .B2(\u_cpu.ALU.u_wallace._0801_ ),
    .Y(\u_cpu.ALU.u_wallace._0828_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6598_  (.A1(\u_cpu.ALU.u_wallace._0636_ ),
    .A2(\u_cpu.ALU.u_wallace._0806_ ),
    .B1(\u_cpu.ALU.u_wallace._0816_ ),
    .Y(\u_cpu.ALU.u_wallace._0830_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._6599_  (.A(\u_cpu.ALU.u_wallace._0800_ ),
    .B(\u_cpu.ALU.u_wallace._0803_ ),
    .Y(\u_cpu.ALU.u_wallace._0831_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._6600_  (.A1(\u_cpu.ALU.u_wallace._4923_ ),
    .A2(\u_cpu.ALU.u_wallace._0635_ ),
    .A3(\u_cpu.ALU.u_wallace._0627_ ),
    .B1(\u_cpu.ALU.u_wallace._0641_ ),
    .X(\u_cpu.ALU.u_wallace._0832_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6601_  (.A1(\u_cpu.ALU.u_wallace._0828_ ),
    .A2(\u_cpu.ALU.u_wallace._0831_ ),
    .B1(\u_cpu.ALU.u_wallace._0832_ ),
    .Y(\u_cpu.ALU.u_wallace._0833_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._6602_  (.A1(\u_cpu.ALU.u_wallace._0827_ ),
    .A2(\u_cpu.ALU.u_wallace._0823_ ),
    .B1(\u_cpu.ALU.u_wallace._0828_ ),
    .B2(\u_cpu.ALU.u_wallace._0830_ ),
    .C1(\u_cpu.ALU.u_wallace._0833_ ),
    .Y(\u_cpu.ALU.u_wallace._0834_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6603_  (.A1(\u_cpu.ALU.u_wallace._0655_ ),
    .A2(\u_cpu.ALU.u_wallace._0663_ ),
    .B1(\u_cpu.ALU.u_wallace._0825_ ),
    .B2(\u_cpu.ALU.u_wallace._0834_ ),
    .Y(\u_cpu.ALU.u_wallace._0835_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6604_  (.A1(\u_cpu.ALU.u_wallace._1497_ ),
    .A2(\u_cpu.ALU.u_wallace._4909_ ),
    .B1(\u_cpu.ALU.u_wallace._0313_ ),
    .B2(\u_cpu.ALU.u_wallace._1465_ ),
    .Y(\u_cpu.ALU.u_wallace._0836_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6605_  (.A(\u_cpu.ALU.u_wallace._1026_ ),
    .B(\u_cpu.ALU.u_wallace._1541_ ),
    .C(\u_cpu.ALU.u_wallace._4920_ ),
    .D(\u_cpu.ALU.u_wallace._0182_ ),
    .X(\u_cpu.ALU.u_wallace._0837_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6606_  (.A1(\u_cpu.ALU.u_wallace._4470_ ),
    .A2(\u_cpu.ALU.u_wallace._0169_ ),
    .B1(\u_cpu.ALU.u_wallace._0836_ ),
    .B2(\u_cpu.ALU.u_wallace._0837_ ),
    .Y(\u_cpu.ALU.u_wallace._0838_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6607_  (.A1(\u_cpu.ALU.u_wallace._1541_ ),
    .A2(\u_cpu.ALU.u_wallace._4920_ ),
    .B1(\u_cpu.ALU.u_wallace._0182_ ),
    .B2(\u_cpu.ALU.u_wallace._2144_ ),
    .X(\u_cpu.ALU.u_wallace._0839_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6608_  (.A(\u_cpu.ALU.u_wallace._4467_ ),
    .B(\u_cpu.ALU.u_wallace._1497_ ),
    .C(\u_cpu.ALU.u_wallace._4907_ ),
    .D(\u_cpu.ALU.u_wallace._0177_ ),
    .Y(\u_cpu.ALU.u_wallace._0841_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6609_  (.A(\u_cpu.ALU.u_wallace._0839_ ),
    .B(\u_cpu.ALU.u_wallace._0841_ ),
    .C(\u_cpu.ALU.u_wallace._3404_ ),
    .D(\u_cpu.ALU.u_wallace._4794_ ),
    .Y(\u_cpu.ALU.u_wallace._0842_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6610_  (.A(\u_cpu.ALU.u_wallace._0457_ ),
    .B(\u_cpu.ALU.u_wallace._0313_ ),
    .Y(\u_cpu.ALU.u_wallace._0843_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6611_  (.A1(\u_cpu.ALU.u_wallace._4658_ ),
    .A2(\u_cpu.ALU.u_wallace._0330_ ),
    .B1(\u_cpu.ALU.u_wallace._0448_ ),
    .B2(\u_cpu.ALU.u_wallace._4657_ ),
    .Y(\u_cpu.ALU.u_wallace._0844_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6612_  (.A1(\u_cpu.ALU.u_wallace._0843_ ),
    .A2(\u_cpu.ALU.u_wallace._0844_ ),
    .B1(\u_cpu.ALU.u_wallace._0646_ ),
    .Y(\u_cpu.ALU.u_wallace._0845_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6613_  (.A1(\u_cpu.ALU.u_wallace._0838_ ),
    .A2(\u_cpu.ALU.u_wallace._0842_ ),
    .B1(\u_cpu.ALU.u_wallace._0845_ ),
    .X(\u_cpu.ALU.u_wallace._0846_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6614_  (.A(\u_cpu.ALU.u_wallace._4554_ ),
    .X(\u_cpu.ALU.u_wallace._0847_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._6615_  (.A1(\u_cpu.ALU.u_wallace._0611_ ),
    .A2(\u_cpu.ALU.u_wallace._0847_ ),
    .A3(\u_cpu.ALU.u_wallace._3481_ ),
    .B1(\u_cpu.ALU.u_wallace._0615_ ),
    .X(\u_cpu.ALU.u_wallace._0848_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6616_  (.A(\u_cpu.ALU.u_wallace._0846_ ),
    .B(\u_cpu.ALU.u_wallace._0848_ ),
    .Y(\u_cpu.ALU.u_wallace._0849_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6617_  (.A(\u_cpu.ALU.u_wallace._0447_ ),
    .X(\u_cpu.ALU.u_wallace._0850_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6618_  (.A(\u_cpu.ALU.u_wallace._0523_ ),
    .B(\u_cpu.ALU.u_wallace._0545_ ),
    .C(\u_cpu.ALU.u_wallace._0330_ ),
    .D(\u_cpu.ALU.u_wallace._0850_ ),
    .X(\u_cpu.ALU.u_wallace._0852_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._6619_  (.A(\u_cpu.ALU.u_wallace._0843_ ),
    .B(\u_cpu.ALU.u_wallace._0844_ ),
    .Y(\u_cpu.ALU.u_wallace._0853_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6620_  (.A1(\u_cpu.ALU.u_wallace._0852_ ),
    .A2(\u_cpu.ALU.u_wallace._0853_ ),
    .B1(\u_cpu.ALU.u_wallace._0842_ ),
    .C1(\u_cpu.ALU.u_wallace._0838_ ),
    .X(\u_cpu.ALU.u_wallace._0854_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6621_  (.A1(\u_cpu.ALU.u_wallace._0838_ ),
    .A2(\u_cpu.ALU.u_wallace._0842_ ),
    .B1(\u_cpu.ALU.u_wallace._0845_ ),
    .Y(\u_cpu.ALU.u_wallace._0855_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._6622_  (.A1(\u_cpu.ALU.u_wallace._4539_ ),
    .A2(\u_cpu.ALU.u_wallace._4904_ ),
    .A3(\u_cpu.ALU.u_wallace._0614_ ),
    .B1(\u_cpu.ALU.u_wallace._0612_ ),
    .X(\u_cpu.ALU.u_wallace._0856_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6623_  (.A1(\u_cpu.ALU.u_wallace._0855_ ),
    .A2(\u_cpu.ALU.u_wallace._0854_ ),
    .B1(\u_cpu.ALU.u_wallace._0856_ ),
    .Y(\u_cpu.ALU.u_wallace._0857_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6624_  (.A1(\u_cpu.ALU.u_wallace._0656_ ),
    .A2(\u_cpu.ALU.u_wallace._0650_ ),
    .B1(\u_cpu.ALU.u_wallace._0638_ ),
    .Y(\u_cpu.ALU.u_wallace._0858_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6625_  (.A(\u_cpu.ALU.u_wallace._0825_ ),
    .B(\u_cpu.ALU.u_wallace._0834_ ),
    .C(\u_cpu.ALU.u_wallace._0858_ ),
    .Y(\u_cpu.ALU.u_wallace._0859_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6626_  (.A1(\u_cpu.ALU.u_wallace._0849_ ),
    .A2(\u_cpu.ALU.u_wallace._0854_ ),
    .B1(\u_cpu.ALU.u_wallace._0857_ ),
    .C1(\u_cpu.ALU.u_wallace._0859_ ),
    .Y(\u_cpu.ALU.u_wallace._0860_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6627_  (.A1(\u_cpu.ALU.u_wallace._0638_ ),
    .A2(\u_cpu.ALU.u_wallace._0663_ ),
    .B1(\u_cpu.ALU.u_wallace._0664_ ),
    .Y(\u_cpu.ALU.u_wallace._0861_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._6628_  (.A1_N(\u_cpu.ALU.u_wallace._0620_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0625_ ),
    .B1(\u_cpu.ALU.u_wallace._0658_ ),
    .B2(\u_cpu.ALU.u_wallace._0861_ ),
    .Y(\u_cpu.ALU.u_wallace._0863_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6629_  (.A1(\u_cpu.ALU.u_wallace._0852_ ),
    .A2(\u_cpu.ALU.u_wallace._0853_ ),
    .B1(\u_cpu.ALU.u_wallace._0842_ ),
    .C1(\u_cpu.ALU.u_wallace._0838_ ),
    .Y(\u_cpu.ALU.u_wallace._0864_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6630_  (.A1(\u_cpu.ALU.u_wallace._0846_ ),
    .A2(\u_cpu.ALU.u_wallace._0864_ ),
    .B1(\u_cpu.ALU.u_wallace._0848_ ),
    .Y(\u_cpu.ALU.u_wallace._0865_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6631_  (.A(\u_cpu.ALU.u_wallace._0846_ ),
    .B(\u_cpu.ALU.u_wallace._0864_ ),
    .C(\u_cpu.ALU.u_wallace._0848_ ),
    .X(\u_cpu.ALU.u_wallace._0866_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6632_  (.A1(\u_cpu.ALU.u_wallace._0828_ ),
    .A2(\u_cpu.ALU.u_wallace._0830_ ),
    .B1(\u_cpu.ALU.u_wallace._0824_ ),
    .C1(\u_cpu.ALU.u_wallace._0833_ ),
    .Y(\u_cpu.ALU.u_wallace._0867_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6633_  (.A1(\u_cpu.ALU.u_wallace._0827_ ),
    .A2(\u_cpu.ALU.u_wallace._0823_ ),
    .B1(\u_cpu.ALU.u_wallace._0812_ ),
    .B2(\u_cpu.ALU.u_wallace._0819_ ),
    .Y(\u_cpu.ALU.u_wallace._0868_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._6634_  (.A1(\u_cpu.ALU.u_wallace._0451_ ),
    .A2(\u_cpu.ALU.u_wallace._0644_ ),
    .A3(\u_cpu.ALU.u_wallace._0637_ ),
    .B1(\u_cpu.ALU.u_wallace._0656_ ),
    .B2(\u_cpu.ALU.u_wallace._0650_ ),
    .X(\u_cpu.ALU.u_wallace._0869_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6635_  (.A1(\u_cpu.ALU.u_wallace._0867_ ),
    .A2(\u_cpu.ALU.u_wallace._0868_ ),
    .B1(\u_cpu.ALU.u_wallace._0869_ ),
    .Y(\u_cpu.ALU.u_wallace._0870_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6636_  (.A1(\u_cpu.ALU.u_wallace._0865_ ),
    .A2(\u_cpu.ALU.u_wallace._0866_ ),
    .B1(\u_cpu.ALU.u_wallace._0835_ ),
    .B2(\u_cpu.ALU.u_wallace._0870_ ),
    .Y(\u_cpu.ALU.u_wallace._0871_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._6637_  (.A1(\u_cpu.ALU.u_wallace._0835_ ),
    .A2(\u_cpu.ALU.u_wallace._0860_ ),
    .B1(\u_cpu.ALU.u_wallace._0666_ ),
    .B2(\u_cpu.ALU.u_wallace._0863_ ),
    .C1(\u_cpu.ALU.u_wallace._0871_ ),
    .X(\u_cpu.ALU.u_wallace._0872_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6638_  (.A1(\u_cpu.ALU.u_wallace._0459_ ),
    .A2(\u_cpu.ALU.u_wallace._0609_ ),
    .B1(\u_cpu.ALU.u_wallace._0613_ ),
    .C1(\u_cpu.ALU.u_wallace._0616_ ),
    .X(\u_cpu.ALU.u_wallace._0874_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6639_  (.A(\u_cpu.ALU.u_wallace._0613_ ),
    .B(\u_cpu.ALU.u_wallace._0616_ ),
    .Y(\u_cpu.ALU.u_wallace._0875_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._6640_  (.A1(\u_cpu.ALU.u_wallace._4678_ ),
    .A2(\u_cpu.ALU.u_wallace._0458_ ),
    .A3(\u_cpu.ALU.u_wallace._0440_ ),
    .B1(\u_cpu.ALU.u_wallace._0454_ ),
    .X(\u_cpu.ALU.u_wallace._0876_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._6641_  (.A1(\u_cpu.ALU.u_wallace._0875_ ),
    .A2(\u_cpu.ALU.u_wallace._0876_ ),
    .B1_N(\u_cpu.ALU.u_wallace._0623_ ),
    .Y(\u_cpu.ALU.u_wallace._0877_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6642_  (.A(\u_cpu.ALU.u_wallace._4561_ ),
    .B(\u_cpu.ALU.u_wallace._0041_ ),
    .Y(\u_cpu.ALU.u_wallace._0878_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._6643_  (.A1(\u_cpu.ALU.u_wallace._4717_ ),
    .A2(\u_cpu.ALU.u_wallace._4783_ ),
    .A3(\u_cpu.ALU.u_wallace._4599_ ),
    .A4(\u_cpu.ALU.u_wallace._4554_ ),
    .B1(\u_cpu.ALU.u_wallace._0878_ ),
    .X(\u_cpu.ALU.u_wallace._0879_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6644_  (.A1(\u_cpu.ALU.u_wallace._4401_ ),
    .A2(\u_cpu.ALU.SrcB[9] ),
    .B1(\u_cpu.ALU.u_wallace._4550_ ),
    .B2(\u_cpu.ALU.SrcB[8] ),
    .Y(\u_cpu.ALU.u_wallace._0880_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6645_  (.A(\u_cpu.ALU.u_wallace._3821_ ),
    .B(\u_cpu.ALU.u_wallace._4609_ ),
    .Y(\u_cpu.ALU.u_wallace._0881_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6646_  (.A1(\u_cpu.ALU.u_wallace._0881_ ),
    .A2(\u_cpu.ALU.u_wallace._0685_ ),
    .B1(\u_cpu.ALU.u_wallace._0683_ ),
    .Y(\u_cpu.ALU.u_wallace._0882_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6647_  (.A(\u_cpu.ALU.u_wallace._4847_ ),
    .B(\u_cpu.ALU.u_wallace._4562_ ),
    .C(\u_cpu.ALU.u_wallace._4598_ ),
    .D(\u_cpu.ALU.u_wallace._4557_ ),
    .X(\u_cpu.ALU.u_wallace._0883_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6648_  (.A1(\u_cpu.ALU.u_wallace._4677_ ),
    .A2(\u_cpu.ALU.u_wallace._4602_ ),
    .B1(\u_cpu.ALU.u_wallace._0880_ ),
    .B2(\u_cpu.ALU.u_wallace._0883_ ),
    .Y(\u_cpu.ALU.u_wallace._0885_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6649_  (.A1(\u_cpu.ALU.u_wallace._0879_ ),
    .A2(\u_cpu.ALU.u_wallace._0880_ ),
    .B1(\u_cpu.ALU.u_wallace._0882_ ),
    .C1(\u_cpu.ALU.u_wallace._0885_ ),
    .X(\u_cpu.ALU.u_wallace._0886_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6650_  (.A1(\u_cpu.ALU.u_wallace._4450_ ),
    .A2(\u_cpu.ALU.u_wallace._4731_ ),
    .B1(\u_cpu.ALU.u_wallace._0144_ ),
    .B2(\u_cpu.ALU.u_wallace._3777_ ),
    .X(\u_cpu.ALU.u_wallace._0887_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6651_  (.A(\u_cpu.ALU.u_wallace._3821_ ),
    .B(\u_cpu.ALU.u_wallace._3832_ ),
    .C(\u_cpu.ALU.u_wallace._4837_ ),
    .D(\u_cpu.ALU.u_wallace._0029_ ),
    .Y(\u_cpu.ALU.u_wallace._0888_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6652_  (.A(\u_cpu.ALU.u_wallace._1322_ ),
    .B(\u_cpu.ALU.u_wallace._0033_ ),
    .Y(\u_cpu.ALU.u_wallace._0889_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6653_  (.A1(\u_cpu.ALU.u_wallace._0887_ ),
    .A2(\u_cpu.ALU.u_wallace._0888_ ),
    .B1(\u_cpu.ALU.u_wallace._0889_ ),
    .X(\u_cpu.ALU.u_wallace._0890_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6654_  (.A1(\u_cpu.ALU.u_wallace._4813_ ),
    .A2(\u_cpu.ALU.u_wallace._0036_ ),
    .B1(\u_cpu.ALU.u_wallace._0887_ ),
    .C1(\u_cpu.ALU.u_wallace._0888_ ),
    .Y(\u_cpu.ALU.u_wallace._0891_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6655_  (.A(\u_cpu.ALU.u_wallace._0890_ ),
    .B(\u_cpu.ALU.u_wallace._0891_ ),
    .Y(\u_cpu.ALU.u_wallace._0892_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._6656_  (.A(\u_cpu.ALU.u_wallace._0878_ ),
    .B(\u_cpu.ALU.u_wallace._0880_ ),
    .C(\u_cpu.ALU.u_wallace._0883_ ),
    .Y(\u_cpu.ALU.u_wallace._0893_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._6657_  (.A1(\u_cpu.ALU.u_wallace._4677_ ),
    .A2(\u_cpu.ALU.u_wallace._4602_ ),
    .B1(\u_cpu.ALU.u_wallace._0880_ ),
    .B2(\u_cpu.ALU.u_wallace._0883_ ),
    .X(\u_cpu.ALU.u_wallace._0894_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._6658_  (.A1(\u_cpu.ALU.u_wallace._0893_ ),
    .A2(\u_cpu.ALU.u_wallace._0894_ ),
    .B1_N(\u_cpu.ALU.u_wallace._0882_ ),
    .Y(\u_cpu.ALU.u_wallace._0896_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6659_  (.A(\u_cpu.ALU.u_wallace._0892_ ),
    .B(\u_cpu.ALU.u_wallace._0896_ ),
    .Y(\u_cpu.ALU.u_wallace._0897_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6660_  (.A(\u_cpu.ALU.u_wallace._4847_ ),
    .B(\u_cpu.ALU.u_wallace._4562_ ),
    .C(\u_cpu.ALU.u_wallace._0045_ ),
    .D(\u_cpu.ALU.u_wallace._4557_ ),
    .Y(\u_cpu.ALU.u_wallace._0898_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._6661_  (.A_N(\u_cpu.ALU.u_wallace._0880_ ),
    .B(\u_cpu.ALU.u_wallace._0898_ ),
    .C(\u_cpu.ALU.u_wallace._4669_ ),
    .D(\u_cpu.ALU.u_wallace._0052_ ),
    .Y(\u_cpu.ALU.u_wallace._0899_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6662_  (.A1(\u_cpu.ALU.u_wallace._0899_ ),
    .A2(\u_cpu.ALU.u_wallace._0885_ ),
    .B1(\u_cpu.ALU.u_wallace._0882_ ),
    .Y(\u_cpu.ALU.u_wallace._0900_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6663_  (.A1(\u_cpu.ALU.u_wallace._0886_ ),
    .A2(\u_cpu.ALU.u_wallace._0900_ ),
    .B1(\u_cpu.ALU.u_wallace._0890_ ),
    .C1(\u_cpu.ALU.u_wallace._0891_ ),
    .Y(\u_cpu.ALU.u_wallace._0901_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._6664_  (.A1(\u_cpu.ALU.u_wallace._0874_ ),
    .A2(\u_cpu.ALU.u_wallace._0877_ ),
    .B1(\u_cpu.ALU.u_wallace._0886_ ),
    .B2(\u_cpu.ALU.u_wallace._0897_ ),
    .C1(\u_cpu.ALU.u_wallace._0901_ ),
    .Y(\u_cpu.ALU.u_wallace._0902_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6665_  (.A1(\u_cpu.ALU.u_wallace._0613_ ),
    .A2(\u_cpu.ALU.u_wallace._0622_ ),
    .B1(\u_cpu.ALU.u_wallace._0619_ ),
    .B2(\u_cpu.ALU.u_wallace._0623_ ),
    .Y(\u_cpu.ALU.u_wallace._0903_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6666_  (.A1(\u_cpu.ALU.u_wallace._0886_ ),
    .A2(\u_cpu.ALU.u_wallace._0900_ ),
    .B1(\u_cpu.ALU.u_wallace._0892_ ),
    .Y(\u_cpu.ALU.u_wallace._0904_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6667_  (.A1(\u_cpu.ALU.u_wallace._0879_ ),
    .A2(\u_cpu.ALU.u_wallace._0880_ ),
    .B1(\u_cpu.ALU.u_wallace._0882_ ),
    .C1(\u_cpu.ALU.u_wallace._0885_ ),
    .Y(\u_cpu.ALU.u_wallace._0905_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._6668_  (.A_N(\u_cpu.ALU.u_wallace._0892_ ),
    .B(\u_cpu.ALU.u_wallace._0905_ ),
    .C(\u_cpu.ALU.u_wallace._0896_ ),
    .Y(\u_cpu.ALU.u_wallace._0907_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6669_  (.A(\u_cpu.ALU.u_wallace._0903_ ),
    .B(\u_cpu.ALU.u_wallace._0904_ ),
    .C(\u_cpu.ALU.u_wallace._0907_ ),
    .Y(\u_cpu.ALU.u_wallace._0908_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._6670_  (.A1(\u_cpu.ALU.u_wallace._0681_ ),
    .A2(\u_cpu.ALU.u_wallace._0684_ ),
    .A3(\u_cpu.ALU.u_wallace._0688_ ),
    .B1(\u_cpu.ALU.u_wallace._0708_ ),
    .X(\u_cpu.ALU.u_wallace._0909_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6671_  (.A1(\u_cpu.ALU.u_wallace._0902_ ),
    .A2(\u_cpu.ALU.u_wallace._0908_ ),
    .B1(\u_cpu.ALU.u_wallace._0909_ ),
    .Y(\u_cpu.ALU.u_wallace._0910_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6672_  (.A(\u_cpu.ALU.u_wallace._0902_ ),
    .B(\u_cpu.ALU.u_wallace._0908_ ),
    .C(\u_cpu.ALU.u_wallace._0909_ ),
    .X(\u_cpu.ALU.u_wallace._0911_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6673_  (.A(\u_cpu.ALU.u_wallace._0869_ ),
    .B(\u_cpu.ALU.u_wallace._0867_ ),
    .C(\u_cpu.ALU.u_wallace._0868_ ),
    .Y(\u_cpu.ALU.u_wallace._0912_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6674_  (.A1(\u_cpu.ALU.u_wallace._0854_ ),
    .A2(\u_cpu.ALU.u_wallace._0849_ ),
    .B1(\u_cpu.ALU.u_wallace._0857_ ),
    .Y(\u_cpu.ALU.u_wallace._0913_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6675_  (.A1(\u_cpu.ALU.u_wallace._0912_ ),
    .A2(\u_cpu.ALU.u_wallace._0859_ ),
    .B1(\u_cpu.ALU.u_wallace._0913_ ),
    .X(\u_cpu.ALU.u_wallace._0914_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6676_  (.A1(\u_cpu.ALU.u_wallace._0865_ ),
    .A2(\u_cpu.ALU.u_wallace._0866_ ),
    .B1(\u_cpu.ALU.u_wallace._0912_ ),
    .C1(\u_cpu.ALU.u_wallace._0859_ ),
    .Y(\u_cpu.ALU.u_wallace._0915_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6677_  (.A1(\u_cpu.ALU.u_wallace._0874_ ),
    .A2(\u_cpu.ALU.u_wallace._0624_ ),
    .B1(\u_cpu.ALU.u_wallace._0623_ ),
    .Y(\u_cpu.ALU.u_wallace._0916_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.ALU.u_wallace._6678_  (.A1(\u_cpu.ALU.u_wallace._0874_ ),
    .A2(\u_cpu.ALU.u_wallace._0624_ ),
    .A3(\u_cpu.ALU.u_wallace._0877_ ),
    .B1(\u_cpu.ALU.u_wallace._0916_ ),
    .Y(\u_cpu.ALU.u_wallace._0918_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6679_  (.A1(\u_cpu.ALU.u_wallace._0918_ ),
    .A2(\u_cpu.ALU.u_wallace._0659_ ),
    .B1(\u_cpu.ALU.u_wallace._0666_ ),
    .Y(\u_cpu.ALU.u_wallace._0919_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6680_  (.A(\u_cpu.ALU.u_wallace._0914_ ),
    .B(\u_cpu.ALU.u_wallace._0915_ ),
    .C(\u_cpu.ALU.u_wallace._0919_ ),
    .Y(\u_cpu.ALU.u_wallace._0920_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6681_  (.A1(\u_cpu.ALU.u_wallace._0910_ ),
    .A2(\u_cpu.ALU.u_wallace._0911_ ),
    .B1(\u_cpu.ALU.u_wallace._0920_ ),
    .Y(\u_cpu.ALU.u_wallace._0921_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._6682_  (.A1(\u_cpu.ALU.u_wallace._0835_ ),
    .A2(\u_cpu.ALU.u_wallace._0860_ ),
    .B1(\u_cpu.ALU.u_wallace._0666_ ),
    .B2(\u_cpu.ALU.u_wallace._0863_ ),
    .C1(\u_cpu.ALU.u_wallace._0871_ ),
    .Y(\u_cpu.ALU.u_wallace._0922_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6683_  (.A1(\u_cpu.ALU.u_wallace._0694_ ),
    .A2(\u_cpu.ALU.u_wallace._0693_ ),
    .B1(\u_cpu.ALU.u_wallace._0707_ ),
    .X(\u_cpu.ALU.u_wallace._0923_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6684_  (.A(\u_cpu.ALU.u_wallace._0923_ ),
    .B(\u_cpu.ALU.u_wallace._0902_ ),
    .C(\u_cpu.ALU.u_wallace._0908_ ),
    .X(\u_cpu.ALU.u_wallace._0924_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6685_  (.A1(\u_cpu.ALU.u_wallace._0902_ ),
    .A2(\u_cpu.ALU.u_wallace._0908_ ),
    .B1(\u_cpu.ALU.u_wallace._0923_ ),
    .Y(\u_cpu.ALU.u_wallace._0925_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6686_  (.A1_N(\u_cpu.ALU.u_wallace._0922_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0920_ ),
    .B1(\u_cpu.ALU.u_wallace._0924_ ),
    .B2(\u_cpu.ALU.u_wallace._0925_ ),
    .Y(\u_cpu.ALU.u_wallace._0926_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6687_  (.A(\u_cpu.ALU.u_wallace._0713_ ),
    .B(\u_cpu.ALU.u_wallace._0712_ ),
    .Y(\u_cpu.ALU.u_wallace._0927_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6688_  (.A1(\u_cpu.ALU.u_wallace._0872_ ),
    .A2(\u_cpu.ALU.u_wallace._0921_ ),
    .B1(\u_cpu.ALU.u_wallace._0926_ ),
    .C1(\u_cpu.ALU.u_wallace._0927_ ),
    .X(\u_cpu.ALU.u_wallace._0929_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6689_  (.A1_N(\u_cpu.ALU.u_wallace._0705_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0704_ ),
    .B1(\u_cpu.ALU.u_wallace._0702_ ),
    .B2(\u_cpu.ALU.u_wallace._0695_ ),
    .Y(\u_cpu.ALU.u_wallace._0930_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._6690_  (.A1(\u_cpu.ALU.u_wallace._0729_ ),
    .A2(\u_cpu.ALU.u_wallace._0551_ ),
    .A3(\u_cpu.ALU.u_wallace._0162_ ),
    .B1(\u_cpu.ALU.u_wallace._0737_ ),
    .Y(\u_cpu.ALU.u_wallace._0931_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6691_  (.A(\u_cpu.ALU.u_wallace._1848_ ),
    .B(\u_cpu.ALU.u_wallace._4529_ ),
    .C(\u_cpu.ALU.u_wallace._4840_ ),
    .D(\u_cpu.ALU.u_wallace._4838_ ),
    .X(\u_cpu.ALU.u_wallace._0932_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6692_  (.A(\u_cpu.ALU.u_wallace._1979_ ),
    .B(\u_cpu.ALU.u_wallace._0365_ ),
    .Y(\u_cpu.ALU.u_wallace._0933_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6693_  (.A(\u_cpu.ALU.u_wallace._1793_ ),
    .B(\u_cpu.ALU.u_wallace._4731_ ),
    .Y(\u_cpu.ALU.u_wallace._0934_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6694_  (.A(\u_cpu.ALU.u_wallace._1180_ ),
    .B(\u_cpu.ALU.u_wallace._0033_ ),
    .Y(\u_cpu.ALU.u_wallace._0935_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6695_  (.A1(\u_cpu.ALU.u_wallace._0933_ ),
    .A2(\u_cpu.ALU.u_wallace._0934_ ),
    .B1(\u_cpu.ALU.u_wallace._0935_ ),
    .Y(\u_cpu.ALU.u_wallace._0936_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6696_  (.A1(\u_cpu.ALU.u_wallace._2922_ ),
    .A2(\u_cpu.ALU.u_wallace._0730_ ),
    .B1(\u_cpu.ALU.u_wallace._0732_ ),
    .B2(\u_cpu.ALU.u_wallace._0600_ ),
    .X(\u_cpu.ALU.u_wallace._0937_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6697_  (.A(\u_cpu.ALU.u_wallace._1180_ ),
    .B(\u_cpu.ALU.u_wallace._1191_ ),
    .C(\u_cpu.ALU.u_wallace._0546_ ),
    .D(\u_cpu.ALU.u_wallace._0547_ ),
    .Y(\u_cpu.ALU.u_wallace._0938_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6698_  (.A(\u_cpu.ALU.u_wallace._0937_ ),
    .B(\u_cpu.ALU.u_wallace._0938_ ),
    .C(\u_cpu.ALU.u_wallace._4597_ ),
    .D(\u_cpu.ALU.u_wallace._0735_ ),
    .Y(\u_cpu.ALU.u_wallace._0940_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6699_  (.A(\u_cpu.ALU.u_wallace._0553_ ),
    .X(\u_cpu.ALU.u_wallace._0941_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6700_  (.A1(\u_cpu.ALU.u_wallace._1180_ ),
    .A2(\u_cpu.ALU.u_wallace._0546_ ),
    .B1(\u_cpu.ALU.u_wallace._0547_ ),
    .B2(\u_cpu.ALU.u_wallace._1191_ ),
    .Y(\u_cpu.ALU.u_wallace._0942_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6701_  (.A(\u_cpu.ALU.u_wallace._4556_ ),
    .B(\u_cpu.ALU.u_wallace._2549_ ),
    .C(\u_cpu.ALU.u_wallace._0120_ ),
    .D(\u_cpu.ALU.u_wallace._0728_ ),
    .X(\u_cpu.ALU.u_wallace._0943_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6702_  (.A1(\u_cpu.ALU.u_wallace._0403_ ),
    .A2(\u_cpu.ALU.u_wallace._0941_ ),
    .B1(\u_cpu.ALU.u_wallace._0942_ ),
    .B2(\u_cpu.ALU.u_wallace._0943_ ),
    .Y(\u_cpu.ALU.u_wallace._0944_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6703_  (.A1(\u_cpu.ALU.u_wallace._0932_ ),
    .A2(\u_cpu.ALU.u_wallace._0936_ ),
    .B1(\u_cpu.ALU.u_wallace._0940_ ),
    .C1(\u_cpu.ALU.u_wallace._0944_ ),
    .Y(\u_cpu.ALU.u_wallace._0945_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6704_  (.A1(\u_cpu.ALU.u_wallace._0933_ ),
    .A2(\u_cpu.ALU.u_wallace._0934_ ),
    .B1(\u_cpu.ALU.u_wallace._0935_ ),
    .X(\u_cpu.ALU.u_wallace._0946_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6705_  (.A1(\u_cpu.ALU.u_wallace._0933_ ),
    .A2(\u_cpu.ALU.u_wallace._0934_ ),
    .B1(\u_cpu.ALU.u_wallace._0946_ ),
    .Y(\u_cpu.ALU.u_wallace._0947_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6706_  (.A1(\u_cpu.ALU.u_wallace._0940_ ),
    .A2(\u_cpu.ALU.u_wallace._0944_ ),
    .B1(\u_cpu.ALU.u_wallace._0947_ ),
    .X(\u_cpu.ALU.u_wallace._0948_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._6707_  (.A_N(\u_cpu.ALU.u_wallace._0931_ ),
    .B(\u_cpu.ALU.u_wallace._0945_ ),
    .C(\u_cpu.ALU.u_wallace._0948_ ),
    .Y(\u_cpu.ALU.u_wallace._0949_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6708_  (.A1(\u_cpu.ALU.u_wallace._0932_ ),
    .A2(\u_cpu.ALU.u_wallace._0936_ ),
    .B1(\u_cpu.ALU.u_wallace._0940_ ),
    .C1(\u_cpu.ALU.u_wallace._0944_ ),
    .X(\u_cpu.ALU.u_wallace._0951_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6709_  (.A1(\u_cpu.ALU.u_wallace._0940_ ),
    .A2(\u_cpu.ALU.u_wallace._0944_ ),
    .B1(\u_cpu.ALU.u_wallace._0947_ ),
    .Y(\u_cpu.ALU.u_wallace._0952_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6710_  (.A1(\u_cpu.ALU.u_wallace._0951_ ),
    .A2(\u_cpu.ALU.u_wallace._0952_ ),
    .B1(\u_cpu.ALU.u_wallace._0931_ ),
    .Y(\u_cpu.ALU.u_wallace._0953_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._6711_  (.A1(\u_cpu.ALU.u_wallace._0558_ ),
    .A2(\u_cpu.ALU.u_wallace._0555_ ),
    .B1(\u_cpu.ALU.u_wallace._0552_ ),
    .X(\u_cpu.ALU.u_wallace._0954_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._6712_  (.A1(\u_cpu.ALU.u_wallace._0954_ ),
    .A2(\u_cpu.ALU.u_wallace._0745_ ),
    .B1_N(\u_cpu.ALU.u_wallace._0739_ ),
    .Y(\u_cpu.ALU.u_wallace._0955_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6713_  (.A1(\u_cpu.ALU.u_wallace._0949_ ),
    .A2(\u_cpu.ALU.u_wallace._0953_ ),
    .B1(\u_cpu.ALU.u_wallace._0955_ ),
    .X(\u_cpu.ALU.u_wallace._0956_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6714_  (.A(\u_cpu.ALU.SrcB[18] ),
    .X(\u_cpu.ALU.u_wallace._0957_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6715_  (.A(\u_cpu.ALU.u_wallace._0957_ ),
    .X(\u_cpu.ALU.u_wallace._0958_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6716_  (.A(\u_cpu.ALU.u_wallace._0958_ ),
    .X(\u_cpu.ALU.u_wallace._0959_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6717_  (.A(\u_cpu.ALU.u_wallace._0734_ ),
    .B(\u_cpu.ALU.u_wallace._0738_ ),
    .Y(\u_cpu.ALU.u_wallace._0960_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._6718_  (.A1(\u_cpu.ALU.u_wallace._0621_ ),
    .A2(\u_cpu.ALU.u_wallace._0124_ ),
    .A3(\u_cpu.ALU.u_wallace._0725_ ),
    .B1(\u_cpu.ALU.u_wallace._0496_ ),
    .X(\u_cpu.ALU.u_wallace._0962_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6719_  (.A1(\u_cpu.ALU.u_wallace._0960_ ),
    .A2(\u_cpu.ALU.u_wallace._0962_ ),
    .B1(\u_cpu.ALU.u_wallace._0954_ ),
    .Y(\u_cpu.ALU.u_wallace._0963_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6720_  (.A1(\u_cpu.ALU.u_wallace._0739_ ),
    .A2(\u_cpu.ALU.u_wallace._0963_ ),
    .B1(\u_cpu.ALU.u_wallace._0949_ ),
    .C1(\u_cpu.ALU.u_wallace._0953_ ),
    .Y(\u_cpu.ALU.u_wallace._0964_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6721_  (.A(\u_cpu.ALU.u_wallace._0956_ ),
    .B(\u_cpu.ALU.u_wallace._0959_ ),
    .C(\u_cpu.ALU.u_wallace._0129_ ),
    .D(\u_cpu.ALU.u_wallace._0964_ ),
    .Y(\u_cpu.ALU.u_wallace._0965_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6722_  (.A1(\u_cpu.ALU.u_wallace._0739_ ),
    .A2(\u_cpu.ALU.u_wallace._0963_ ),
    .B1(\u_cpu.ALU.u_wallace._0949_ ),
    .C1(\u_cpu.ALU.u_wallace._0953_ ),
    .X(\u_cpu.ALU.u_wallace._0966_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6723_  (.A1(\u_cpu.ALU.u_wallace._0949_ ),
    .A2(\u_cpu.ALU.u_wallace._0953_ ),
    .B1(\u_cpu.ALU.u_wallace._0955_ ),
    .Y(\u_cpu.ALU.u_wallace._0967_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6724_  (.A(\u_cpu.ALU.u_wallace._0129_ ),
    .B(\u_cpu.ALU.u_wallace._0959_ ),
    .Y(\u_cpu.ALU.u_wallace._0968_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6725_  (.A1(\u_cpu.ALU.u_wallace._0966_ ),
    .A2(\u_cpu.ALU.u_wallace._0967_ ),
    .B1(\u_cpu.ALU.u_wallace._0968_ ),
    .Y(\u_cpu.ALU.u_wallace._0969_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6726_  (.A(\u_cpu.ALU.u_wallace._0930_ ),
    .B(\u_cpu.ALU.u_wallace._0965_ ),
    .C(\u_cpu.ALU.u_wallace._0969_ ),
    .Y(\u_cpu.ALU.u_wallace._0970_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._6727_  (.A1(\u_cpu.ALU.u_wallace._0966_ ),
    .A2(\u_cpu.ALU.u_wallace._0967_ ),
    .B1_N(\u_cpu.ALU.u_wallace._0968_ ),
    .Y(\u_cpu.ALU.u_wallace._0971_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._6728_  (.A(\u_cpu.ALU.u_wallace._0959_ ),
    .Y(\u_cpu.ALU.u_wallace._0973_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6729_  (.A1(\u_cpu.ALU.u_wallace._0043_ ),
    .A2(\u_cpu.ALU.u_wallace._0973_ ),
    .B1(\u_cpu.ALU.u_wallace._0964_ ),
    .C1(\u_cpu.ALU.u_wallace._0956_ ),
    .Y(\u_cpu.ALU.u_wallace._0974_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._6730_  (.A1_N(\u_cpu.ALU.u_wallace._0702_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0695_ ),
    .B1(\u_cpu.ALU.u_wallace._0705_ ),
    .B2(\u_cpu.ALU.u_wallace._0704_ ),
    .Y(\u_cpu.ALU.u_wallace._0975_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6731_  (.A(\u_cpu.ALU.u_wallace._0971_ ),
    .B(\u_cpu.ALU.u_wallace._0974_ ),
    .C(\u_cpu.ALU.u_wallace._0975_ ),
    .Y(\u_cpu.ALU.u_wallace._0976_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6732_  (.A1(\u_cpu.ALU.u_wallace._0970_ ),
    .A2(\u_cpu.ALU.u_wallace._0976_ ),
    .B1(\u_cpu.ALU.u_wallace._0751_ ),
    .Y(\u_cpu.ALU.u_wallace._0977_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6733_  (.A(\u_cpu.ALU.u_wallace._0751_ ),
    .B(\u_cpu.ALU.u_wallace._0970_ ),
    .C(\u_cpu.ALU.u_wallace._0976_ ),
    .X(\u_cpu.ALU.u_wallace._0978_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6734_  (.A1(\u_cpu.ALU.u_wallace._0910_ ),
    .A2(\u_cpu.ALU.u_wallace._0911_ ),
    .B1(\u_cpu.ALU.u_wallace._0922_ ),
    .C1(\u_cpu.ALU.u_wallace._0920_ ),
    .X(\u_cpu.ALU.u_wallace._0979_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._6735_  (.A1(\u_cpu.ALU.u_wallace._0903_ ),
    .A2(\u_cpu.ALU.u_wallace._0904_ ),
    .A3(\u_cpu.ALU.u_wallace._0907_ ),
    .B1(\u_cpu.ALU.u_wallace._0909_ ),
    .Y(\u_cpu.ALU.u_wallace._0980_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6736_  (.A1(\u_cpu.ALU.u_wallace._0902_ ),
    .A2(\u_cpu.ALU.u_wallace._0980_ ),
    .B1(\u_cpu.ALU.u_wallace._0925_ ),
    .Y(\u_cpu.ALU.u_wallace._0981_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6737_  (.A1(\u_cpu.ALU.u_wallace._0922_ ),
    .A2(\u_cpu.ALU.u_wallace._0920_ ),
    .B1(\u_cpu.ALU.u_wallace._0981_ ),
    .Y(\u_cpu.ALU.u_wallace._0982_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._6738_  (.A1(\u_cpu.ALU.u_wallace._0680_ ),
    .A2(\u_cpu.ALU.u_wallace._0706_ ),
    .A3(\u_cpu.ALU.u_wallace._0711_ ),
    .B1(\u_cpu.ALU.u_wallace._0673_ ),
    .Y(\u_cpu.ALU.u_wallace._0984_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6739_  (.A1(\u_cpu.ALU.u_wallace._0979_ ),
    .A2(\u_cpu.ALU.u_wallace._0982_ ),
    .B1(\u_cpu.ALU.u_wallace._0984_ ),
    .Y(\u_cpu.ALU.u_wallace._0985_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6740_  (.A1(\u_cpu.ALU.u_wallace._0977_ ),
    .A2(\u_cpu.ALU.u_wallace._0978_ ),
    .B1(\u_cpu.ALU.u_wallace._0985_ ),
    .Y(\u_cpu.ALU.u_wallace._0986_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6741_  (.A1(\u_cpu.ALU.u_wallace._0872_ ),
    .A2(\u_cpu.ALU.u_wallace._0921_ ),
    .B1(\u_cpu.ALU.u_wallace._0926_ ),
    .C1(\u_cpu.ALU.u_wallace._0927_ ),
    .Y(\u_cpu.ALU.u_wallace._0987_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6742_  (.A(\u_cpu.ALU.u_wallace._0970_ ),
    .B(\u_cpu.ALU.u_wallace._0976_ ),
    .C(\u_cpu.ALU.u_wallace._0755_ ),
    .X(\u_cpu.ALU.u_wallace._0988_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6743_  (.A1(\u_cpu.ALU.u_wallace._0970_ ),
    .A2(\u_cpu.ALU.u_wallace._0976_ ),
    .B1(\u_cpu.ALU.u_wallace._0755_ ),
    .Y(\u_cpu.ALU.u_wallace._0989_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6744_  (.A1_N(\u_cpu.ALU.u_wallace._0987_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0985_ ),
    .B1(\u_cpu.ALU.u_wallace._0988_ ),
    .B2(\u_cpu.ALU.u_wallace._0989_ ),
    .Y(\u_cpu.ALU.u_wallace._0990_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._6745_  (.A1(\u_cpu.ALU.u_wallace._0776_ ),
    .A2(\u_cpu.ALU.u_wallace._0761_ ),
    .B1(\u_cpu.ALU.u_wallace._0929_ ),
    .B2(\u_cpu.ALU.u_wallace._0986_ ),
    .C1(\u_cpu.ALU.u_wallace._0990_ ),
    .Y(\u_cpu.ALU.u_wallace._0991_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6746_  (.A1(\u_cpu.ALU.u_wallace._0872_ ),
    .A2(\u_cpu.ALU.u_wallace._0921_ ),
    .B1(\u_cpu.ALU.u_wallace._0926_ ),
    .Y(\u_cpu.ALU.u_wallace._0992_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6747_  (.A1(\u_cpu.ALU.u_wallace._0970_ ),
    .A2(\u_cpu.ALU.u_wallace._0976_ ),
    .B1(\u_cpu.ALU.u_wallace._0751_ ),
    .X(\u_cpu.ALU.u_wallace._0993_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6748_  (.A(\u_cpu.ALU.u_wallace._0751_ ),
    .B(\u_cpu.ALU.u_wallace._0970_ ),
    .C(\u_cpu.ALU.u_wallace._0976_ ),
    .Y(\u_cpu.ALU.u_wallace._0995_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6749_  (.A1(\u_cpu.ALU.u_wallace._0993_ ),
    .A2(\u_cpu.ALU.u_wallace._0995_ ),
    .B1(\u_cpu.ALU.u_wallace._0984_ ),
    .B2(\u_cpu.ALU.u_wallace._0992_ ),
    .Y(\u_cpu.ALU.u_wallace._0996_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6750_  (.A1(\u_cpu.ALU.u_wallace._0984_ ),
    .A2(\u_cpu.ALU.u_wallace._0992_ ),
    .B1(\u_cpu.ALU.u_wallace._0996_ ),
    .Y(\u_cpu.ALU.u_wallace._0997_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6751_  (.A1(\u_cpu.ALU.u_wallace._0760_ ),
    .A2(\u_cpu.ALU.u_wallace._0777_ ),
    .B1(\u_cpu.ALU.u_wallace._0718_ ),
    .Y(\u_cpu.ALU.u_wallace._0998_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6752_  (.A1(\u_cpu.ALU.u_wallace._0997_ ),
    .A2(\u_cpu.ALU.u_wallace._0990_ ),
    .B1(\u_cpu.ALU.u_wallace._0998_ ),
    .X(\u_cpu.ALU.u_wallace._0999_ ));
 sky130_fd_sc_hd__and4bb_2 \u_cpu.ALU.u_wallace._6753_  (.A_N(\u_cpu.ALU.u_wallace._0565_ ),
    .B_N(\u_cpu.ALU.u_wallace._0287_ ),
    .C(\u_cpu.ALU.u_wallace._0748_ ),
    .D(\u_cpu.ALU.u_wallace._0756_ ),
    .X(\u_cpu.ALU.u_wallace._1000_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._6754_  (.A(\u_cpu.ALU.u_wallace._1000_ ),
    .Y(\u_cpu.ALU.u_wallace._1001_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6755_  (.A(\u_cpu.ALU.u_wallace._0752_ ),
    .B(\u_cpu.ALU.u_wallace._1001_ ),
    .Y(\u_cpu.ALU.u_wallace._1002_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6756_  (.A(\u_cpu.ALU.u_wallace._0991_ ),
    .B(\u_cpu.ALU.u_wallace._0999_ ),
    .C(\u_cpu.ALU.u_wallace._1002_ ),
    .Y(\u_cpu.ALU.u_wallace._1003_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._6757_  (.A1(\u_cpu.ALU.u_wallace._0776_ ),
    .A2(\u_cpu.ALU.u_wallace._0761_ ),
    .B1(\u_cpu.ALU.u_wallace._0929_ ),
    .B2(\u_cpu.ALU.u_wallace._0986_ ),
    .C1(\u_cpu.ALU.u_wallace._0990_ ),
    .X(\u_cpu.ALU.u_wallace._1004_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6758_  (.A1(\u_cpu.ALU.u_wallace._0997_ ),
    .A2(\u_cpu.ALU.u_wallace._0990_ ),
    .B1(\u_cpu.ALU.u_wallace._0998_ ),
    .Y(\u_cpu.ALU.u_wallace._1006_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._6759_  (.A(\u_cpu.ALU.u_wallace._1002_ ),
    .Y(\u_cpu.ALU.u_wallace._1007_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6760_  (.A1(\u_cpu.ALU.u_wallace._1004_ ),
    .A2(\u_cpu.ALU.u_wallace._1006_ ),
    .B1(\u_cpu.ALU.u_wallace._1007_ ),
    .Y(\u_cpu.ALU.u_wallace._1008_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6761_  (.A(\u_cpu.ALU.u_wallace._0799_ ),
    .B(\u_cpu.ALU.u_wallace._1003_ ),
    .C(\u_cpu.ALU.u_wallace._1008_ ),
    .Y(\u_cpu.ALU.u_wallace._1009_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6762_  (.A1(\u_cpu.ALU.u_wallace._1003_ ),
    .A2(\u_cpu.ALU.u_wallace._1008_ ),
    .B1(\u_cpu.ALU.u_wallace._0799_ ),
    .X(\u_cpu.ALU.u_wallace._1010_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6763_  (.A(\u_cpu.ALU.u_wallace._0787_ ),
    .B(\u_cpu.ALU.u_wallace._0798_ ),
    .C(\u_cpu.ALU.u_wallace._1009_ ),
    .D(\u_cpu.ALU.u_wallace._1010_ ),
    .Y(\u_cpu.ALU.u_wallace._1011_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6764_  (.A(\u_cpu.ALU.u_wallace._0799_ ),
    .B(\u_cpu.ALU.u_wallace._1003_ ),
    .C(\u_cpu.ALU.u_wallace._1008_ ),
    .X(\u_cpu.ALU.u_wallace._1012_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6765_  (.A1(\u_cpu.ALU.u_wallace._1003_ ),
    .A2(\u_cpu.ALU.u_wallace._1008_ ),
    .B1(\u_cpu.ALU.u_wallace._0799_ ),
    .Y(\u_cpu.ALU.u_wallace._1013_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6766_  (.A1_N(\u_cpu.ALU.u_wallace._0787_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0798_ ),
    .B1(\u_cpu.ALU.u_wallace._1012_ ),
    .B2(\u_cpu.ALU.u_wallace._1013_ ),
    .Y(\u_cpu.ALU.u_wallace._1014_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6767_  (.A(\u_cpu.ALU.u_wallace._1011_ ),
    .B(\u_cpu.ALU.u_wallace._1014_ ),
    .Y(\u_cpu.ALU.u_wallace._1015_ ));
 sky130_fd_sc_hd__nor4_2 \u_cpu.ALU.u_wallace._6768_  (.A(\u_cpu.ALU.u_wallace._0434_ ),
    .B(\u_cpu.ALU.u_wallace._0603_ ),
    .C(\u_cpu.ALU.u_wallace._0602_ ),
    .D(\u_cpu.ALU.u_wallace._0793_ ),
    .Y(\u_cpu.ALU.u_wallace._1017_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6769_  (.A1(\u_cpu.ALU.u_wallace._0795_ ),
    .A2(\u_cpu.ALU.u_wallace._0796_ ),
    .B1(\u_cpu.ALU.u_wallace._1017_ ),
    .X(\u_cpu.ALU.u_wallace._1018_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._6770_  (.A(\u_cpu.ALU.u_wallace._1015_ ),
    .B(\u_cpu.ALU.u_wallace._1018_ ),
    .X(\u_cpu.ALU.Product_Wallace[18] ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6771_  (.A1(\u_cpu.ALU.u_wallace._0752_ ),
    .A2(\u_cpu.ALU.u_wallace._1001_ ),
    .B1(\u_cpu.ALU.u_wallace._1006_ ),
    .Y(\u_cpu.ALU.u_wallace._1019_ ));
 sky130_fd_sc_hd__a32oi_2 \u_cpu.ALU.u_wallace._6772_  (.A1(\u_cpu.ALU.u_wallace._0930_ ),
    .A2(\u_cpu.ALU.u_wallace._0965_ ),
    .A3(\u_cpu.ALU.u_wallace._0969_ ),
    .B1(\u_cpu.ALU.u_wallace._0976_ ),
    .B2(\u_cpu.ALU.u_wallace._0755_ ),
    .Y(\u_cpu.ALU.u_wallace._1020_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._6773_  (.A(\u_cpu.ALU.u_wallace._1020_ ),
    .Y(\u_cpu.ALU.u_wallace._1021_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6774_  (.A(\u_cpu.ALU.u_wallace._0912_ ),
    .B(\u_cpu.ALU.u_wallace._0859_ ),
    .Y(\u_cpu.ALU.u_wallace._1022_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6775_  (.A1_N(\u_cpu.ALU.u_wallace._0913_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1022_ ),
    .B1(\u_cpu.ALU.u_wallace._0835_ ),
    .B2(\u_cpu.ALU.u_wallace._0860_ ),
    .Y(\u_cpu.ALU.u_wallace._1023_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._6776_  (.A1_N(\u_cpu.ALU.u_wallace._0910_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0911_ ),
    .B1(\u_cpu.ALU.u_wallace._0919_ ),
    .B2(\u_cpu.ALU.u_wallace._1023_ ),
    .Y(\u_cpu.ALU.u_wallace._1024_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6777_  (.A(\u_cpu.ALU.u_wallace._4007_ ),
    .B(\u_cpu.ALU.u_wallace._4291_ ),
    .C(\u_cpu.ALU.u_wallace._4550_ ),
    .D(\u_cpu.ALU.u_wallace._4650_ ),
    .Y(\u_cpu.ALU.u_wallace._1025_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6778_  (.A(\u_cpu.ALU.u_wallace._1025_ ),
    .B(\u_cpu.ALU.u_wallace._4609_ ),
    .C(\u_cpu.ALU.u_wallace._4567_ ),
    .Y(\u_cpu.ALU.u_wallace._1027_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6779_  (.A1(\u_cpu.ALU.SrcB[9] ),
    .A2(\u_cpu.ALU.u_wallace._4550_ ),
    .B1(\u_cpu.ALU.u_wallace._4646_ ),
    .B2(\u_cpu.ALU.SrcB[8] ),
    .Y(\u_cpu.ALU.u_wallace._1028_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6780_  (.A1(\u_cpu.ALU.u_wallace._0878_ ),
    .A2(\u_cpu.ALU.u_wallace._0880_ ),
    .B1(\u_cpu.ALU.u_wallace._0898_ ),
    .Y(\u_cpu.ALU.u_wallace._1029_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6781_  (.A(\u_cpu.ALU.SrcB[8] ),
    .B(\u_cpu.ALU.u_wallace._4291_ ),
    .C(\u_cpu.ALU.u_wallace._4550_ ),
    .D(\u_cpu.ALU.u_wallace._4646_ ),
    .X(\u_cpu.ALU.u_wallace._1030_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6782_  (.A1(\u_cpu.ALU.u_wallace._4573_ ),
    .A2(\u_cpu.ALU.u_wallace._4601_ ),
    .B1(\u_cpu.ALU.u_wallace._1028_ ),
    .B2(\u_cpu.ALU.u_wallace._1030_ ),
    .Y(\u_cpu.ALU.u_wallace._1031_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6783_  (.A1(\u_cpu.ALU.u_wallace._1027_ ),
    .A2(\u_cpu.ALU.u_wallace._1028_ ),
    .B1(\u_cpu.ALU.u_wallace._1029_ ),
    .C1(\u_cpu.ALU.u_wallace._1031_ ),
    .Y(\u_cpu.ALU.u_wallace._1032_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6784_  (.A(\u_cpu.ALU.u_wallace._3623_ ),
    .B(\u_cpu.ALU.u_wallace._4447_ ),
    .C(\u_cpu.ALU.u_wallace._4731_ ),
    .D(\u_cpu.ALU.u_wallace._0365_ ),
    .Y(\u_cpu.ALU.u_wallace._1033_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6785_  (.A1(\u_cpu.ALU.u_wallace._3645_ ),
    .A2(\u_cpu.ALU.u_wallace._4836_ ),
    .B1(\u_cpu.ALU.u_wallace._4841_ ),
    .B2(\u_cpu.ALU.u_wallace._2790_ ),
    .X(\u_cpu.ALU.u_wallace._1034_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6786_  (.A(\u_cpu.ALU.u_wallace._3777_ ),
    .B(\u_cpu.ALU.SrcB[13] ),
    .Y(\u_cpu.ALU.u_wallace._1035_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6787_  (.A1(\u_cpu.ALU.u_wallace._1033_ ),
    .A2(\u_cpu.ALU.u_wallace._1034_ ),
    .B1(\u_cpu.ALU.u_wallace._1035_ ),
    .X(\u_cpu.ALU.u_wallace._1036_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6788_  (.A1(\u_cpu.ALU.u_wallace._4454_ ),
    .A2(\u_cpu.ALU.u_wallace._0037_ ),
    .B1(\u_cpu.ALU.u_wallace._1033_ ),
    .C1(\u_cpu.ALU.u_wallace._1034_ ),
    .Y(\u_cpu.ALU.u_wallace._1038_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6789_  (.A1(\u_cpu.ALU.u_wallace._1028_ ),
    .A2(\u_cpu.ALU.u_wallace._1027_ ),
    .B1(\u_cpu.ALU.u_wallace._1031_ ),
    .Y(\u_cpu.ALU.u_wallace._1039_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._6790_  (.A1(\u_cpu.ALU.u_wallace._4676_ ),
    .A2(\u_cpu.ALU.u_wallace._4601_ ),
    .A3(\u_cpu.ALU.u_wallace._0880_ ),
    .B1(\u_cpu.ALU.u_wallace._0898_ ),
    .X(\u_cpu.ALU.u_wallace._1040_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6791_  (.A1(\u_cpu.ALU.u_wallace._1036_ ),
    .A2(\u_cpu.ALU.u_wallace._1038_ ),
    .B1(\u_cpu.ALU.u_wallace._1039_ ),
    .B2(\u_cpu.ALU.u_wallace._1040_ ),
    .Y(\u_cpu.ALU.u_wallace._1041_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6792_  (.A(\u_cpu.ALU.u_wallace._0846_ ),
    .B(\u_cpu.ALU.u_wallace._0864_ ),
    .C(\u_cpu.ALU.u_wallace._0848_ ),
    .Y(\u_cpu.ALU.u_wallace._1042_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._6793_  (.A(\u_cpu.ALU.u_wallace._1028_ ),
    .B(\u_cpu.ALU.u_wallace._1027_ ),
    .Y(\u_cpu.ALU.u_wallace._1043_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6794_  (.A1(\u_cpu.ALU.u_wallace._4595_ ),
    .A2(\u_cpu.ALU.u_wallace._4642_ ),
    .B1(\u_cpu.ALU.u_wallace._4653_ ),
    .B2(\u_cpu.ALU.u_wallace._4594_ ),
    .X(\u_cpu.ALU.u_wallace._1044_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6795_  (.A1(\u_cpu.ALU.u_wallace._4783_ ),
    .A2(\u_cpu.ALU.u_wallace._0052_ ),
    .B1(\u_cpu.ALU.u_wallace._1044_ ),
    .B2(\u_cpu.ALU.u_wallace._1025_ ),
    .Y(\u_cpu.ALU.u_wallace._1045_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6796_  (.A1(\u_cpu.ALU.u_wallace._1043_ ),
    .A2(\u_cpu.ALU.u_wallace._1045_ ),
    .B1(\u_cpu.ALU.u_wallace._1040_ ),
    .Y(\u_cpu.ALU.u_wallace._1046_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6797_  (.A1(\u_cpu.ALU.u_wallace._4449_ ),
    .A2(\u_cpu.ALU.u_wallace._0028_ ),
    .B1(\u_cpu.ALU.u_wallace._4838_ ),
    .B2(\u_cpu.ALU.u_wallace._2725_ ),
    .Y(\u_cpu.ALU.u_wallace._1047_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._6798_  (.A1(\u_cpu.ALU.u_wallace._4660_ ),
    .A2(\u_cpu.ALU.u_wallace._3821_ ),
    .A3(\u_cpu.ALU.u_wallace._4840_ ),
    .A4(\u_cpu.ALU.u_wallace._4838_ ),
    .B1(\u_cpu.ALU.u_wallace._1035_ ),
    .X(\u_cpu.ALU.u_wallace._1049_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6799_  (.A1(\u_cpu.ALU.u_wallace._4452_ ),
    .A2(\u_cpu.ALU.u_wallace._0033_ ),
    .B1(\u_cpu.ALU.u_wallace._1033_ ),
    .B2(\u_cpu.ALU.u_wallace._1034_ ),
    .X(\u_cpu.ALU.u_wallace._1050_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6800_  (.A1(\u_cpu.ALU.u_wallace._1047_ ),
    .A2(\u_cpu.ALU.u_wallace._1049_ ),
    .B1(\u_cpu.ALU.u_wallace._1050_ ),
    .Y(\u_cpu.ALU.u_wallace._1051_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._6801_  (.A1(\u_cpu.ALU.u_wallace._1032_ ),
    .A2(\u_cpu.ALU.u_wallace._1046_ ),
    .B1_N(\u_cpu.ALU.u_wallace._1051_ ),
    .Y(\u_cpu.ALU.u_wallace._1052_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.ALU.u_wallace._6802_  (.A1(\u_cpu.ALU.u_wallace._1032_ ),
    .A2(\u_cpu.ALU.u_wallace._1041_ ),
    .B1(\u_cpu.ALU.u_wallace._0864_ ),
    .B2(\u_cpu.ALU.u_wallace._1042_ ),
    .C1(\u_cpu.ALU.u_wallace._1052_ ),
    .Y(\u_cpu.ALU.u_wallace._1053_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6803_  (.A1(\u_cpu.ALU.u_wallace._0890_ ),
    .A2(\u_cpu.ALU.u_wallace._0891_ ),
    .B1(\u_cpu.ALU.u_wallace._0900_ ),
    .Y(\u_cpu.ALU.u_wallace._1054_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6804_  (.A1(\u_cpu.ALU.u_wallace._0855_ ),
    .A2(\u_cpu.ALU.u_wallace._0856_ ),
    .B1(\u_cpu.ALU.u_wallace._0864_ ),
    .Y(\u_cpu.ALU.u_wallace._1055_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6805_  (.A(\u_cpu.ALU.u_wallace._1032_ ),
    .B(\u_cpu.ALU.u_wallace._1046_ ),
    .Y(\u_cpu.ALU.u_wallace._1056_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6806_  (.A1(\u_cpu.ALU.u_wallace._1032_ ),
    .A2(\u_cpu.ALU.u_wallace._1041_ ),
    .B1(\u_cpu.ALU.u_wallace._1056_ ),
    .B2(\u_cpu.ALU.u_wallace._1051_ ),
    .Y(\u_cpu.ALU.u_wallace._1057_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6807_  (.A1(\u_cpu.ALU.u_wallace._0886_ ),
    .A2(\u_cpu.ALU.u_wallace._1054_ ),
    .B1(\u_cpu.ALU.u_wallace._1055_ ),
    .B2(\u_cpu.ALU.u_wallace._1057_ ),
    .Y(\u_cpu.ALU.u_wallace._1058_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6808_  (.A1(\u_cpu.ALU.u_wallace._1027_ ),
    .A2(\u_cpu.ALU.u_wallace._1028_ ),
    .B1(\u_cpu.ALU.u_wallace._1029_ ),
    .C1(\u_cpu.ALU.u_wallace._1031_ ),
    .X(\u_cpu.ALU.u_wallace._1060_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.ALU.u_wallace._6809_  (.A1(\u_cpu.ALU.u_wallace._1036_ ),
    .A2(\u_cpu.ALU.u_wallace._1038_ ),
    .B1(\u_cpu.ALU.u_wallace._1040_ ),
    .B2(\u_cpu.ALU.u_wallace._1039_ ),
    .C1(\u_cpu.ALU.u_wallace._1060_ ),
    .Y(\u_cpu.ALU.u_wallace._1061_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._6810_  (.A(\u_cpu.ALU.u_wallace._0855_ ),
    .B(\u_cpu.ALU.u_wallace._0856_ ),
    .Y(\u_cpu.ALU.u_wallace._1062_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6811_  (.A(\u_cpu.ALU.u_wallace._1044_ ),
    .B(\u_cpu.ALU.u_wallace._1025_ ),
    .C(\u_cpu.ALU.u_wallace._0607_ ),
    .D(\u_cpu.ALU.u_wallace._4610_ ),
    .Y(\u_cpu.ALU.u_wallace._1063_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6812_  (.A1(\u_cpu.ALU.u_wallace._1063_ ),
    .A2(\u_cpu.ALU.u_wallace._1031_ ),
    .B1(\u_cpu.ALU.u_wallace._1029_ ),
    .Y(\u_cpu.ALU.u_wallace._1064_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6813_  (.A1(\u_cpu.ALU.u_wallace._1060_ ),
    .A2(\u_cpu.ALU.u_wallace._1064_ ),
    .B1(\u_cpu.ALU.u_wallace._1051_ ),
    .Y(\u_cpu.ALU.u_wallace._1065_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6814_  (.A1(\u_cpu.ALU.u_wallace._0854_ ),
    .A2(\u_cpu.ALU.u_wallace._1062_ ),
    .B1(\u_cpu.ALU.u_wallace._1065_ ),
    .Y(\u_cpu.ALU.u_wallace._1066_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._6815_  (.A1(\u_cpu.ALU.u_wallace._1061_ ),
    .A2(\u_cpu.ALU.u_wallace._1052_ ),
    .B1_N(\u_cpu.ALU.u_wallace._1055_ ),
    .Y(\u_cpu.ALU.u_wallace._1067_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6816_  (.A1(\u_cpu.ALU.u_wallace._1061_ ),
    .A2(\u_cpu.ALU.u_wallace._1066_ ),
    .B1(\u_cpu.ALU.u_wallace._1067_ ),
    .Y(\u_cpu.ALU.u_wallace._1068_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6817_  (.A1(\u_cpu.ALU.u_wallace._0892_ ),
    .A2(\u_cpu.ALU.u_wallace._0896_ ),
    .B1(\u_cpu.ALU.u_wallace._0886_ ),
    .Y(\u_cpu.ALU.u_wallace._1069_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._6818_  (.A1_N(\u_cpu.ALU.u_wallace._1053_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1058_ ),
    .B1(\u_cpu.ALU.u_wallace._1068_ ),
    .B2(\u_cpu.ALU.u_wallace._1069_ ),
    .Y(\u_cpu.ALU.u_wallace._1071_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6819_  (.A1(\u_cpu.ALU.u_wallace._0800_ ),
    .A2(\u_cpu.ALU.u_wallace._0803_ ),
    .B1(\u_cpu.ALU.u_wallace._0811_ ),
    .Y(\u_cpu.ALU.u_wallace._1072_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6820_  (.A(\u_cpu.ALU.SrcA[17] ),
    .X(\u_cpu.ALU.u_wallace._1073_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6821_  (.A1(\u_cpu.ALU.u_wallace._0490_ ),
    .A2(\u_cpu.ALU.u_wallace._0441_ ),
    .B1(\u_cpu.ALU.u_wallace._1073_ ),
    .B2(\u_cpu.ALU.u_wallace._0206_ ),
    .Y(\u_cpu.ALU.u_wallace._1074_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6822_  (.A(\u_cpu.ALU.u_wallace._0448_ ),
    .X(\u_cpu.ALU.u_wallace._1075_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6823_  (.A(\u_cpu.ALU.u_wallace._0457_ ),
    .B(\u_cpu.ALU.u_wallace._0330_ ),
    .Y(\u_cpu.ALU.u_wallace._1076_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._6824_  (.A1(\u_cpu.ALU.u_wallace._0217_ ),
    .A2(\u_cpu.ALU.u_wallace._4796_ ),
    .A3(\u_cpu.ALU.u_wallace._1075_ ),
    .A4(\u_cpu.ALU.u_wallace._0642_ ),
    .B1(\u_cpu.ALU.u_wallace._1076_ ),
    .X(\u_cpu.ALU.u_wallace._1077_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6825_  (.A1(\u_cpu.ALU.u_wallace._0578_ ),
    .A2(\u_cpu.ALU.u_wallace._0826_ ),
    .B1(\u_cpu.ALU.u_wallace._0822_ ),
    .B2(\u_cpu.ALU.u_wallace._0820_ ),
    .X(\u_cpu.ALU.u_wallace._1078_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6826_  (.A1(\u_cpu.ALU.u_wallace._1074_ ),
    .A2(\u_cpu.ALU.u_wallace._1077_ ),
    .B1(\u_cpu.ALU.u_wallace._1078_ ),
    .Y(\u_cpu.ALU.u_wallace._1079_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6827_  (.A1(\u_cpu.ALU.u_wallace._1072_ ),
    .A2(\u_cpu.ALU.u_wallace._0832_ ),
    .B1(\u_cpu.ALU.u_wallace._1079_ ),
    .Y(\u_cpu.ALU.u_wallace._1080_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6828_  (.A(\u_cpu.ALU.u_wallace._0457_ ),
    .B(\u_cpu.ALU.u_wallace._0448_ ),
    .Y(\u_cpu.ALU.u_wallace._1082_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._6829_  (.A1(\u_cpu.ALU.u_wallace._1158_ ),
    .A2(\u_cpu.ALU.u_wallace._1169_ ),
    .A3(\u_cpu.ALU.u_wallace._0642_ ),
    .A4(\u_cpu.ALU.u_wallace._0802_ ),
    .B1(\u_cpu.ALU.u_wallace._1082_ ),
    .X(\u_cpu.ALU.u_wallace._1083_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6830_  (.A(\u_cpu.ALU.SrcA[18] ),
    .X(\u_cpu.ALU.u_wallace._1084_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6831_  (.A1(\u_cpu.ALU.u_wallace._0490_ ),
    .A2(\u_cpu.ALU.u_wallace._1073_ ),
    .B1(\u_cpu.ALU.u_wallace._1084_ ),
    .B2(\u_cpu.ALU.u_wallace._0206_ ),
    .Y(\u_cpu.ALU.u_wallace._1085_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6832_  (.A1(\u_cpu.ALU.u_wallace._0293_ ),
    .A2(\u_cpu.ALU.u_wallace._0630_ ),
    .B1(\u_cpu.ALU.u_wallace._0808_ ),
    .B2(\u_cpu.ALU.u_wallace._0797_ ),
    .X(\u_cpu.ALU.u_wallace._1086_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6833_  (.A(\u_cpu.ALU.u_wallace._0206_ ),
    .B(\u_cpu.ALU.u_wallace._1914_ ),
    .C(\u_cpu.ALU.u_wallace._0630_ ),
    .D(\u_cpu.ALU.u_wallace._1084_ ),
    .Y(\u_cpu.ALU.u_wallace._1087_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6834_  (.A1(\u_cpu.ALU.u_wallace._0840_ ),
    .A2(\u_cpu.ALU.u_wallace._0850_ ),
    .B1(\u_cpu.ALU.u_wallace._1086_ ),
    .B2(\u_cpu.ALU.u_wallace._1087_ ),
    .X(\u_cpu.ALU.u_wallace._1088_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6835_  (.A(\u_cpu.ALU.u_wallace._2768_ ),
    .B(\u_cpu.ALU.SrcA[2] ),
    .C(\u_cpu.ALU.u_wallace._4920_ ),
    .D(\u_cpu.ALU.u_wallace._0813_ ),
    .Y(\u_cpu.ALU.u_wallace._1089_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6836_  (.A(\u_cpu.ALU.SrcA[19] ),
    .X(\u_cpu.ALU.u_wallace._1090_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6837_  (.A(\u_cpu.ALU.u_wallace._1089_ ),
    .B(\u_cpu.ALU.u_wallace._1090_ ),
    .C(\u_cpu.ALU.u_wallace._0873_ ),
    .Y(\u_cpu.ALU.u_wallace._1091_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6838_  (.A1(\u_cpu.ALU.u_wallace._1760_ ),
    .A2(\u_cpu.ALU.SrcA[13] ),
    .B1(\u_cpu.ALU.u_wallace._0626_ ),
    .B2(\u_cpu.ALU.SrcA[2] ),
    .Y(\u_cpu.ALU.u_wallace._1093_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6839_  (.A(\u_cpu.ALU.u_wallace._0075_ ),
    .B(\u_cpu.ALU.u_wallace._1084_ ),
    .Y(\u_cpu.ALU.u_wallace._1094_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6840_  (.A1(\u_cpu.ALU.u_wallace._1094_ ),
    .A2(\u_cpu.ALU.u_wallace._0800_ ),
    .B1(\u_cpu.ALU.u_wallace._0801_ ),
    .Y(\u_cpu.ALU.u_wallace._1095_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._6841_  (.A(\u_cpu.ALU.SrcA[19] ),
    .Y(\u_cpu.ALU.u_wallace._1096_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6842_  (.A(\u_cpu.ALU.u_wallace._4649_ ),
    .B(\u_cpu.ALU.SrcA[2] ),
    .C(\u_cpu.ALU.u_wallace._4920_ ),
    .D(\u_cpu.ALU.u_wallace._0628_ ),
    .X(\u_cpu.ALU.u_wallace._1097_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6843_  (.A1(\u_cpu.ALU.u_wallace._0634_ ),
    .A2(\u_cpu.ALU.u_wallace._1096_ ),
    .B1(\u_cpu.ALU.u_wallace._1093_ ),
    .B2(\u_cpu.ALU.u_wallace._1097_ ),
    .Y(\u_cpu.ALU.u_wallace._1098_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6844_  (.A1(\u_cpu.ALU.u_wallace._1091_ ),
    .A2(\u_cpu.ALU.u_wallace._1093_ ),
    .B1(\u_cpu.ALU.u_wallace._1095_ ),
    .C1(\u_cpu.ALU.u_wallace._1098_ ),
    .Y(\u_cpu.ALU.u_wallace._1099_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6845_  (.A(\u_cpu.ALU.SrcA[19] ),
    .X(\u_cpu.ALU.u_wallace._1100_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6846_  (.A(\u_cpu.ALU.u_wallace._1100_ ),
    .X(\u_cpu.ALU.u_wallace._1101_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6847_  (.A(\u_cpu.ALU.SrcB[17] ),
    .X(\u_cpu.ALU.u_wallace._1102_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6848_  (.A1(\u_cpu.ALU.u_wallace._4645_ ),
    .A2(\u_cpu.ALU.u_wallace._4907_ ),
    .B1(\u_cpu.ALU.u_wallace._1102_ ),
    .B2(\u_cpu.ALU.u_wallace._0348_ ),
    .X(\u_cpu.ALU.u_wallace._1104_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6849_  (.A1(\u_cpu.ALU.u_wallace._2757_ ),
    .A2(\u_cpu.ALU.u_wallace._1101_ ),
    .B1(\u_cpu.ALU.u_wallace._1104_ ),
    .B2(\u_cpu.ALU.u_wallace._1089_ ),
    .Y(\u_cpu.ALU.u_wallace._1105_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._6850_  (.A(\u_cpu.ALU.u_wallace._1093_ ),
    .B(\u_cpu.ALU.u_wallace._1091_ ),
    .Y(\u_cpu.ALU.u_wallace._1106_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._6851_  (.A1(\u_cpu.ALU.u_wallace._1105_ ),
    .A2(\u_cpu.ALU.u_wallace._1106_ ),
    .B1_N(\u_cpu.ALU.u_wallace._1095_ ),
    .Y(\u_cpu.ALU.u_wallace._1107_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._6852_  (.A1(\u_cpu.ALU.u_wallace._1083_ ),
    .A2(\u_cpu.ALU.u_wallace._1085_ ),
    .B1(\u_cpu.ALU.u_wallace._1088_ ),
    .C1(\u_cpu.ALU.u_wallace._1099_ ),
    .D1(\u_cpu.ALU.u_wallace._1107_ ),
    .Y(\u_cpu.ALU.u_wallace._1108_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6853_  (.A1(\u_cpu.ALU.u_wallace._0468_ ),
    .A2(\u_cpu.ALU.u_wallace._1075_ ),
    .B1(\u_cpu.ALU.u_wallace._1086_ ),
    .B2(\u_cpu.ALU.u_wallace._1087_ ),
    .Y(\u_cpu.ALU.u_wallace._1109_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6854_  (.A(\u_cpu.ALU.u_wallace._1086_ ),
    .B(\u_cpu.ALU.u_wallace._1087_ ),
    .C(\u_cpu.ALU.u_wallace._4662_ ),
    .D(\u_cpu.ALU.u_wallace._1075_ ),
    .X(\u_cpu.ALU.u_wallace._1110_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6855_  (.A1(\u_cpu.ALU.u_wallace._1091_ ),
    .A2(\u_cpu.ALU.u_wallace._1093_ ),
    .B1(\u_cpu.ALU.u_wallace._1095_ ),
    .C1(\u_cpu.ALU.u_wallace._1098_ ),
    .X(\u_cpu.ALU.u_wallace._1111_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6856_  (.A(\u_cpu.ALU.u_wallace._1104_ ),
    .B(\u_cpu.ALU.u_wallace._1089_ ),
    .C(\u_cpu.ALU.u_wallace._0086_ ),
    .D(\u_cpu.ALU.u_wallace._1101_ ),
    .Y(\u_cpu.ALU.u_wallace._1112_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6857_  (.A1(\u_cpu.ALU.u_wallace._1098_ ),
    .A2(\u_cpu.ALU.u_wallace._1112_ ),
    .B1(\u_cpu.ALU.u_wallace._1095_ ),
    .Y(\u_cpu.ALU.u_wallace._1113_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6858_  (.A1(\u_cpu.ALU.u_wallace._1109_ ),
    .A2(\u_cpu.ALU.u_wallace._1110_ ),
    .B1(\u_cpu.ALU.u_wallace._1111_ ),
    .B2(\u_cpu.ALU.u_wallace._1113_ ),
    .Y(\u_cpu.ALU.u_wallace._1115_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6859_  (.A1(\u_cpu.ALU.u_wallace._0812_ ),
    .A2(\u_cpu.ALU.u_wallace._1080_ ),
    .B1(\u_cpu.ALU.u_wallace._1108_ ),
    .C1(\u_cpu.ALU.u_wallace._1115_ ),
    .Y(\u_cpu.ALU.u_wallace._1116_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6860_  (.A1(\u_cpu.ALU.u_wallace._1085_ ),
    .A2(\u_cpu.ALU.u_wallace._1083_ ),
    .B1(\u_cpu.ALU.u_wallace._1088_ ),
    .Y(\u_cpu.ALU.u_wallace._1117_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._6861_  (.A1(\u_cpu.ALU.u_wallace._1111_ ),
    .A2(\u_cpu.ALU.u_wallace._1113_ ),
    .B1_N(\u_cpu.ALU.u_wallace._1117_ ),
    .Y(\u_cpu.ALU.u_wallace._1118_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6862_  (.A1(\u_cpu.ALU.u_wallace._1109_ ),
    .A2(\u_cpu.ALU.u_wallace._1110_ ),
    .B1(\u_cpu.ALU.u_wallace._1099_ ),
    .C1(\u_cpu.ALU.u_wallace._1107_ ),
    .Y(\u_cpu.ALU.u_wallace._1119_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._6863_  (.A1_N(\u_cpu.ALU.u_wallace._0828_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0830_ ),
    .B1(\u_cpu.ALU.u_wallace._0824_ ),
    .B2(\u_cpu.ALU.u_wallace._0833_ ),
    .Y(\u_cpu.ALU.u_wallace._1120_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6864_  (.A(\u_cpu.ALU.u_wallace._1118_ ),
    .B(\u_cpu.ALU.u_wallace._1119_ ),
    .C(\u_cpu.ALU.u_wallace._1120_ ),
    .Y(\u_cpu.ALU.u_wallace._1121_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6865_  (.A(\u_cpu.ALU.u_wallace._2144_ ),
    .B(\u_cpu.ALU.u_wallace._2538_ ),
    .C(\u_cpu.ALU.u_wallace._0182_ ),
    .D(\u_cpu.ALU.u_wallace._0332_ ),
    .Y(\u_cpu.ALU.u_wallace._1122_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6866_  (.A1(\u_cpu.ALU.u_wallace._1541_ ),
    .A2(\u_cpu.ALU.u_wallace._0182_ ),
    .B1(\u_cpu.ALU.u_wallace._0332_ ),
    .B2(\u_cpu.ALU.u_wallace._1026_ ),
    .X(\u_cpu.ALU.u_wallace._1123_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6867_  (.A1_N(\u_cpu.ALU.u_wallace._1122_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1123_ ),
    .B1(\u_cpu.ALU.u_wallace._4471_ ),
    .B2(\u_cpu.ALU.u_wallace._4913_ ),
    .Y(\u_cpu.ALU.u_wallace._1124_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6868_  (.A(\u_cpu.ALU.u_wallace._1123_ ),
    .B(\u_cpu.ALU.u_wallace._4917_ ),
    .C(\u_cpu.ALU.u_wallace._3404_ ),
    .D(\u_cpu.ALU.u_wallace._1122_ ),
    .Y(\u_cpu.ALU.u_wallace._1126_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6869_  (.A1(\u_cpu.ALU.u_wallace._1076_ ),
    .A2(\u_cpu.ALU.u_wallace._1074_ ),
    .B1(\u_cpu.ALU.u_wallace._0820_ ),
    .Y(\u_cpu.ALU.u_wallace._1127_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6870_  (.A(\u_cpu.ALU.u_wallace._1124_ ),
    .B(\u_cpu.ALU.u_wallace._1126_ ),
    .C(\u_cpu.ALU.u_wallace._1127_ ),
    .X(\u_cpu.ALU.u_wallace._1128_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6871_  (.A(\u_cpu.ALU.u_wallace._4794_ ),
    .X(\u_cpu.ALU.u_wallace._1129_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._6872_  (.A1(\u_cpu.ALU.u_wallace._0839_ ),
    .A2(\u_cpu.ALU.u_wallace._1129_ ),
    .A3(\u_cpu.ALU.u_wallace._3481_ ),
    .B1(\u_cpu.ALU.u_wallace._0837_ ),
    .X(\u_cpu.ALU.u_wallace._1130_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6873_  (.A1(\u_cpu.ALU.u_wallace._1124_ ),
    .A2(\u_cpu.ALU.u_wallace._1126_ ),
    .B1(\u_cpu.ALU.u_wallace._1127_ ),
    .X(\u_cpu.ALU.u_wallace._1131_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6874_  (.A(\u_cpu.ALU.u_wallace._1130_ ),
    .B(\u_cpu.ALU.u_wallace._1131_ ),
    .Y(\u_cpu.ALU.u_wallace._1132_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6875_  (.A1(\u_cpu.ALU.u_wallace._1124_ ),
    .A2(\u_cpu.ALU.u_wallace._1126_ ),
    .B1(\u_cpu.ALU.u_wallace._1127_ ),
    .Y(\u_cpu.ALU.u_wallace._1133_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._6876_  (.A1(\u_cpu.ALU.u_wallace._4539_ ),
    .A2(\u_cpu.ALU.u_wallace._0169_ ),
    .A3(\u_cpu.ALU.u_wallace._0836_ ),
    .B1(\u_cpu.ALU.u_wallace._0841_ ),
    .X(\u_cpu.ALU.u_wallace._1134_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6877_  (.A1(\u_cpu.ALU.u_wallace._1133_ ),
    .A2(\u_cpu.ALU.u_wallace._1128_ ),
    .B1(\u_cpu.ALU.u_wallace._1134_ ),
    .Y(\u_cpu.ALU.u_wallace._1135_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6878_  (.A1(\u_cpu.ALU.u_wallace._1128_ ),
    .A2(\u_cpu.ALU.u_wallace._1132_ ),
    .B1(\u_cpu.ALU.u_wallace._1135_ ),
    .Y(\u_cpu.ALU.u_wallace._1137_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6879_  (.A1(\u_cpu.ALU.u_wallace._1116_ ),
    .A2(\u_cpu.ALU.u_wallace._1121_ ),
    .B1(\u_cpu.ALU.u_wallace._1137_ ),
    .X(\u_cpu.ALU.u_wallace._1138_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6880_  (.A(\u_cpu.ALU.u_wallace._1124_ ),
    .B(\u_cpu.ALU.u_wallace._1126_ ),
    .C(\u_cpu.ALU.u_wallace._1127_ ),
    .Y(\u_cpu.ALU.u_wallace._1139_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6881_  (.A1(\u_cpu.ALU.u_wallace._1131_ ),
    .A2(\u_cpu.ALU.u_wallace._1139_ ),
    .B1(\u_cpu.ALU.u_wallace._1130_ ),
    .Y(\u_cpu.ALU.u_wallace._1140_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6882_  (.A(\u_cpu.ALU.u_wallace._1130_ ),
    .B(\u_cpu.ALU.u_wallace._1131_ ),
    .C(\u_cpu.ALU.u_wallace._1139_ ),
    .X(\u_cpu.ALU.u_wallace._1141_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6883_  (.A(\u_cpu.ALU.u_wallace._1087_ ),
    .B(\u_cpu.ALU.u_wallace._0850_ ),
    .C(\u_cpu.ALU.u_wallace._0840_ ),
    .X(\u_cpu.ALU.u_wallace._1142_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6884_  (.A1(\u_cpu.ALU.u_wallace._1142_ ),
    .A2(\u_cpu.ALU.u_wallace._1086_ ),
    .B1(\u_cpu.ALU.u_wallace._1109_ ),
    .Y(\u_cpu.ALU.u_wallace._1143_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6885_  (.A(\u_cpu.ALU.u_wallace._1107_ ),
    .B(\u_cpu.ALU.u_wallace._1143_ ),
    .C(\u_cpu.ALU.u_wallace._1099_ ),
    .X(\u_cpu.ALU.u_wallace._1144_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6886_  (.A1(\u_cpu.ALU.u_wallace._0812_ ),
    .A2(\u_cpu.ALU.u_wallace._1080_ ),
    .B1(\u_cpu.ALU.u_wallace._1115_ ),
    .Y(\u_cpu.ALU.u_wallace._1145_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._6887_  (.A1(\u_cpu.ALU.u_wallace._1140_ ),
    .A2(\u_cpu.ALU.u_wallace._1141_ ),
    .B1(\u_cpu.ALU.u_wallace._1144_ ),
    .B2(\u_cpu.ALU.u_wallace._1145_ ),
    .C1(\u_cpu.ALU.u_wallace._1121_ ),
    .Y(\u_cpu.ALU.u_wallace._1146_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6888_  (.A1(\u_cpu.ALU.u_wallace._1062_ ),
    .A2(\u_cpu.ALU.u_wallace._0864_ ),
    .B1(\u_cpu.ALU.u_wallace._0865_ ),
    .Y(\u_cpu.ALU.u_wallace._1148_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6889_  (.A1(\u_cpu.ALU.u_wallace._1148_ ),
    .A2(\u_cpu.ALU.u_wallace._0859_ ),
    .B1(\u_cpu.ALU.u_wallace._0835_ ),
    .Y(\u_cpu.ALU.u_wallace._1149_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6890_  (.A(\u_cpu.ALU.u_wallace._1138_ ),
    .B(\u_cpu.ALU.u_wallace._1146_ ),
    .C(\u_cpu.ALU.u_wallace._1149_ ),
    .Y(\u_cpu.ALU.u_wallace._1150_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6891_  (.A1(\u_cpu.ALU.u_wallace._1118_ ),
    .A2(\u_cpu.ALU.u_wallace._1119_ ),
    .B1(\u_cpu.ALU.u_wallace._1120_ ),
    .Y(\u_cpu.ALU.u_wallace._1151_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6892_  (.A1(\u_cpu.ALU.u_wallace._1132_ ),
    .A2(\u_cpu.ALU.u_wallace._1128_ ),
    .B1(\u_cpu.ALU.u_wallace._1135_ ),
    .C1(\u_cpu.ALU.u_wallace._1121_ ),
    .Y(\u_cpu.ALU.u_wallace._1152_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._6893_  (.A1(\u_cpu.ALU.u_wallace._0858_ ),
    .A2(\u_cpu.ALU.u_wallace._0825_ ),
    .A3(\u_cpu.ALU.u_wallace._0834_ ),
    .B1(\u_cpu.ALU.u_wallace._0913_ ),
    .Y(\u_cpu.ALU.u_wallace._1153_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._6894_  (.A1(\u_cpu.ALU.u_wallace._0817_ ),
    .A2(\u_cpu.ALU.u_wallace._0811_ ),
    .A3(\u_cpu.ALU.u_wallace._0816_ ),
    .B1(\u_cpu.ALU.u_wallace._0833_ ),
    .B2(\u_cpu.ALU.u_wallace._0824_ ),
    .X(\u_cpu.ALU.u_wallace._1154_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6895_  (.A1(\u_cpu.ALU.u_wallace._1108_ ),
    .A2(\u_cpu.ALU.u_wallace._1115_ ),
    .B1(\u_cpu.ALU.u_wallace._1154_ ),
    .Y(\u_cpu.ALU.u_wallace._1155_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6896_  (.A1(\u_cpu.ALU.u_wallace._1140_ ),
    .A2(\u_cpu.ALU.u_wallace._1141_ ),
    .B1(\u_cpu.ALU.u_wallace._1151_ ),
    .B2(\u_cpu.ALU.u_wallace._1155_ ),
    .Y(\u_cpu.ALU.u_wallace._1156_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._6897_  (.A1(\u_cpu.ALU.u_wallace._1151_ ),
    .A2(\u_cpu.ALU.u_wallace._1152_ ),
    .B1(\u_cpu.ALU.u_wallace._0835_ ),
    .B2(\u_cpu.ALU.u_wallace._1153_ ),
    .C1(\u_cpu.ALU.u_wallace._1156_ ),
    .Y(\u_cpu.ALU.u_wallace._1157_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6898_  (.A(\u_cpu.ALU.u_wallace._1071_ ),
    .B(\u_cpu.ALU.u_wallace._1150_ ),
    .C(\u_cpu.ALU.u_wallace._1157_ ),
    .Y(\u_cpu.ALU.u_wallace._1159_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._6899_  (.A1(\u_cpu.ALU.u_wallace._0886_ ),
    .A2(\u_cpu.ALU.u_wallace._1054_ ),
    .B1(\u_cpu.ALU.u_wallace._1061_ ),
    .B2(\u_cpu.ALU.u_wallace._1066_ ),
    .C1(\u_cpu.ALU.u_wallace._1067_ ),
    .X(\u_cpu.ALU.u_wallace._1160_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU.u_wallace._6900_  (.A1(\u_cpu.ALU.u_wallace._1032_ ),
    .A2(\u_cpu.ALU.u_wallace._1041_ ),
    .B1(\u_cpu.ALU.u_wallace._0864_ ),
    .B2(\u_cpu.ALU.u_wallace._1042_ ),
    .C1(\u_cpu.ALU.u_wallace._1052_ ),
    .X(\u_cpu.ALU.u_wallace._1161_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._6901_  (.A1(\u_cpu.ALU.u_wallace._0882_ ),
    .A2(\u_cpu.ALU.u_wallace._0899_ ),
    .A3(\u_cpu.ALU.u_wallace._0885_ ),
    .B1(\u_cpu.ALU.u_wallace._1054_ ),
    .X(\u_cpu.ALU.u_wallace._1162_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6902_  (.A1(\u_cpu.ALU.u_wallace._1161_ ),
    .A2(\u_cpu.ALU.u_wallace._1067_ ),
    .B1(\u_cpu.ALU.u_wallace._1162_ ),
    .Y(\u_cpu.ALU.u_wallace._1163_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6903_  (.A1_N(\u_cpu.ALU.u_wallace._1157_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1150_ ),
    .B1(\u_cpu.ALU.u_wallace._1160_ ),
    .B2(\u_cpu.ALU.u_wallace._1163_ ),
    .Y(\u_cpu.ALU.u_wallace._1164_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6904_  (.A1(\u_cpu.ALU.u_wallace._0872_ ),
    .A2(\u_cpu.ALU.u_wallace._1024_ ),
    .B1(\u_cpu.ALU.u_wallace._1159_ ),
    .C1(\u_cpu.ALU.u_wallace._1164_ ),
    .X(\u_cpu.ALU.u_wallace._1165_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6905_  (.A1(\u_cpu.ALU.u_wallace._1116_ ),
    .A2(\u_cpu.ALU.u_wallace._1121_ ),
    .B1(\u_cpu.ALU.u_wallace._1137_ ),
    .Y(\u_cpu.ALU.u_wallace._1166_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6906_  (.A1(\u_cpu.ALU.u_wallace._1140_ ),
    .A2(\u_cpu.ALU.u_wallace._1141_ ),
    .B1(\u_cpu.ALU.u_wallace._1116_ ),
    .C1(\u_cpu.ALU.u_wallace._1121_ ),
    .X(\u_cpu.ALU.u_wallace._1167_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._6907_  (.A1(\u_cpu.ALU.u_wallace._0857_ ),
    .A2(\u_cpu.ALU.u_wallace._1042_ ),
    .A3(\u_cpu.ALU.u_wallace._0859_ ),
    .B1(\u_cpu.ALU.u_wallace._0835_ ),
    .X(\u_cpu.ALU.u_wallace._1168_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU.u_wallace._6908_  (.A1(\u_cpu.ALU.u_wallace._1166_ ),
    .A2(\u_cpu.ALU.u_wallace._1167_ ),
    .A3(\u_cpu.ALU.u_wallace._1168_ ),
    .B1(\u_cpu.ALU.u_wallace._1157_ ),
    .C1(\u_cpu.ALU.u_wallace._1071_ ),
    .X(\u_cpu.ALU.u_wallace._1170_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6909_  (.A1(\u_cpu.ALU.u_wallace._1157_ ),
    .A2(\u_cpu.ALU.u_wallace._1150_ ),
    .B1(\u_cpu.ALU.u_wallace._1071_ ),
    .Y(\u_cpu.ALU.u_wallace._1171_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6910_  (.A1(\u_cpu.ALU.u_wallace._0920_ ),
    .A2(\u_cpu.ALU.u_wallace._0981_ ),
    .B1(\u_cpu.ALU.u_wallace._0872_ ),
    .Y(\u_cpu.ALU.u_wallace._1172_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6911_  (.A1(\u_cpu.ALU.u_wallace._1170_ ),
    .A2(\u_cpu.ALU.u_wallace._1171_ ),
    .B1(\u_cpu.ALU.u_wallace._1172_ ),
    .Y(\u_cpu.ALU.u_wallace._1173_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._6912_  (.A1(\u_cpu.ALU.u_wallace._0874_ ),
    .A2(\u_cpu.ALU.u_wallace._0877_ ),
    .B1(\u_cpu.ALU.u_wallace._0886_ ),
    .B2(\u_cpu.ALU.u_wallace._0897_ ),
    .C1(\u_cpu.ALU.u_wallace._0901_ ),
    .X(\u_cpu.ALU.u_wallace._1174_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6913_  (.A(\u_cpu.ALU.SrcB[19] ),
    .X(\u_cpu.ALU.u_wallace._1175_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6914_  (.A(\u_cpu.ALU.u_wallace._1175_ ),
    .X(\u_cpu.ALU.u_wallace._1176_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6915_  (.A(\u_cpu.ALU.u_wallace._1070_ ),
    .B(\u_cpu.ALU.u_wallace._1176_ ),
    .Y(\u_cpu.ALU.u_wallace._1177_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6916_  (.A(\u_cpu.ALU.u_wallace._1177_ ),
    .B(\u_cpu.ALU.u_wallace._0959_ ),
    .C(\u_cpu.ALU.u_wallace._0184_ ),
    .X(\u_cpu.ALU.u_wallace._1178_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6917_  (.A(\u_cpu.ALU.u_wallace._0162_ ),
    .B(\u_cpu.ALU.u_wallace._0959_ ),
    .Y(\u_cpu.ALU.u_wallace._1179_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6918_  (.A(\u_cpu.ALU.u_wallace._1179_ ),
    .B(\u_cpu.ALU.u_wallace._1176_ ),
    .C(\u_cpu.ALU.u_wallace._3996_ ),
    .X(\u_cpu.ALU.u_wallace._1181_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6919_  (.A1(\u_cpu.ALU.u_wallace._3821_ ),
    .A2(\u_cpu.ALU.u_wallace._4837_ ),
    .B1(\u_cpu.ALU.u_wallace._4838_ ),
    .B2(\u_cpu.ALU.u_wallace._1848_ ),
    .Y(\u_cpu.ALU.u_wallace._1182_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._6920_  (.A1(\u_cpu.ALU.u_wallace._4813_ ),
    .A2(\u_cpu.ALU.u_wallace._0037_ ),
    .A3(\u_cpu.ALU.u_wallace._1182_ ),
    .B1(\u_cpu.ALU.u_wallace._0888_ ),
    .X(\u_cpu.ALU.u_wallace._1183_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._6921_  (.A1(\u_cpu.ALU.u_wallace._1311_ ),
    .A2(\u_cpu.ALU.u_wallace._0120_ ),
    .B1(\u_cpu.ALU.u_wallace._0728_ ),
    .B2(\u_cpu.ALU.u_wallace._4556_ ),
    .X(\u_cpu.ALU.u_wallace._1184_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6922_  (.A(\u_cpu.ALU.u_wallace._1125_ ),
    .B(\u_cpu.ALU.u_wallace._1267_ ),
    .C(\u_cpu.ALU.u_wallace._0730_ ),
    .D(\u_cpu.ALU.u_wallace._0732_ ),
    .Y(\u_cpu.ALU.u_wallace._1185_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._6923_  (.A(\u_cpu.ALU.u_wallace._1184_ ),
    .B(\u_cpu.ALU.u_wallace._1185_ ),
    .C(\u_cpu.ALU.u_wallace._1421_ ),
    .D(\u_cpu.ALU.u_wallace._0550_ ),
    .Y(\u_cpu.ALU.u_wallace._1186_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6924_  (.A1(\u_cpu.ALU.u_wallace._1125_ ),
    .A2(\u_cpu.ALU.u_wallace._0730_ ),
    .B1(\u_cpu.ALU.u_wallace._0547_ ),
    .B2(\u_cpu.ALU.u_wallace._1267_ ),
    .Y(\u_cpu.ALU.u_wallace._1187_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6925_  (.A(\u_cpu.ALU.u_wallace._2955_ ),
    .B(\u_cpu.ALU.u_wallace._4556_ ),
    .C(\u_cpu.ALU.u_wallace._0120_ ),
    .D(\u_cpu.ALU.u_wallace._0728_ ),
    .X(\u_cpu.ALU.u_wallace._1188_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6926_  (.A1(\u_cpu.ALU.u_wallace._0610_ ),
    .A2(\u_cpu.ALU.u_wallace._0941_ ),
    .B1(\u_cpu.ALU.u_wallace._1187_ ),
    .B2(\u_cpu.ALU.u_wallace._1188_ ),
    .Y(\u_cpu.ALU.u_wallace._1189_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6927_  (.A(\u_cpu.ALU.u_wallace._1186_ ),
    .B(\u_cpu.ALU.u_wallace._1189_ ),
    .Y(\u_cpu.ALU.u_wallace._1190_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._6928_  (.A(\u_cpu.ALU.u_wallace._0937_ ),
    .B(\u_cpu.ALU.u_wallace._0735_ ),
    .C(\u_cpu.ALU.u_wallace._4545_ ),
    .X(\u_cpu.ALU.u_wallace._1192_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._6929_  (.A1_N(\u_cpu.ALU.u_wallace._1183_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1190_ ),
    .B1(\u_cpu.ALU.u_wallace._0943_ ),
    .B2(\u_cpu.ALU.u_wallace._1192_ ),
    .Y(\u_cpu.ALU.u_wallace._1193_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6930_  (.A(\u_cpu.ALU.u_wallace._4450_ ),
    .B(\u_cpu.ALU.u_wallace._1793_ ),
    .C(\u_cpu.ALU.u_wallace._4731_ ),
    .D(\u_cpu.ALU.u_wallace._0365_ ),
    .X(\u_cpu.ALU.u_wallace._1194_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._6931_  (.A(\u_cpu.ALU.u_wallace._0889_ ),
    .B(\u_cpu.ALU.u_wallace._1182_ ),
    .Y(\u_cpu.ALU.u_wallace._1195_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6932_  (.A1(\u_cpu.ALU.u_wallace._1194_ ),
    .A2(\u_cpu.ALU.u_wallace._1195_ ),
    .B1(\u_cpu.ALU.u_wallace._1186_ ),
    .C1(\u_cpu.ALU.u_wallace._1189_ ),
    .X(\u_cpu.ALU.u_wallace._1196_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6933_  (.A1(\u_cpu.ALU.u_wallace._0931_ ),
    .A2(\u_cpu.ALU.u_wallace._0952_ ),
    .B1(\u_cpu.ALU.u_wallace._0945_ ),
    .Y(\u_cpu.ALU.u_wallace._1197_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._6934_  (.A1(\u_cpu.ALU.u_wallace._0887_ ),
    .A2(\u_cpu.ALU.u_wallace._0057_ ),
    .A3(\u_cpu.ALU.u_wallace._1136_ ),
    .B1(\u_cpu.ALU.u_wallace._1194_ ),
    .X(\u_cpu.ALU.u_wallace._1198_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6935_  (.A1(\u_cpu.ALU.u_wallace._1186_ ),
    .A2(\u_cpu.ALU.u_wallace._1189_ ),
    .B1(\u_cpu.ALU.u_wallace._1198_ ),
    .Y(\u_cpu.ALU.u_wallace._1199_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._6936_  (.A1(\u_cpu.ALU.u_wallace._0414_ ),
    .A2(\u_cpu.ALU.u_wallace._0554_ ),
    .A3(\u_cpu.ALU.u_wallace._0942_ ),
    .B1(\u_cpu.ALU.u_wallace._0938_ ),
    .X(\u_cpu.ALU.u_wallace._1200_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6937_  (.A1(\u_cpu.ALU.u_wallace._1196_ ),
    .A2(\u_cpu.ALU.u_wallace._1199_ ),
    .B1(\u_cpu.ALU.u_wallace._1200_ ),
    .Y(\u_cpu.ALU.u_wallace._1201_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6938_  (.A1(\u_cpu.ALU.u_wallace._1193_ ),
    .A2(\u_cpu.ALU.u_wallace._1196_ ),
    .B1(\u_cpu.ALU.u_wallace._1197_ ),
    .C1(\u_cpu.ALU.u_wallace._1201_ ),
    .Y(\u_cpu.ALU.u_wallace._1203_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._6939_  (.A1(\u_cpu.ALU.u_wallace._1194_ ),
    .A2(\u_cpu.ALU.u_wallace._1195_ ),
    .B1(\u_cpu.ALU.u_wallace._1189_ ),
    .X(\u_cpu.ALU.u_wallace._1204_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._6940_  (.A1(\u_cpu.ALU.u_wallace._1204_ ),
    .A2(\u_cpu.ALU.u_wallace._1186_ ),
    .B1(\u_cpu.ALU.u_wallace._1200_ ),
    .C1(\u_cpu.ALU.u_wallace._1199_ ),
    .X(\u_cpu.ALU.u_wallace._1205_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6941_  (.A1(\u_cpu.ALU.u_wallace._1205_ ),
    .A2(\u_cpu.ALU.u_wallace._1201_ ),
    .B1(\u_cpu.ALU.u_wallace._1197_ ),
    .X(\u_cpu.ALU.u_wallace._1206_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6942_  (.A1(\u_cpu.ALU.u_wallace._1178_ ),
    .A2(\u_cpu.ALU.u_wallace._1181_ ),
    .B1(\u_cpu.ALU.u_wallace._1203_ ),
    .C1(\u_cpu.ALU.u_wallace._1206_ ),
    .Y(\u_cpu.ALU.u_wallace._1207_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6943_  (.A(\u_cpu.ALU.SrcB[19] ),
    .X(\u_cpu.ALU.u_wallace._1208_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6944_  (.A(\u_cpu.ALU.u_wallace._0446_ ),
    .B(\u_cpu.ALU.u_wallace._1454_ ),
    .C(\u_cpu.ALU.u_wallace._0958_ ),
    .D(\u_cpu.ALU.u_wallace._1208_ ),
    .X(\u_cpu.ALU.u_wallace._1209_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._6945_  (.A(\u_cpu.ALU.SrcB[19] ),
    .X(\u_cpu.ALU.u_wallace._1210_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._6946_  (.A(\u_cpu.ALU.u_wallace._1210_ ),
    .Y(\u_cpu.ALU.u_wallace._1211_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU.u_wallace._6947_  (.A1_N(\u_cpu.ALU.u_wallace._0184_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0959_ ),
    .B1(\u_cpu.ALU.u_wallace._1211_ ),
    .B2(\u_cpu.ALU.u_wallace._0043_ ),
    .X(\u_cpu.ALU.u_wallace._1212_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._6948_  (.A1(\u_cpu.ALU.u_wallace._1193_ ),
    .A2(\u_cpu.ALU.u_wallace._1196_ ),
    .B1(\u_cpu.ALU.u_wallace._1197_ ),
    .C1(\u_cpu.ALU.u_wallace._1201_ ),
    .X(\u_cpu.ALU.u_wallace._1214_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6949_  (.A1(\u_cpu.ALU.u_wallace._1205_ ),
    .A2(\u_cpu.ALU.u_wallace._1201_ ),
    .B1(\u_cpu.ALU.u_wallace._1197_ ),
    .Y(\u_cpu.ALU.u_wallace._1215_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6950_  (.A1(\u_cpu.ALU.u_wallace._1209_ ),
    .A2(\u_cpu.ALU.u_wallace._1212_ ),
    .B1(\u_cpu.ALU.u_wallace._1214_ ),
    .B2(\u_cpu.ALU.u_wallace._1215_ ),
    .Y(\u_cpu.ALU.u_wallace._1216_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6951_  (.A1(\u_cpu.ALU.u_wallace._1174_ ),
    .A2(\u_cpu.ALU.u_wallace._0980_ ),
    .B1(\u_cpu.ALU.u_wallace._1207_ ),
    .C1(\u_cpu.ALU.u_wallace._1216_ ),
    .Y(\u_cpu.ALU.u_wallace._1217_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6952_  (.A1(\u_cpu.ALU.u_wallace._1178_ ),
    .A2(\u_cpu.ALU.u_wallace._1181_ ),
    .B1(\u_cpu.ALU.u_wallace._1214_ ),
    .B2(\u_cpu.ALU.u_wallace._1215_ ),
    .Y(\u_cpu.ALU.u_wallace._1218_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6953_  (.A1(\u_cpu.ALU.u_wallace._1209_ ),
    .A2(\u_cpu.ALU.u_wallace._1212_ ),
    .B1(\u_cpu.ALU.u_wallace._1203_ ),
    .C1(\u_cpu.ALU.u_wallace._1206_ ),
    .Y(\u_cpu.ALU.u_wallace._1219_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6954_  (.A1(\u_cpu.ALU.u_wallace._0923_ ),
    .A2(\u_cpu.ALU.u_wallace._0908_ ),
    .B1(\u_cpu.ALU.u_wallace._1174_ ),
    .Y(\u_cpu.ALU.u_wallace._1220_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._6955_  (.A1(\u_cpu.ALU.u_wallace._0043_ ),
    .A2(\u_cpu.ALU.u_wallace._0973_ ),
    .A3(\u_cpu.ALU.u_wallace._0967_ ),
    .B1(\u_cpu.ALU.u_wallace._0964_ ),
    .X(\u_cpu.ALU.u_wallace._1221_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._6956_  (.A1(\u_cpu.ALU.u_wallace._1218_ ),
    .A2(\u_cpu.ALU.u_wallace._1219_ ),
    .A3(\u_cpu.ALU.u_wallace._1220_ ),
    .B1(\u_cpu.ALU.u_wallace._1221_ ),
    .Y(\u_cpu.ALU.u_wallace._1222_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6957_  (.A(\u_cpu.ALU.u_wallace._1218_ ),
    .B(\u_cpu.ALU.u_wallace._1219_ ),
    .C(\u_cpu.ALU.u_wallace._1220_ ),
    .Y(\u_cpu.ALU.u_wallace._1223_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6958_  (.A(\u_cpu.ALU.u_wallace._1217_ ),
    .B(\u_cpu.ALU.u_wallace._1223_ ),
    .Y(\u_cpu.ALU.u_wallace._1225_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6959_  (.A1(\u_cpu.ALU.u_wallace._1217_ ),
    .A2(\u_cpu.ALU.u_wallace._1222_ ),
    .B1(\u_cpu.ALU.u_wallace._1225_ ),
    .B2(\u_cpu.ALU.u_wallace._1221_ ),
    .Y(\u_cpu.ALU.u_wallace._1226_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6960_  (.A(\u_cpu.ALU.u_wallace._1173_ ),
    .B(\u_cpu.ALU.u_wallace._1226_ ),
    .Y(\u_cpu.ALU.u_wallace._1227_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6961_  (.A1(\u_cpu.ALU.u_wallace._0919_ ),
    .A2(\u_cpu.ALU.u_wallace._1023_ ),
    .B1(\u_cpu.ALU.u_wallace._0921_ ),
    .Y(\u_cpu.ALU.u_wallace._1228_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6962_  (.A1(\u_cpu.ALU.u_wallace._1159_ ),
    .A2(\u_cpu.ALU.u_wallace._1164_ ),
    .B1(\u_cpu.ALU.u_wallace._1228_ ),
    .Y(\u_cpu.ALU.u_wallace._1229_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._6963_  (.A1(\u_cpu.ALU.u_wallace._1165_ ),
    .A2(\u_cpu.ALU.u_wallace._1229_ ),
    .B1_N(\u_cpu.ALU.u_wallace._1226_ ),
    .Y(\u_cpu.ALU.u_wallace._1230_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._6964_  (.A1(\u_cpu.ALU.u_wallace._0929_ ),
    .A2(\u_cpu.ALU.u_wallace._0996_ ),
    .B1(\u_cpu.ALU.u_wallace._1165_ ),
    .B2(\u_cpu.ALU.u_wallace._1227_ ),
    .C1(\u_cpu.ALU.u_wallace._1230_ ),
    .Y(\u_cpu.ALU.u_wallace._1231_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.ALU.u_wallace._6965_  (.A1(\u_cpu.ALU.u_wallace._1172_ ),
    .A2(\u_cpu.ALU.u_wallace._1170_ ),
    .A3(\u_cpu.ALU.u_wallace._1171_ ),
    .B1(\u_cpu.ALU.u_wallace._1173_ ),
    .C1(\u_cpu.ALU.u_wallace._1226_ ),
    .Y(\u_cpu.ALU.u_wallace._1232_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6966_  (.A1(\u_cpu.ALU.u_wallace._0984_ ),
    .A2(\u_cpu.ALU.u_wallace._0992_ ),
    .B1(\u_cpu.ALU.u_wallace._0986_ ),
    .Y(\u_cpu.ALU.u_wallace._1233_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6967_  (.A1(\u_cpu.ALU.u_wallace._1232_ ),
    .A2(\u_cpu.ALU.u_wallace._1230_ ),
    .B1(\u_cpu.ALU.u_wallace._1233_ ),
    .X(\u_cpu.ALU.u_wallace._1234_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._6968_  (.A(\u_cpu.ALU.u_wallace._1021_ ),
    .B(\u_cpu.ALU.u_wallace._1231_ ),
    .C(\u_cpu.ALU.u_wallace._1234_ ),
    .Y(\u_cpu.ALU.u_wallace._1236_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._6969_  (.A1(\u_cpu.ALU.u_wallace._0929_ ),
    .A2(\u_cpu.ALU.u_wallace._0996_ ),
    .B1(\u_cpu.ALU.u_wallace._1165_ ),
    .B2(\u_cpu.ALU.u_wallace._1227_ ),
    .C1(\u_cpu.ALU.u_wallace._1230_ ),
    .X(\u_cpu.ALU.u_wallace._1237_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6970_  (.A1(\u_cpu.ALU.u_wallace._1232_ ),
    .A2(\u_cpu.ALU.u_wallace._1230_ ),
    .B1(\u_cpu.ALU.u_wallace._1233_ ),
    .Y(\u_cpu.ALU.u_wallace._1238_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._6971_  (.A1(\u_cpu.ALU.u_wallace._1237_ ),
    .A2(\u_cpu.ALU.u_wallace._1238_ ),
    .B1_N(\u_cpu.ALU.u_wallace._1021_ ),
    .Y(\u_cpu.ALU.u_wallace._1239_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6972_  (.A1(\u_cpu.ALU.u_wallace._1004_ ),
    .A2(\u_cpu.ALU.u_wallace._1019_ ),
    .B1(\u_cpu.ALU.u_wallace._1236_ ),
    .C1(\u_cpu.ALU.u_wallace._1239_ ),
    .Y(\u_cpu.ALU.u_wallace._1240_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6973_  (.A1(\u_cpu.ALU.u_wallace._1006_ ),
    .A2(\u_cpu.ALU.u_wallace._1007_ ),
    .B1(\u_cpu.ALU.u_wallace._0991_ ),
    .Y(\u_cpu.ALU.u_wallace._1241_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._6974_  (.A1(\u_cpu.ALU.u_wallace._1236_ ),
    .A2(\u_cpu.ALU.u_wallace._1239_ ),
    .B1(\u_cpu.ALU.u_wallace._1241_ ),
    .X(\u_cpu.ALU.u_wallace._1242_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._6975_  (.A1(\u_cpu.ALU.u_wallace._0787_ ),
    .A2(\u_cpu.ALU.u_wallace._1013_ ),
    .B1(\u_cpu.ALU.u_wallace._1240_ ),
    .C1(\u_cpu.ALU.u_wallace._1242_ ),
    .Y(\u_cpu.ALU.u_wallace._1243_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6976_  (.A(\u_cpu.ALU.u_wallace._1003_ ),
    .B(\u_cpu.ALU.u_wallace._1008_ ),
    .Y(\u_cpu.ALU.u_wallace._1244_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._6977_  (.A1(\u_cpu.ALU.u_wallace._0784_ ),
    .A2(\u_cpu.ALU.u_wallace._0780_ ),
    .B1(\u_cpu.ALU.u_wallace._0767_ ),
    .X(\u_cpu.ALU.u_wallace._1245_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6978_  (.A1(\u_cpu.ALU.u_wallace._1244_ ),
    .A2(\u_cpu.ALU.u_wallace._1245_ ),
    .B1(\u_cpu.ALU.u_wallace._0787_ ),
    .Y(\u_cpu.ALU.u_wallace._1247_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6979_  (.A(\u_cpu.ALU.u_wallace._1240_ ),
    .B(\u_cpu.ALU.u_wallace._1242_ ),
    .Y(\u_cpu.ALU.u_wallace._1248_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6980_  (.A1(\u_cpu.ALU.u_wallace._1012_ ),
    .A2(\u_cpu.ALU.u_wallace._1247_ ),
    .B1(\u_cpu.ALU.u_wallace._1248_ ),
    .Y(\u_cpu.ALU.u_wallace._1249_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6981_  (.A1(\u_cpu.ALU.u_wallace._1012_ ),
    .A2(\u_cpu.ALU.u_wallace._1243_ ),
    .B1(\u_cpu.ALU.u_wallace._1249_ ),
    .Y(\u_cpu.ALU.u_wallace._1250_ ));
 sky130_fd_sc_hd__nor4_2 \u_cpu.ALU.u_wallace._6982_  (.A(\u_cpu.ALU.u_wallace._1013_ ),
    .B(\u_cpu.ALU.u_wallace._0593_ ),
    .C(\u_cpu.ALU.u_wallace._1012_ ),
    .D(\u_cpu.ALU.u_wallace._0793_ ),
    .Y(\u_cpu.ALU.u_wallace._1251_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6983_  (.A1(\u_cpu.ALU.u_wallace._1015_ ),
    .A2(\u_cpu.ALU.u_wallace._1018_ ),
    .B1(\u_cpu.ALU.u_wallace._1251_ ),
    .Y(\u_cpu.ALU.u_wallace._1252_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu.ALU.u_wallace._6984_  (.A(\u_cpu.ALU.u_wallace._1250_ ),
    .B(\u_cpu.ALU.u_wallace._1252_ ),
    .Y(\u_cpu.ALU.Product_Wallace[19] ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._6985_  (.A1(\u_cpu.ALU.u_wallace._1236_ ),
    .A2(\u_cpu.ALU.u_wallace._1239_ ),
    .B1(\u_cpu.ALU.u_wallace._1241_ ),
    .Y(\u_cpu.ALU.u_wallace._1253_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6986_  (.A1(\u_cpu.ALU.u_wallace._1020_ ),
    .A2(\u_cpu.ALU.u_wallace._1238_ ),
    .B1(\u_cpu.ALU.u_wallace._1231_ ),
    .Y(\u_cpu.ALU.u_wallace._1254_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._6987_  (.A(\u_cpu.ALU.u_wallace._1217_ ),
    .Y(\u_cpu.ALU.u_wallace._1255_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._6988_  (.A1(\u_cpu.ALU.u_wallace._1228_ ),
    .A2(\u_cpu.ALU.u_wallace._1159_ ),
    .A3(\u_cpu.ALU.u_wallace._1164_ ),
    .B1(\u_cpu.ALU.u_wallace._1173_ ),
    .B2(\u_cpu.ALU.u_wallace._1226_ ),
    .X(\u_cpu.ALU.u_wallace._1257_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6989_  (.A1(\u_cpu.ALU.u_wallace._1117_ ),
    .A2(\u_cpu.ALU.u_wallace._1113_ ),
    .B1(\u_cpu.ALU.u_wallace._1099_ ),
    .Y(\u_cpu.ALU.u_wallace._1258_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6990_  (.A(\u_cpu.ALU.u_wallace._0742_ ),
    .B(\u_cpu.ALU.u_wallace._1073_ ),
    .Y(\u_cpu.ALU.u_wallace._1259_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._6991_  (.A1(\u_cpu.ALU.u_wallace._1158_ ),
    .A2(\u_cpu.ALU.u_wallace._0545_ ),
    .A3(\u_cpu.ALU.u_wallace._0802_ ),
    .A4(\u_cpu.ALU.u_wallace._1090_ ),
    .B1(\u_cpu.ALU.u_wallace._1259_ ),
    .X(\u_cpu.ALU.u_wallace._1260_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6992_  (.A1(\u_cpu.ALU.u_wallace._0534_ ),
    .A2(\u_cpu.ALU.u_wallace._0808_ ),
    .B1(\u_cpu.ALU.u_wallace._1100_ ),
    .B2(\u_cpu.ALU.u_wallace._0775_ ),
    .Y(\u_cpu.ALU.u_wallace._1261_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._6993_  (.A(\u_cpu.ALU.u_wallace._0797_ ),
    .B(\u_cpu.ALU.u_wallace._0293_ ),
    .C(\u_cpu.ALU.u_wallace._0808_ ),
    .D(\u_cpu.ALU.u_wallace._1100_ ),
    .X(\u_cpu.ALU.u_wallace._1262_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._6994_  (.A1(\u_cpu.ALU.u_wallace._1224_ ),
    .A2(\u_cpu.ALU.u_wallace._0635_ ),
    .B1(\u_cpu.ALU.u_wallace._1261_ ),
    .B2(\u_cpu.ALU.u_wallace._1262_ ),
    .Y(\u_cpu.ALU.u_wallace._1263_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._6995_  (.A1(\u_cpu.ALU.u_wallace._1760_ ),
    .A2(\u_cpu.ALU.SrcA[14] ),
    .B1(\u_cpu.ALU.u_wallace._0628_ ),
    .B2(\u_cpu.ALU.SrcA[3] ),
    .Y(\u_cpu.ALU.u_wallace._1264_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6996_  (.A(\u_cpu.ALU.u_wallace._0064_ ),
    .B(\u_cpu.ALU.SrcA[20] ),
    .Y(\u_cpu.ALU.u_wallace._1265_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._6997_  (.A1(\u_cpu.ALU.u_wallace._4431_ ),
    .A2(\u_cpu.ALU.u_wallace._0600_ ),
    .A3(\u_cpu.ALU.u_wallace._0313_ ),
    .A4(\u_cpu.ALU.u_wallace._1102_ ),
    .B1(\u_cpu.ALU.u_wallace._1265_ ),
    .X(\u_cpu.ALU.u_wallace._1266_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._6998_  (.A(\u_cpu.ALU.u_wallace._0075_ ),
    .B(\u_cpu.ALU.u_wallace._1090_ ),
    .Y(\u_cpu.ALU.u_wallace._1268_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._6999_  (.A1(\u_cpu.ALU.u_wallace._1268_ ),
    .A2(\u_cpu.ALU.u_wallace._1093_ ),
    .B1(\u_cpu.ALU.u_wallace._1089_ ),
    .Y(\u_cpu.ALU.u_wallace._1269_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7000_  (.A(\u_cpu.ALU.SrcA[20] ),
    .X(\u_cpu.ALU.u_wallace._1270_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7001_  (.A(\u_cpu.ALU.u_wallace._1270_ ),
    .Y(\u_cpu.ALU.u_wallace._1271_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7002_  (.A(\u_cpu.ALU.u_wallace._1760_ ),
    .B(\u_cpu.ALU.SrcA[3] ),
    .C(\u_cpu.ALU.SrcA[14] ),
    .D(\u_cpu.ALU.SrcB[17] ),
    .X(\u_cpu.ALU.u_wallace._1272_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7003_  (.A1(\u_cpu.ALU.u_wallace._0634_ ),
    .A2(\u_cpu.ALU.u_wallace._1271_ ),
    .B1(\u_cpu.ALU.u_wallace._1264_ ),
    .B2(\u_cpu.ALU.u_wallace._1272_ ),
    .Y(\u_cpu.ALU.u_wallace._1273_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7004_  (.A1(\u_cpu.ALU.u_wallace._1264_ ),
    .A2(\u_cpu.ALU.u_wallace._1266_ ),
    .B1(\u_cpu.ALU.u_wallace._1269_ ),
    .C1(\u_cpu.ALU.u_wallace._1273_ ),
    .Y(\u_cpu.ALU.u_wallace._1274_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7005_  (.A(\u_cpu.ALU.u_wallace._1270_ ),
    .X(\u_cpu.ALU.u_wallace._1275_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7006_  (.A1(\u_cpu.ALU.u_wallace._3678_ ),
    .A2(\u_cpu.ALU.u_wallace._0182_ ),
    .B1(\u_cpu.ALU.u_wallace._0813_ ),
    .B2(\u_cpu.ALU.u_wallace._2549_ ),
    .X(\u_cpu.ALU.u_wallace._1276_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7007_  (.A(\u_cpu.ALU.u_wallace._4645_ ),
    .B(\u_cpu.ALU.u_wallace._2549_ ),
    .C(\u_cpu.ALU.u_wallace._0177_ ),
    .D(\u_cpu.ALU.u_wallace._0639_ ),
    .Y(\u_cpu.ALU.u_wallace._1277_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7008_  (.A1(\u_cpu.ALU.u_wallace._0873_ ),
    .A2(\u_cpu.ALU.u_wallace._1275_ ),
    .B1(\u_cpu.ALU.u_wallace._1276_ ),
    .B2(\u_cpu.ALU.u_wallace._1277_ ),
    .Y(\u_cpu.ALU.u_wallace._1279_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._7009_  (.A(\u_cpu.ALU.u_wallace._1265_ ),
    .B(\u_cpu.ALU.u_wallace._1264_ ),
    .C(\u_cpu.ALU.u_wallace._1272_ ),
    .Y(\u_cpu.ALU.u_wallace._1280_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._7010_  (.A1(\u_cpu.ALU.u_wallace._0634_ ),
    .A2(\u_cpu.ALU.u_wallace._1096_ ),
    .A3(\u_cpu.ALU.u_wallace._1093_ ),
    .B1(\u_cpu.ALU.u_wallace._1089_ ),
    .X(\u_cpu.ALU.u_wallace._1281_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7011_  (.A1(\u_cpu.ALU.u_wallace._1279_ ),
    .A2(\u_cpu.ALU.u_wallace._1280_ ),
    .B1(\u_cpu.ALU.u_wallace._1281_ ),
    .Y(\u_cpu.ALU.u_wallace._1282_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._7012_  (.A1(\u_cpu.ALU.u_wallace._1260_ ),
    .A2(\u_cpu.ALU.u_wallace._1261_ ),
    .B1(\u_cpu.ALU.u_wallace._1263_ ),
    .C1(\u_cpu.ALU.u_wallace._1274_ ),
    .D1(\u_cpu.ALU.u_wallace._1282_ ),
    .Y(\u_cpu.ALU.u_wallace._1283_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._7013_  (.A1(\u_cpu.ALU.u_wallace._1892_ ),
    .A2(\u_cpu.ALU.u_wallace._0635_ ),
    .B1(\u_cpu.ALU.u_wallace._1261_ ),
    .B2(\u_cpu.ALU.u_wallace._1262_ ),
    .X(\u_cpu.ALU.u_wallace._1284_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7014_  (.A(\u_cpu.ALU.u_wallace._4657_ ),
    .B(\u_cpu.ALU.u_wallace._4658_ ),
    .C(\u_cpu.ALU.u_wallace._1084_ ),
    .D(\u_cpu.ALU.u_wallace._1090_ ),
    .Y(\u_cpu.ALU.u_wallace._1285_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7015_  (.A(\u_cpu.ALU.u_wallace._1073_ ),
    .X(\u_cpu.ALU.u_wallace._1286_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.ALU.u_wallace._7016_  (.A_N(\u_cpu.ALU.u_wallace._1261_ ),
    .B(\u_cpu.ALU.u_wallace._1285_ ),
    .C(\u_cpu.ALU.u_wallace._0578_ ),
    .D(\u_cpu.ALU.u_wallace._1286_ ),
    .X(\u_cpu.ALU.u_wallace._1287_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7017_  (.A1(\u_cpu.ALU.u_wallace._1264_ ),
    .A2(\u_cpu.ALU.u_wallace._1266_ ),
    .B1(\u_cpu.ALU.u_wallace._1269_ ),
    .C1(\u_cpu.ALU.u_wallace._1273_ ),
    .X(\u_cpu.ALU.u_wallace._1288_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7018_  (.A(\u_cpu.ALU.u_wallace._1276_ ),
    .B(\u_cpu.ALU.u_wallace._1277_ ),
    .C(\u_cpu.ALU.u_wallace._0086_ ),
    .D(\u_cpu.ALU.u_wallace._1275_ ),
    .Y(\u_cpu.ALU.u_wallace._1290_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7019_  (.A1(\u_cpu.ALU.u_wallace._1273_ ),
    .A2(\u_cpu.ALU.u_wallace._1290_ ),
    .B1(\u_cpu.ALU.u_wallace._1269_ ),
    .Y(\u_cpu.ALU.u_wallace._1291_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7020_  (.A1(\u_cpu.ALU.u_wallace._1284_ ),
    .A2(\u_cpu.ALU.u_wallace._1287_ ),
    .B1(\u_cpu.ALU.u_wallace._1288_ ),
    .B2(\u_cpu.ALU.u_wallace._1291_ ),
    .Y(\u_cpu.ALU.u_wallace._1292_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7021_  (.A(\u_cpu.ALU.u_wallace._1258_ ),
    .B(\u_cpu.ALU.u_wallace._1283_ ),
    .C(\u_cpu.ALU.u_wallace._1292_ ),
    .Y(\u_cpu.ALU.u_wallace._1293_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._7022_  (.A1(\u_cpu.ALU.u_wallace._1261_ ),
    .A2(\u_cpu.ALU.u_wallace._1260_ ),
    .B1(\u_cpu.ALU.u_wallace._1263_ ),
    .X(\u_cpu.ALU.u_wallace._1294_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7023_  (.A1(\u_cpu.ALU.u_wallace._1288_ ),
    .A2(\u_cpu.ALU.u_wallace._1291_ ),
    .B1(\u_cpu.ALU.u_wallace._1294_ ),
    .Y(\u_cpu.ALU.u_wallace._1295_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7024_  (.A1(\u_cpu.ALU.u_wallace._1284_ ),
    .A2(\u_cpu.ALU.u_wallace._1287_ ),
    .B1(\u_cpu.ALU.u_wallace._1274_ ),
    .C1(\u_cpu.ALU.u_wallace._1282_ ),
    .Y(\u_cpu.ALU.u_wallace._1296_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._7025_  (.A1(\u_cpu.ALU.u_wallace._1268_ ),
    .A2(\u_cpu.ALU.u_wallace._1093_ ),
    .A3(\u_cpu.ALU.u_wallace._1097_ ),
    .B1(\u_cpu.ALU.u_wallace._1095_ ),
    .X(\u_cpu.ALU.u_wallace._1297_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7026_  (.A1(\u_cpu.ALU.u_wallace._1098_ ),
    .A2(\u_cpu.ALU.u_wallace._1297_ ),
    .B1(\u_cpu.ALU.u_wallace._1107_ ),
    .B2(\u_cpu.ALU.u_wallace._1143_ ),
    .Y(\u_cpu.ALU.u_wallace._1298_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7027_  (.A(\u_cpu.ALU.u_wallace._1295_ ),
    .B(\u_cpu.ALU.u_wallace._1296_ ),
    .C(\u_cpu.ALU.u_wallace._1298_ ),
    .Y(\u_cpu.ALU.u_wallace._1299_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7028_  (.A(\u_cpu.ALU.u_wallace._1123_ ),
    .B(\u_cpu.ALU.u_wallace._0475_ ),
    .C(\u_cpu.ALU.u_wallace._2626_ ),
    .Y(\u_cpu.ALU.u_wallace._1301_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7029_  (.A(\u_cpu.ALU.u_wallace._1122_ ),
    .B(\u_cpu.ALU.u_wallace._1301_ ),
    .Y(\u_cpu.ALU.u_wallace._1302_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7030_  (.A(\u_cpu.ALU.u_wallace._0479_ ),
    .B(\u_cpu.ALU.u_wallace._1914_ ),
    .C(\u_cpu.ALU.u_wallace._0630_ ),
    .D(\u_cpu.ALU.u_wallace._1084_ ),
    .X(\u_cpu.ALU.u_wallace._1303_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7031_  (.A(\u_cpu.ALU.u_wallace._1082_ ),
    .B(\u_cpu.ALU.u_wallace._1085_ ),
    .Y(\u_cpu.ALU.u_wallace._1304_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7032_  (.A1(\u_cpu.ALU.u_wallace._1541_ ),
    .A2(\u_cpu.ALU.u_wallace._0324_ ),
    .B1(\u_cpu.ALU.u_wallace._0441_ ),
    .B2(\u_cpu.ALU.u_wallace._2144_ ),
    .X(\u_cpu.ALU.u_wallace._1305_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7033_  (.A(\u_cpu.ALU.u_wallace._2571_ ),
    .B(\u_cpu.ALU.u_wallace._1497_ ),
    .C(\u_cpu.ALU.u_wallace._0332_ ),
    .D(\u_cpu.ALU.u_wallace._0448_ ),
    .Y(\u_cpu.ALU.u_wallace._1306_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7034_  (.A(\u_cpu.ALU.u_wallace._1305_ ),
    .B(\u_cpu.ALU.u_wallace._1306_ ),
    .C(\u_cpu.ALU.u_wallace._3404_ ),
    .D(\u_cpu.ALU.u_wallace._0319_ ),
    .Y(\u_cpu.ALU.u_wallace._1307_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7035_  (.A1(\u_cpu.ALU.u_wallace._1497_ ),
    .A2(\u_cpu.ALU.u_wallace._0332_ ),
    .B1(\u_cpu.ALU.u_wallace._0448_ ),
    .B2(\u_cpu.ALU.u_wallace._4467_ ),
    .Y(\u_cpu.ALU.u_wallace._1308_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7036_  (.A(\u_cpu.ALU.u_wallace._1026_ ),
    .B(\u_cpu.ALU.u_wallace._1541_ ),
    .C(\u_cpu.ALU.u_wallace._0324_ ),
    .D(\u_cpu.ALU.u_wallace._0447_ ),
    .X(\u_cpu.ALU.u_wallace._1309_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7037_  (.A1(\u_cpu.ALU.u_wallace._4470_ ),
    .A2(\u_cpu.ALU.u_wallace._0458_ ),
    .B1(\u_cpu.ALU.u_wallace._1308_ ),
    .B2(\u_cpu.ALU.u_wallace._1309_ ),
    .Y(\u_cpu.ALU.u_wallace._1310_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7038_  (.A1(\u_cpu.ALU.u_wallace._1303_ ),
    .A2(\u_cpu.ALU.u_wallace._1304_ ),
    .B1(\u_cpu.ALU.u_wallace._1307_ ),
    .C1(\u_cpu.ALU.u_wallace._1310_ ),
    .Y(\u_cpu.ALU.u_wallace._1312_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7039_  (.A1(\u_cpu.ALU.u_wallace._1086_ ),
    .A2(\u_cpu.ALU.u_wallace._1075_ ),
    .A3(\u_cpu.ALU.u_wallace._0468_ ),
    .B1(\u_cpu.ALU.u_wallace._1303_ ),
    .X(\u_cpu.ALU.u_wallace._1313_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7040_  (.A1(\u_cpu.ALU.u_wallace._1307_ ),
    .A2(\u_cpu.ALU.u_wallace._1310_ ),
    .B1(\u_cpu.ALU.u_wallace._1313_ ),
    .X(\u_cpu.ALU.u_wallace._1314_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7041_  (.A(\u_cpu.ALU.u_wallace._1302_ ),
    .B(\u_cpu.ALU.u_wallace._1312_ ),
    .C(\u_cpu.ALU.u_wallace._1314_ ),
    .X(\u_cpu.ALU.u_wallace._1315_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7042_  (.A1(\u_cpu.ALU.u_wallace._1303_ ),
    .A2(\u_cpu.ALU.u_wallace._1304_ ),
    .B1(\u_cpu.ALU.u_wallace._1307_ ),
    .C1(\u_cpu.ALU.u_wallace._1310_ ),
    .X(\u_cpu.ALU.u_wallace._1316_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7043_  (.A1(\u_cpu.ALU.u_wallace._1307_ ),
    .A2(\u_cpu.ALU.u_wallace._1310_ ),
    .B1(\u_cpu.ALU.u_wallace._1313_ ),
    .Y(\u_cpu.ALU.u_wallace._1317_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7044_  (.A1(\u_cpu.ALU.u_wallace._1316_ ),
    .A2(\u_cpu.ALU.u_wallace._1317_ ),
    .B1(\u_cpu.ALU.u_wallace._1122_ ),
    .C1(\u_cpu.ALU.u_wallace._1301_ ),
    .X(\u_cpu.ALU.u_wallace._1318_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7045_  (.A1_N(\u_cpu.ALU.u_wallace._1293_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1299_ ),
    .B1(\u_cpu.ALU.u_wallace._1315_ ),
    .B2(\u_cpu.ALU.u_wallace._1318_ ),
    .Y(\u_cpu.ALU.u_wallace._1319_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7046_  (.A1(\u_cpu.ALU.u_wallace._1316_ ),
    .A2(\u_cpu.ALU.u_wallace._1317_ ),
    .B1(\u_cpu.ALU.u_wallace._1302_ ),
    .Y(\u_cpu.ALU.u_wallace._1320_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7047_  (.A(\u_cpu.ALU.u_wallace._2056_ ),
    .Y(\u_cpu.ALU.u_wallace._1321_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7048_  (.A(\u_cpu.ALU.u_wallace._0177_ ),
    .Y(\u_cpu.ALU.u_wallace._1323_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7049_  (.A(\u_cpu.ALU.SrcA[15] ),
    .Y(\u_cpu.ALU.u_wallace._1324_ ));
 sky130_fd_sc_hd__o41a_2 \u_cpu.ALU.u_wallace._7050_  (.A1(\u_cpu.ALU.u_wallace._1037_ ),
    .A2(\u_cpu.ALU.u_wallace._1321_ ),
    .A3(\u_cpu.ALU.u_wallace._1323_ ),
    .A4(\u_cpu.ALU.u_wallace._1324_ ),
    .B1(\u_cpu.ALU.u_wallace._1301_ ),
    .X(\u_cpu.ALU.u_wallace._1325_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7051_  (.A(\u_cpu.ALU.u_wallace._1314_ ),
    .B(\u_cpu.ALU.u_wallace._1325_ ),
    .C(\u_cpu.ALU.u_wallace._1312_ ),
    .Y(\u_cpu.ALU.u_wallace._1326_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7052_  (.A(\u_cpu.ALU.u_wallace._1320_ ),
    .B(\u_cpu.ALU.u_wallace._1326_ ),
    .Y(\u_cpu.ALU.u_wallace._1327_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7053_  (.A(\u_cpu.ALU.u_wallace._1293_ ),
    .B(\u_cpu.ALU.u_wallace._1299_ ),
    .C(\u_cpu.ALU.u_wallace._1327_ ),
    .Y(\u_cpu.ALU.u_wallace._1328_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7054_  (.A1(\u_cpu.ALU.u_wallace._1144_ ),
    .A2(\u_cpu.ALU.u_wallace._1145_ ),
    .B1(\u_cpu.ALU.u_wallace._1137_ ),
    .B2(\u_cpu.ALU.u_wallace._1155_ ),
    .Y(\u_cpu.ALU.u_wallace._1329_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7055_  (.A1(\u_cpu.ALU.u_wallace._1319_ ),
    .A2(\u_cpu.ALU.u_wallace._1328_ ),
    .B1(\u_cpu.ALU.u_wallace._1329_ ),
    .Y(\u_cpu.ALU.u_wallace._1330_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7056_  (.A(\u_cpu.ALU.u_wallace._4007_ ),
    .B(\u_cpu.ALU.u_wallace._4291_ ),
    .C(\u_cpu.ALU.u_wallace._4646_ ),
    .D(\u_cpu.ALU.u_wallace._4790_ ),
    .Y(\u_cpu.ALU.u_wallace._1331_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7057_  (.A(\u_cpu.ALU.u_wallace._1331_ ),
    .B(\u_cpu.ALU.u_wallace._4609_ ),
    .C(\u_cpu.ALU.u_wallace._4551_ ),
    .Y(\u_cpu.ALU.u_wallace._1332_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7058_  (.A1(\u_cpu.ALU.u_wallace._0045_ ),
    .A2(\u_cpu.ALU.u_wallace._4797_ ),
    .B1(\u_cpu.ALU.u_wallace._4900_ ),
    .B2(\u_cpu.ALU.u_wallace._4716_ ),
    .Y(\u_cpu.ALU.u_wallace._1334_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7059_  (.A(\u_cpu.ALU.u_wallace._4567_ ),
    .B(\u_cpu.ALU.u_wallace._0041_ ),
    .Y(\u_cpu.ALU.u_wallace._1335_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7060_  (.A1(\u_cpu.ALU.u_wallace._1335_ ),
    .A2(\u_cpu.ALU.u_wallace._1028_ ),
    .B1(\u_cpu.ALU.u_wallace._1025_ ),
    .Y(\u_cpu.ALU.u_wallace._1336_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7061_  (.A1(\u_cpu.ALU.u_wallace._0045_ ),
    .A2(\u_cpu.ALU.u_wallace._4797_ ),
    .B1(\u_cpu.ALU.u_wallace._4900_ ),
    .B2(\u_cpu.ALU.u_wallace._4847_ ),
    .X(\u_cpu.ALU.u_wallace._1337_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7062_  (.A1(\u_cpu.ALU.u_wallace._4643_ ),
    .A2(\u_cpu.ALU.u_wallace._0052_ ),
    .B1(\u_cpu.ALU.u_wallace._1331_ ),
    .B2(\u_cpu.ALU.u_wallace._1337_ ),
    .X(\u_cpu.ALU.u_wallace._1338_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7063_  (.A1(\u_cpu.ALU.u_wallace._1332_ ),
    .A2(\u_cpu.ALU.u_wallace._1334_ ),
    .B1(\u_cpu.ALU.u_wallace._1336_ ),
    .C1(\u_cpu.ALU.u_wallace._1338_ ),
    .X(\u_cpu.ALU.u_wallace._1339_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._7064_  (.A1_N(\u_cpu.ALU.u_wallace._4904_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4601_ ),
    .B1(\u_cpu.ALU.u_wallace._1331_ ),
    .B2(\u_cpu.ALU.u_wallace._1337_ ),
    .Y(\u_cpu.ALU.u_wallace._1340_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7065_  (.A(\u_cpu.ALU.u_wallace._1334_ ),
    .B(\u_cpu.ALU.u_wallace._1332_ ),
    .Y(\u_cpu.ALU.u_wallace._1341_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._7066_  (.A1(\u_cpu.ALU.u_wallace._1335_ ),
    .A2(\u_cpu.ALU.u_wallace._1028_ ),
    .B1(\u_cpu.ALU.u_wallace._1025_ ),
    .X(\u_cpu.ALU.u_wallace._1342_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7067_  (.A1(\u_cpu.ALU.u_wallace._1340_ ),
    .A2(\u_cpu.ALU.u_wallace._1341_ ),
    .B1(\u_cpu.ALU.u_wallace._1342_ ),
    .Y(\u_cpu.ALU.u_wallace._1343_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7068_  (.A1(\u_cpu.ALU.u_wallace._4412_ ),
    .A2(\u_cpu.ALU.u_wallace._0364_ ),
    .B1(\u_cpu.ALU.u_wallace._0365_ ),
    .B2(\u_cpu.ALU.u_wallace._3689_ ),
    .X(\u_cpu.ALU.u_wallace._1345_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7069_  (.A(\u_cpu.ALU.u_wallace._4561_ ),
    .B(\u_cpu.ALU.u_wallace._4412_ ),
    .C(\u_cpu.ALU.u_wallace._0364_ ),
    .D(\u_cpu.ALU.u_wallace._0365_ ),
    .Y(\u_cpu.ALU.u_wallace._1346_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7070_  (.A(\u_cpu.ALU.u_wallace._2725_ ),
    .B(\u_cpu.ALU.SrcB[13] ),
    .Y(\u_cpu.ALU.u_wallace._1347_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7071_  (.A1(\u_cpu.ALU.u_wallace._1345_ ),
    .A2(\u_cpu.ALU.u_wallace._1346_ ),
    .B1(\u_cpu.ALU.u_wallace._1347_ ),
    .X(\u_cpu.ALU.u_wallace._1348_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7072_  (.A1(\u_cpu.ALU.u_wallace._0203_ ),
    .A2(\u_cpu.ALU.u_wallace._0036_ ),
    .B1(\u_cpu.ALU.u_wallace._1345_ ),
    .C1(\u_cpu.ALU.u_wallace._1346_ ),
    .Y(\u_cpu.ALU.u_wallace._1349_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7073_  (.A(\u_cpu.ALU.u_wallace._1348_ ),
    .B(\u_cpu.ALU.u_wallace._1349_ ),
    .Y(\u_cpu.ALU.u_wallace._1350_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7074_  (.A(\u_cpu.ALU.u_wallace._1343_ ),
    .B(\u_cpu.ALU.u_wallace._1350_ ),
    .Y(\u_cpu.ALU.u_wallace._1351_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7075_  (.A1(\u_cpu.ALU.u_wallace._1332_ ),
    .A2(\u_cpu.ALU.u_wallace._1334_ ),
    .B1(\u_cpu.ALU.u_wallace._1336_ ),
    .C1(\u_cpu.ALU.u_wallace._1338_ ),
    .Y(\u_cpu.ALU.u_wallace._1352_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU.u_wallace._7076_  (.A1_N(\u_cpu.ALU.u_wallace._1345_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1346_ ),
    .B1(\u_cpu.ALU.u_wallace._0203_ ),
    .B2(\u_cpu.ALU.u_wallace._0124_ ),
    .X(\u_cpu.ALU.u_wallace._1353_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7077_  (.A(\u_cpu.ALU.u_wallace._1345_ ),
    .B(\u_cpu.ALU.u_wallace._1346_ ),
    .C(\u_cpu.ALU.u_wallace._4698_ ),
    .D(\u_cpu.ALU.u_wallace._0034_ ),
    .X(\u_cpu.ALU.u_wallace._1354_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7078_  (.A1_N(\u_cpu.ALU.u_wallace._1352_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1343_ ),
    .B1(\u_cpu.ALU.u_wallace._1353_ ),
    .B2(\u_cpu.ALU.u_wallace._1354_ ),
    .Y(\u_cpu.ALU.u_wallace._1356_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7079_  (.A1(\u_cpu.ALU.u_wallace._1339_ ),
    .A2(\u_cpu.ALU.u_wallace._1351_ ),
    .B1(\u_cpu.ALU.u_wallace._1356_ ),
    .Y(\u_cpu.ALU.u_wallace._1357_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._7080_  (.A1(\u_cpu.ALU.u_wallace._1134_ ),
    .A2(\u_cpu.ALU.u_wallace._1133_ ),
    .B1(\u_cpu.ALU.u_wallace._1139_ ),
    .X(\u_cpu.ALU.u_wallace._1358_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.ALU.u_wallace._7081_  (.A1(\u_cpu.ALU.u_wallace._1040_ ),
    .A2(\u_cpu.ALU.u_wallace._1043_ ),
    .A3(\u_cpu.ALU.u_wallace._1045_ ),
    .B1(\u_cpu.ALU.u_wallace._1051_ ),
    .B2(\u_cpu.ALU.u_wallace._1064_ ),
    .X(\u_cpu.ALU.u_wallace._1359_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7082_  (.A1(\u_cpu.ALU.u_wallace._1357_ ),
    .A2(\u_cpu.ALU.u_wallace._1358_ ),
    .B1(\u_cpu.ALU.u_wallace._1359_ ),
    .Y(\u_cpu.ALU.u_wallace._1360_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU.u_wallace._7083_  (.A1(\u_cpu.ALU.u_wallace._1342_ ),
    .A2(\u_cpu.ALU.u_wallace._1340_ ),
    .A3(\u_cpu.ALU.u_wallace._1341_ ),
    .B1(\u_cpu.ALU.u_wallace._1350_ ),
    .C1(\u_cpu.ALU.u_wallace._1343_ ),
    .X(\u_cpu.ALU.u_wallace._1361_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7084_  (.A1(\u_cpu.ALU.u_wallace._1352_ ),
    .A2(\u_cpu.ALU.u_wallace._1343_ ),
    .B1(\u_cpu.ALU.u_wallace._1350_ ),
    .Y(\u_cpu.ALU.u_wallace._1362_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._7085_  (.A1(\u_cpu.ALU.u_wallace._1139_ ),
    .A2(\u_cpu.ALU.u_wallace._1132_ ),
    .B1(\u_cpu.ALU.u_wallace._1361_ ),
    .C1(\u_cpu.ALU.u_wallace._1362_ ),
    .X(\u_cpu.ALU.u_wallace._1363_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7086_  (.A1(\u_cpu.ALU.u_wallace._1134_ ),
    .A2(\u_cpu.ALU.u_wallace._1133_ ),
    .B1(\u_cpu.ALU.u_wallace._1139_ ),
    .Y(\u_cpu.ALU.u_wallace._1364_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7087_  (.A(\u_cpu.ALU.u_wallace._1364_ ),
    .B(\u_cpu.ALU.u_wallace._1356_ ),
    .Y(\u_cpu.ALU.u_wallace._1365_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7088_  (.A1(\u_cpu.ALU.u_wallace._1361_ ),
    .A2(\u_cpu.ALU.u_wallace._1362_ ),
    .B1(\u_cpu.ALU.u_wallace._1358_ ),
    .Y(\u_cpu.ALU.u_wallace._1367_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7089_  (.A1(\u_cpu.ALU.u_wallace._1361_ ),
    .A2(\u_cpu.ALU.u_wallace._1365_ ),
    .B1(\u_cpu.ALU.u_wallace._1367_ ),
    .Y(\u_cpu.ALU.u_wallace._1368_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7090_  (.A1(\u_cpu.ALU.u_wallace._1360_ ),
    .A2(\u_cpu.ALU.u_wallace._1363_ ),
    .B1(\u_cpu.ALU.u_wallace._1359_ ),
    .B2(\u_cpu.ALU.u_wallace._1368_ ),
    .Y(\u_cpu.ALU.u_wallace._1369_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7091_  (.A(\u_cpu.ALU.u_wallace._1258_ ),
    .B(\u_cpu.ALU.u_wallace._1283_ ),
    .C(\u_cpu.ALU.u_wallace._1292_ ),
    .X(\u_cpu.ALU.u_wallace._1370_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7092_  (.A(\u_cpu.ALU.u_wallace._1299_ ),
    .B(\u_cpu.ALU.u_wallace._1327_ ),
    .Y(\u_cpu.ALU.u_wallace._1371_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7093_  (.A1(\u_cpu.ALU.u_wallace._1370_ ),
    .A2(\u_cpu.ALU.u_wallace._1371_ ),
    .B1(\u_cpu.ALU.u_wallace._1319_ ),
    .C1(\u_cpu.ALU.u_wallace._1329_ ),
    .Y(\u_cpu.ALU.u_wallace._1372_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7094_  (.A(\u_cpu.ALU.u_wallace._1369_ ),
    .B(\u_cpu.ALU.u_wallace._1372_ ),
    .Y(\u_cpu.ALU.u_wallace._1373_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7095_  (.A1(\u_cpu.ALU.u_wallace._1029_ ),
    .A2(\u_cpu.ALU.u_wallace._1063_ ),
    .A3(\u_cpu.ALU.u_wallace._1031_ ),
    .B1(\u_cpu.ALU.u_wallace._1041_ ),
    .X(\u_cpu.ALU.u_wallace._1374_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7096_  (.A1(\u_cpu.ALU.u_wallace._1363_ ),
    .A2(\u_cpu.ALU.u_wallace._1367_ ),
    .B1(\u_cpu.ALU.u_wallace._1374_ ),
    .Y(\u_cpu.ALU.u_wallace._1375_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._7097_  (.A1(\u_cpu.ALU.u_wallace._1060_ ),
    .A2(\u_cpu.ALU.u_wallace._1041_ ),
    .B1(\u_cpu.ALU.u_wallace._1361_ ),
    .B2(\u_cpu.ALU.u_wallace._1365_ ),
    .C1(\u_cpu.ALU.u_wallace._1367_ ),
    .X(\u_cpu.ALU.u_wallace._1376_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7098_  (.A1(\u_cpu.ALU.u_wallace._1370_ ),
    .A2(\u_cpu.ALU.u_wallace._1371_ ),
    .B1(\u_cpu.ALU.u_wallace._1319_ ),
    .C1(\u_cpu.ALU.u_wallace._1329_ ),
    .X(\u_cpu.ALU.u_wallace._1378_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7099_  (.A1(\u_cpu.ALU.u_wallace._1375_ ),
    .A2(\u_cpu.ALU.u_wallace._1376_ ),
    .B1(\u_cpu.ALU.u_wallace._1330_ ),
    .B2(\u_cpu.ALU.u_wallace._1378_ ),
    .Y(\u_cpu.ALU.u_wallace._1379_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7100_  (.A1(\u_cpu.ALU.u_wallace._1154_ ),
    .A2(\u_cpu.ALU.u_wallace._1108_ ),
    .A3(\u_cpu.ALU.u_wallace._1115_ ),
    .B1(\u_cpu.ALU.u_wallace._1152_ ),
    .X(\u_cpu.ALU.u_wallace._1380_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._7101_  (.A1(\u_cpu.ALU.u_wallace._1168_ ),
    .A2(\u_cpu.ALU.u_wallace._1380_ ),
    .A3(\u_cpu.ALU.u_wallace._1156_ ),
    .B1(\u_cpu.ALU.u_wallace._1150_ ),
    .B2(\u_cpu.ALU.u_wallace._1071_ ),
    .X(\u_cpu.ALU.u_wallace._1381_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7102_  (.A1(\u_cpu.ALU.u_wallace._1330_ ),
    .A2(\u_cpu.ALU.u_wallace._1373_ ),
    .B1(\u_cpu.ALU.u_wallace._1379_ ),
    .C1(\u_cpu.ALU.u_wallace._1381_ ),
    .X(\u_cpu.ALU.u_wallace._1382_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._7103_  (.A_N(\u_cpu.ALU.u_wallace._1330_ ),
    .B(\u_cpu.ALU.u_wallace._1372_ ),
    .C(\u_cpu.ALU.u_wallace._1369_ ),
    .Y(\u_cpu.ALU.u_wallace._1383_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7104_  (.A1(\u_cpu.ALU.u_wallace._1383_ ),
    .A2(\u_cpu.ALU.u_wallace._1379_ ),
    .B1(\u_cpu.ALU.u_wallace._1381_ ),
    .Y(\u_cpu.ALU.u_wallace._1384_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.ALU.u_wallace._7105_  (.A1_N(\u_cpu.ALU.u_wallace._1061_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1066_ ),
    .B1(\u_cpu.ALU.u_wallace._1067_ ),
    .B2(\u_cpu.ALU.u_wallace._1162_ ),
    .X(\u_cpu.ALU.u_wallace._1385_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7106_  (.A(\u_cpu.ALU.SrcB[20] ),
    .X(\u_cpu.ALU.u_wallace._1386_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7107_  (.A(\u_cpu.ALU.SrcB[18] ),
    .X(\u_cpu.ALU.u_wallace._1387_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7108_  (.A(\u_cpu.ALU.u_wallace._1410_ ),
    .B(\u_cpu.ALU.u_wallace._0731_ ),
    .C(\u_cpu.ALU.u_wallace._1387_ ),
    .D(\u_cpu.ALU.u_wallace._1175_ ),
    .Y(\u_cpu.ALU.u_wallace._1389_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7109_  (.A1(\u_cpu.ALU.u_wallace._0348_ ),
    .A2(\u_cpu.ALU.u_wallace._0957_ ),
    .B1(\u_cpu.ALU.u_wallace._1210_ ),
    .B2(\u_cpu.ALU.u_wallace._0250_ ),
    .X(\u_cpu.ALU.u_wallace._1390_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7110_  (.A1(\u_cpu.ALU.u_wallace._0446_ ),
    .A2(\u_cpu.ALU.u_wallace._1386_ ),
    .B1(\u_cpu.ALU.u_wallace._1389_ ),
    .B2(\u_cpu.ALU.u_wallace._1390_ ),
    .X(\u_cpu.ALU.u_wallace._1391_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7111_  (.A(\u_cpu.ALU.SrcB[20] ),
    .X(\u_cpu.ALU.u_wallace._1392_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7112_  (.A(\u_cpu.ALU.u_wallace._1390_ ),
    .B(\u_cpu.ALU.u_wallace._1392_ ),
    .C(\u_cpu.ALU.u_wallace._0108_ ),
    .D(\u_cpu.ALU.u_wallace._1389_ ),
    .Y(\u_cpu.ALU.u_wallace._1393_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7113_  (.A(\u_cpu.ALU.u_wallace._1391_ ),
    .B(\u_cpu.ALU.u_wallace._1209_ ),
    .C(\u_cpu.ALU.u_wallace._1393_ ),
    .X(\u_cpu.ALU.u_wallace._1394_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.ALU.u_wallace._7114_  (.A1_N(\u_cpu.ALU.u_wallace._1179_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1177_ ),
    .B1(\u_cpu.ALU.u_wallace._1393_ ),
    .B2(\u_cpu.ALU.u_wallace._1391_ ),
    .X(\u_cpu.ALU.u_wallace._1395_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.ALU.u_wallace._7115_  (.A(\u_cpu.ALU.u_wallace._1394_ ),
    .B_N(\u_cpu.ALU.u_wallace._1395_ ),
    .X(\u_cpu.ALU.u_wallace._1396_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7116_  (.A(\u_cpu.ALU.u_wallace._4561_ ),
    .B(\u_cpu.ALU.u_wallace._4447_ ),
    .C(\u_cpu.ALU.u_wallace._0364_ ),
    .D(\u_cpu.ALU.u_wallace._4841_ ),
    .X(\u_cpu.ALU.u_wallace._1397_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7117_  (.A(\u_cpu.ALU.u_wallace._1035_ ),
    .B(\u_cpu.ALU.u_wallace._1047_ ),
    .Y(\u_cpu.ALU.u_wallace._1398_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7118_  (.A1(\u_cpu.ALU.u_wallace._2834_ ),
    .A2(\u_cpu.ALU.u_wallace._0120_ ),
    .B1(\u_cpu.ALU.u_wallace._0732_ ),
    .B2(\u_cpu.ALU.u_wallace._2955_ ),
    .Y(\u_cpu.ALU.u_wallace._1400_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7119_  (.A(\u_cpu.ALU.u_wallace._3832_ ),
    .B(\u_cpu.ALU.u_wallace._1125_ ),
    .C(\u_cpu.ALU.u_wallace._0546_ ),
    .D(\u_cpu.ALU.u_wallace._0547_ ),
    .Y(\u_cpu.ALU.u_wallace._1401_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._7120_  (.A_N(\u_cpu.ALU.u_wallace._1400_ ),
    .B(\u_cpu.ALU.u_wallace._1401_ ),
    .C(\u_cpu.ALU.u_wallace._2933_ ),
    .D(\u_cpu.ALU.u_wallace._0735_ ),
    .Y(\u_cpu.ALU.u_wallace._1402_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7121_  (.A(\u_cpu.ALU.u_wallace._1793_ ),
    .B(\u_cpu.ALU.u_wallace._2955_ ),
    .C(\u_cpu.ALU.u_wallace._0120_ ),
    .D(\u_cpu.ALU.u_wallace._0728_ ),
    .X(\u_cpu.ALU.u_wallace._1403_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7122_  (.A1(\u_cpu.ALU.u_wallace._0939_ ),
    .A2(\u_cpu.ALU.u_wallace._0941_ ),
    .B1(\u_cpu.ALU.u_wallace._1400_ ),
    .B2(\u_cpu.ALU.u_wallace._1403_ ),
    .Y(\u_cpu.ALU.u_wallace._1404_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7123_  (.A1(\u_cpu.ALU.u_wallace._1397_ ),
    .A2(\u_cpu.ALU.u_wallace._1398_ ),
    .B1(\u_cpu.ALU.u_wallace._1402_ ),
    .C1(\u_cpu.ALU.u_wallace._1404_ ),
    .X(\u_cpu.ALU.u_wallace._1405_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7124_  (.A1(\u_cpu.ALU.u_wallace._1184_ ),
    .A2(\u_cpu.ALU.u_wallace._0551_ ),
    .A3(\u_cpu.ALU.u_wallace._4541_ ),
    .B1(\u_cpu.ALU.u_wallace._1188_ ),
    .X(\u_cpu.ALU.u_wallace._1406_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7125_  (.A1(\u_cpu.ALU.u_wallace._1034_ ),
    .A2(\u_cpu.ALU.u_wallace._0363_ ),
    .A3(\u_cpu.ALU.u_wallace._4452_ ),
    .B1(\u_cpu.ALU.u_wallace._1397_ ),
    .X(\u_cpu.ALU.u_wallace._1407_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7126_  (.A1(\u_cpu.ALU.u_wallace._1402_ ),
    .A2(\u_cpu.ALU.u_wallace._1404_ ),
    .B1(\u_cpu.ALU.u_wallace._1407_ ),
    .X(\u_cpu.ALU.u_wallace._1408_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7127_  (.A(\u_cpu.ALU.u_wallace._1406_ ),
    .B(\u_cpu.ALU.u_wallace._1408_ ),
    .Y(\u_cpu.ALU.u_wallace._1409_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7128_  (.A1(\u_cpu.ALU.u_wallace._1186_ ),
    .A2(\u_cpu.ALU.u_wallace._1204_ ),
    .B1(\u_cpu.ALU.u_wallace._1193_ ),
    .Y(\u_cpu.ALU.u_wallace._1411_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7129_  (.A1(\u_cpu.ALU.u_wallace._1402_ ),
    .A2(\u_cpu.ALU.u_wallace._1404_ ),
    .B1(\u_cpu.ALU.u_wallace._1407_ ),
    .Y(\u_cpu.ALU.u_wallace._1412_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._7130_  (.A1(\u_cpu.ALU.u_wallace._0621_ ),
    .A2(\u_cpu.ALU.u_wallace._0554_ ),
    .A3(\u_cpu.ALU.u_wallace._1187_ ),
    .B1(\u_cpu.ALU.u_wallace._1185_ ),
    .X(\u_cpu.ALU.u_wallace._1413_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7131_  (.A1(\u_cpu.ALU.u_wallace._1405_ ),
    .A2(\u_cpu.ALU.u_wallace._1412_ ),
    .B1(\u_cpu.ALU.u_wallace._1413_ ),
    .Y(\u_cpu.ALU.u_wallace._1414_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._7132_  (.A1(\u_cpu.ALU.u_wallace._1405_ ),
    .A2(\u_cpu.ALU.u_wallace._1409_ ),
    .B1(\u_cpu.ALU.u_wallace._1196_ ),
    .B2(\u_cpu.ALU.u_wallace._1411_ ),
    .C1(\u_cpu.ALU.u_wallace._1414_ ),
    .Y(\u_cpu.ALU.u_wallace._1415_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7133_  (.A1(\u_cpu.ALU.u_wallace._1397_ ),
    .A2(\u_cpu.ALU.u_wallace._1398_ ),
    .B1(\u_cpu.ALU.u_wallace._1402_ ),
    .C1(\u_cpu.ALU.u_wallace._1404_ ),
    .Y(\u_cpu.ALU.u_wallace._1416_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7134_  (.A(\u_cpu.ALU.u_wallace._1406_ ),
    .B(\u_cpu.ALU.u_wallace._1416_ ),
    .C(\u_cpu.ALU.u_wallace._1408_ ),
    .Y(\u_cpu.ALU.u_wallace._1417_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7135_  (.A1(\u_cpu.ALU.u_wallace._1183_ ),
    .A2(\u_cpu.ALU.u_wallace._1190_ ),
    .B1(\u_cpu.ALU.u_wallace._1193_ ),
    .Y(\u_cpu.ALU.u_wallace._1418_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7136_  (.A1(\u_cpu.ALU.u_wallace._1417_ ),
    .A2(\u_cpu.ALU.u_wallace._1414_ ),
    .B1(\u_cpu.ALU.u_wallace._1418_ ),
    .X(\u_cpu.ALU.u_wallace._1419_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._7137_  (.A_N(\u_cpu.ALU.u_wallace._1396_ ),
    .B(\u_cpu.ALU.u_wallace._1415_ ),
    .C(\u_cpu.ALU.u_wallace._1419_ ),
    .Y(\u_cpu.ALU.u_wallace._1420_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7138_  (.A(\u_cpu.ALU.u_wallace._1393_ ),
    .B(\u_cpu.ALU.u_wallace._1391_ ),
    .Y(\u_cpu.ALU.u_wallace._1422_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._7139_  (.A1(\u_cpu.ALU.u_wallace._0043_ ),
    .A2(\u_cpu.ALU.u_wallace._1211_ ),
    .A3(\u_cpu.ALU.u_wallace._1179_ ),
    .B1(\u_cpu.ALU.u_wallace._1422_ ),
    .X(\u_cpu.ALU.u_wallace._1423_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7140_  (.A1(\u_cpu.ALU.u_wallace._1405_ ),
    .A2(\u_cpu.ALU.u_wallace._1409_ ),
    .B1(\u_cpu.ALU.u_wallace._1414_ ),
    .C1(\u_cpu.ALU.u_wallace._1418_ ),
    .X(\u_cpu.ALU.u_wallace._1424_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7141_  (.A1(\u_cpu.ALU.u_wallace._1417_ ),
    .A2(\u_cpu.ALU.u_wallace._1414_ ),
    .B1(\u_cpu.ALU.u_wallace._1418_ ),
    .Y(\u_cpu.ALU.u_wallace._1425_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7142_  (.A1(\u_cpu.ALU.u_wallace._1394_ ),
    .A2(\u_cpu.ALU.u_wallace._1423_ ),
    .B1(\u_cpu.ALU.u_wallace._1424_ ),
    .B2(\u_cpu.ALU.u_wallace._1425_ ),
    .Y(\u_cpu.ALU.u_wallace._1426_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7143_  (.A(\u_cpu.ALU.u_wallace._1385_ ),
    .B(\u_cpu.ALU.u_wallace._1420_ ),
    .C(\u_cpu.ALU.u_wallace._1426_ ),
    .Y(\u_cpu.ALU.u_wallace._1427_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7144_  (.A(\u_cpu.ALU.u_wallace._1427_ ),
    .Y(\u_cpu.ALU.u_wallace._1428_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU.u_wallace._7145_  (.A1_N(\u_cpu.ALU.u_wallace._1162_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1067_ ),
    .B1(\u_cpu.ALU.u_wallace._1066_ ),
    .B2(\u_cpu.ALU.u_wallace._1061_ ),
    .X(\u_cpu.ALU.u_wallace._1429_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._7146_  (.A1(\u_cpu.ALU.u_wallace._1424_ ),
    .A2(\u_cpu.ALU.u_wallace._1425_ ),
    .B1_N(\u_cpu.ALU.u_wallace._1396_ ),
    .Y(\u_cpu.ALU.u_wallace._1430_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7147_  (.A1(\u_cpu.ALU.u_wallace._1394_ ),
    .A2(\u_cpu.ALU.u_wallace._1423_ ),
    .B1(\u_cpu.ALU.u_wallace._1415_ ),
    .C1(\u_cpu.ALU.u_wallace._1419_ ),
    .Y(\u_cpu.ALU.u_wallace._1431_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._7148_  (.A1(\u_cpu.ALU.u_wallace._1209_ ),
    .A2(\u_cpu.ALU.u_wallace._1212_ ),
    .A3(\u_cpu.ALU.u_wallace._1215_ ),
    .B1(\u_cpu.ALU.u_wallace._1203_ ),
    .X(\u_cpu.ALU.u_wallace._1433_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7149_  (.A1(\u_cpu.ALU.u_wallace._1429_ ),
    .A2(\u_cpu.ALU.u_wallace._1430_ ),
    .A3(\u_cpu.ALU.u_wallace._1431_ ),
    .B1(\u_cpu.ALU.u_wallace._1433_ ),
    .X(\u_cpu.ALU.u_wallace._1434_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7150_  (.A1(\u_cpu.ALU.u_wallace._1396_ ),
    .A2(\u_cpu.ALU.u_wallace._1425_ ),
    .B1(\u_cpu.ALU.u_wallace._1415_ ),
    .Y(\u_cpu.ALU.u_wallace._1435_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7151_  (.A1(\u_cpu.ALU.u_wallace._1425_ ),
    .A2(\u_cpu.ALU.u_wallace._1435_ ),
    .B1(\u_cpu.ALU.u_wallace._1430_ ),
    .C1(\u_cpu.ALU.u_wallace._1429_ ),
    .Y(\u_cpu.ALU.u_wallace._1436_ ));
 sky130_fd_sc_hd__a21bo_2 \u_cpu.ALU.u_wallace._7152_  (.A1(\u_cpu.ALU.u_wallace._1436_ ),
    .A2(\u_cpu.ALU.u_wallace._1427_ ),
    .B1_N(\u_cpu.ALU.u_wallace._1433_ ),
    .X(\u_cpu.ALU.u_wallace._1437_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7153_  (.A1(\u_cpu.ALU.u_wallace._1428_ ),
    .A2(\u_cpu.ALU.u_wallace._1434_ ),
    .B1(\u_cpu.ALU.u_wallace._1437_ ),
    .Y(\u_cpu.ALU.u_wallace._1438_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7154_  (.A1(\u_cpu.ALU.u_wallace._1382_ ),
    .A2(\u_cpu.ALU.u_wallace._1384_ ),
    .B1(\u_cpu.ALU.u_wallace._1438_ ),
    .Y(\u_cpu.ALU.u_wallace._1439_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7155_  (.A1(\u_cpu.ALU.u_wallace._1330_ ),
    .A2(\u_cpu.ALU.u_wallace._1373_ ),
    .B1(\u_cpu.ALU.u_wallace._1379_ ),
    .C1(\u_cpu.ALU.u_wallace._1381_ ),
    .Y(\u_cpu.ALU.u_wallace._1440_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7156_  (.A1(\u_cpu.ALU.u_wallace._1330_ ),
    .A2(\u_cpu.ALU.u_wallace._1373_ ),
    .B1(\u_cpu.ALU.u_wallace._1379_ ),
    .Y(\u_cpu.ALU.u_wallace._1441_ ));
 sky130_fd_sc_hd__a32oi_2 \u_cpu.ALU.u_wallace._7157_  (.A1(\u_cpu.ALU.u_wallace._1168_ ),
    .A2(\u_cpu.ALU.u_wallace._1380_ ),
    .A3(\u_cpu.ALU.u_wallace._1156_ ),
    .B1(\u_cpu.ALU.u_wallace._1150_ ),
    .B2(\u_cpu.ALU.u_wallace._1071_ ),
    .Y(\u_cpu.ALU.u_wallace._1442_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7158_  (.A(\u_cpu.ALU.u_wallace._1441_ ),
    .B(\u_cpu.ALU.u_wallace._1442_ ),
    .Y(\u_cpu.ALU.u_wallace._1444_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._7159_  (.A1(\u_cpu.ALU.u_wallace._1434_ ),
    .A2(\u_cpu.ALU.u_wallace._1428_ ),
    .B1(\u_cpu.ALU.u_wallace._1437_ ),
    .C1(\u_cpu.ALU.u_wallace._1440_ ),
    .D1(\u_cpu.ALU.u_wallace._1444_ ),
    .Y(\u_cpu.ALU.u_wallace._1445_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7160_  (.A(\u_cpu.ALU.u_wallace._1257_ ),
    .B(\u_cpu.ALU.u_wallace._1439_ ),
    .C(\u_cpu.ALU.u_wallace._1445_ ),
    .Y(\u_cpu.ALU.u_wallace._1446_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._7161_  (.A1(\u_cpu.ALU.u_wallace._1436_ ),
    .A2(\u_cpu.ALU.u_wallace._1427_ ),
    .B1_N(\u_cpu.ALU.u_wallace._1433_ ),
    .Y(\u_cpu.ALU.u_wallace._1447_ ));
 sky130_fd_sc_hd__and3b_2 \u_cpu.ALU.u_wallace._7162_  (.A_N(\u_cpu.ALU.u_wallace._1433_ ),
    .B(\u_cpu.ALU.u_wallace._1436_ ),
    .C(\u_cpu.ALU.u_wallace._1427_ ),
    .X(\u_cpu.ALU.u_wallace._1448_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._7163_  (.A1_N(\u_cpu.ALU.u_wallace._1447_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1448_ ),
    .B1(\u_cpu.ALU.u_wallace._1440_ ),
    .B2(\u_cpu.ALU.u_wallace._1444_ ),
    .Y(\u_cpu.ALU.u_wallace._1449_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._7164_  (.A1(\u_cpu.ALU.u_wallace._1434_ ),
    .A2(\u_cpu.ALU.u_wallace._1428_ ),
    .B1(\u_cpu.ALU.u_wallace._1437_ ),
    .C1(\u_cpu.ALU.u_wallace._1440_ ),
    .D1(\u_cpu.ALU.u_wallace._1444_ ),
    .X(\u_cpu.ALU.u_wallace._1450_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._7165_  (.A1(\u_cpu.ALU.u_wallace._1172_ ),
    .A2(\u_cpu.ALU.u_wallace._1170_ ),
    .A3(\u_cpu.ALU.u_wallace._1171_ ),
    .B1(\u_cpu.ALU.u_wallace._1227_ ),
    .X(\u_cpu.ALU.u_wallace._1451_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7166_  (.A1(\u_cpu.ALU.u_wallace._1449_ ),
    .A2(\u_cpu.ALU.u_wallace._1450_ ),
    .B1(\u_cpu.ALU.u_wallace._1451_ ),
    .Y(\u_cpu.ALU.u_wallace._1452_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7167_  (.A1(\u_cpu.ALU.u_wallace._1255_ ),
    .A2(\u_cpu.ALU.u_wallace._1222_ ),
    .B1(\u_cpu.ALU.u_wallace._1446_ ),
    .C1(\u_cpu.ALU.u_wallace._1452_ ),
    .Y(\u_cpu.ALU.u_wallace._1453_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7168_  (.A(\u_cpu.ALU.u_wallace._1255_ ),
    .B(\u_cpu.ALU.u_wallace._1222_ ),
    .Y(\u_cpu.ALU.u_wallace._1455_ ));
 sky130_fd_sc_hd__a21bo_2 \u_cpu.ALU.u_wallace._7169_  (.A1(\u_cpu.ALU.u_wallace._1446_ ),
    .A2(\u_cpu.ALU.u_wallace._1452_ ),
    .B1_N(\u_cpu.ALU.u_wallace._1455_ ),
    .X(\u_cpu.ALU.u_wallace._1456_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7170_  (.A(\u_cpu.ALU.u_wallace._1254_ ),
    .B(\u_cpu.ALU.u_wallace._1453_ ),
    .C(\u_cpu.ALU.u_wallace._1456_ ),
    .Y(\u_cpu.ALU.u_wallace._1457_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7171_  (.A1(\u_cpu.ALU.u_wallace._1255_ ),
    .A2(\u_cpu.ALU.u_wallace._1222_ ),
    .B1(\u_cpu.ALU.u_wallace._1446_ ),
    .C1(\u_cpu.ALU.u_wallace._1452_ ),
    .X(\u_cpu.ALU.u_wallace._1458_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._7172_  (.A1(\u_cpu.ALU.u_wallace._1446_ ),
    .A2(\u_cpu.ALU.u_wallace._1452_ ),
    .B1_N(\u_cpu.ALU.u_wallace._1455_ ),
    .Y(\u_cpu.ALU.u_wallace._1459_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._7173_  (.A1(\u_cpu.ALU.u_wallace._1458_ ),
    .A2(\u_cpu.ALU.u_wallace._1459_ ),
    .B1_N(\u_cpu.ALU.u_wallace._1254_ ),
    .Y(\u_cpu.ALU.u_wallace._1460_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._7174_  (.A1(\u_cpu.ALU.u_wallace._1009_ ),
    .A2(\u_cpu.ALU.u_wallace._1253_ ),
    .B1(\u_cpu.ALU.u_wallace._1457_ ),
    .C1(\u_cpu.ALU.u_wallace._1460_ ),
    .D1(\u_cpu.ALU.u_wallace._1240_ ),
    .Y(\u_cpu.ALU.u_wallace._1461_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7175_  (.A1(\u_cpu.ALU.u_wallace._1004_ ),
    .A2(\u_cpu.ALU.u_wallace._1019_ ),
    .B1(\u_cpu.ALU.u_wallace._1236_ ),
    .C1(\u_cpu.ALU.u_wallace._1239_ ),
    .X(\u_cpu.ALU.u_wallace._1462_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7176_  (.A(\u_cpu.ALU.u_wallace._1009_ ),
    .B(\u_cpu.ALU.u_wallace._1253_ ),
    .Y(\u_cpu.ALU.u_wallace._1463_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7177_  (.A(\u_cpu.ALU.u_wallace._1457_ ),
    .B(\u_cpu.ALU.u_wallace._1460_ ),
    .Y(\u_cpu.ALU.u_wallace._1464_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7178_  (.A1(\u_cpu.ALU.u_wallace._1462_ ),
    .A2(\u_cpu.ALU.u_wallace._1463_ ),
    .B1(\u_cpu.ALU.u_wallace._1464_ ),
    .Y(\u_cpu.ALU.u_wallace._1466_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._7179_  (.A(\u_cpu.ALU.u_wallace._1461_ ),
    .B(\u_cpu.ALU.u_wallace._1466_ ),
    .X(\u_cpu.ALU.u_wallace._1467_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7180_  (.A(\u_cpu.ALU.u_wallace._0795_ ),
    .B(\u_cpu.ALU.u_wallace._1015_ ),
    .C(\u_cpu.ALU.u_wallace._1250_ ),
    .X(\u_cpu.ALU.u_wallace._1468_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.ALU.u_wallace._7181_  (.A_N(\u_cpu.ALU.u_wallace._0427_ ),
    .B(\u_cpu.ALU.u_wallace._0591_ ),
    .C(\u_cpu.ALU.u_wallace._0593_ ),
    .D(\u_cpu.ALU.u_wallace._0429_ ),
    .X(\u_cpu.ALU.u_wallace._1469_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7182_  (.A1(\u_cpu.ALU.u_wallace._0795_ ),
    .A2(\u_cpu.ALU.u_wallace._1469_ ),
    .B1(\u_cpu.ALU.u_wallace._1017_ ),
    .Y(\u_cpu.ALU.u_wallace._1470_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7183_  (.A(\u_cpu.ALU.u_wallace._1015_ ),
    .B(\u_cpu.ALU.u_wallace._1250_ ),
    .Y(\u_cpu.ALU.u_wallace._1471_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7184_  (.A(\u_cpu.ALU.u_wallace._1247_ ),
    .B(\u_cpu.ALU.u_wallace._1240_ ),
    .C(\u_cpu.ALU.u_wallace._1242_ ),
    .D(\u_cpu.ALU.u_wallace._1009_ ),
    .X(\u_cpu.ALU.u_wallace._1472_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7185_  (.A1(\u_cpu.ALU.u_wallace._1250_ ),
    .A2(\u_cpu.ALU.u_wallace._1251_ ),
    .B1(\u_cpu.ALU.u_wallace._1472_ ),
    .Y(\u_cpu.ALU.u_wallace._1473_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7186_  (.A1(\u_cpu.ALU.u_wallace._1470_ ),
    .A2(\u_cpu.ALU.u_wallace._1471_ ),
    .B1(\u_cpu.ALU.u_wallace._1473_ ),
    .Y(\u_cpu.ALU.u_wallace._1474_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._7187_  (.A1(\u_cpu.ALU.u_wallace._1468_ ),
    .A2(\u_cpu.ALU.u_wallace._0601_ ),
    .A3(\u_cpu.ALU.u_wallace._0595_ ),
    .B1(\u_cpu.ALU.u_wallace._1474_ ),
    .Y(\u_cpu.ALU.u_wallace._1475_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._7188_  (.A(\u_cpu.ALU.u_wallace._1467_ ),
    .B(\u_cpu.ALU.u_wallace._1475_ ),
    .X(\u_cpu.ALU.Product_Wallace[20] ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7189_  (.A(\u_cpu.ALU.u_wallace._1457_ ),
    .Y(\u_cpu.ALU.u_wallace._1477_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7190_  (.A(\u_cpu.ALU.u_wallace._1460_ ),
    .B(\u_cpu.ALU.u_wallace._1462_ ),
    .Y(\u_cpu.ALU.u_wallace._1478_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._7191_  (.A1(\u_cpu.ALU.u_wallace._1429_ ),
    .A2(\u_cpu.ALU.u_wallace._1430_ ),
    .A3(\u_cpu.ALU.u_wallace._1431_ ),
    .B1(\u_cpu.ALU.u_wallace._1433_ ),
    .Y(\u_cpu.ALU.u_wallace._1479_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.ALU.u_wallace._7192_  (.A1(\u_cpu.ALU.u_wallace._1179_ ),
    .A2(\u_cpu.ALU.u_wallace._1177_ ),
    .A3(\u_cpu.ALU.u_wallace._1422_ ),
    .B1(\u_cpu.ALU.u_wallace._1428_ ),
    .B2(\u_cpu.ALU.u_wallace._1479_ ),
    .X(\u_cpu.ALU.u_wallace._1480_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7193_  (.A(\u_cpu.ALU.u_wallace._1434_ ),
    .B(\u_cpu.ALU.u_wallace._1394_ ),
    .C(\u_cpu.ALU.u_wallace._1427_ ),
    .X(\u_cpu.ALU.u_wallace._1481_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7194_  (.A1(\u_cpu.ALU.u_wallace._1384_ ),
    .A2(\u_cpu.ALU.u_wallace._1438_ ),
    .B1(\u_cpu.ALU.u_wallace._1440_ ),
    .Y(\u_cpu.ALU.u_wallace._1482_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7195_  (.A1(\u_cpu.ALU.u_wallace._1363_ ),
    .A2(\u_cpu.ALU.u_wallace._1360_ ),
    .B1(\u_cpu.ALU.u_wallace._1368_ ),
    .B2(\u_cpu.ALU.u_wallace._1359_ ),
    .X(\u_cpu.ALU.u_wallace._1483_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7196_  (.A1(\u_cpu.ALU.u_wallace._1330_ ),
    .A2(\u_cpu.ALU.u_wallace._1483_ ),
    .B1(\u_cpu.ALU.u_wallace._1372_ ),
    .Y(\u_cpu.ALU.u_wallace._1484_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7197_  (.A(\u_cpu.ALU.u_wallace._1351_ ),
    .Y(\u_cpu.ALU.u_wallace._1485_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7198_  (.A(\u_cpu.ALU.u_wallace._1307_ ),
    .B(\u_cpu.ALU.u_wallace._1310_ ),
    .Y(\u_cpu.ALU.u_wallace._1487_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._7199_  (.A1(\u_cpu.ALU.u_wallace._4678_ ),
    .A2(\u_cpu.ALU.u_wallace._0442_ ),
    .A3(\u_cpu.ALU.u_wallace._1085_ ),
    .B1(\u_cpu.ALU.u_wallace._1087_ ),
    .X(\u_cpu.ALU.u_wallace._1488_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7200_  (.A1(\u_cpu.ALU.u_wallace._1487_ ),
    .A2(\u_cpu.ALU.u_wallace._1488_ ),
    .B1(\u_cpu.ALU.u_wallace._1325_ ),
    .Y(\u_cpu.ALU.u_wallace._1489_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7201_  (.A1(\u_cpu.ALU.u_wallace._4550_ ),
    .A2(\u_cpu.ALU.SrcB[11] ),
    .B1(\u_cpu.ALU.SrcB[12] ),
    .B2(\u_cpu.ALU.u_wallace._4401_ ),
    .Y(\u_cpu.ALU.u_wallace._1490_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7202_  (.A(\u_cpu.ALU.u_wallace._4444_ ),
    .B(\u_cpu.ALU.u_wallace._4553_ ),
    .C(\u_cpu.ALU.u_wallace._4836_ ),
    .D(\u_cpu.ALU.u_wallace._4841_ ),
    .X(\u_cpu.ALU.u_wallace._1491_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7203_  (.A1(\u_cpu.ALU.u_wallace._1490_ ),
    .A2(\u_cpu.ALU.u_wallace._1491_ ),
    .B1(\u_cpu.ALU.u_wallace._4669_ ),
    .C1(\u_cpu.ALU.u_wallace._0034_ ),
    .Y(\u_cpu.ALU.u_wallace._1492_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._7204_  (.A1(\u_cpu.ALU.u_wallace._4669_ ),
    .A2(\u_cpu.ALU.u_wallace._0363_ ),
    .B1(\u_cpu.ALU.u_wallace._1490_ ),
    .C1(\u_cpu.ALU.u_wallace._1491_ ),
    .X(\u_cpu.ALU.u_wallace._1493_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7205_  (.A(\u_cpu.ALU.u_wallace._1492_ ),
    .B(\u_cpu.ALU.u_wallace._1493_ ),
    .Y(\u_cpu.ALU.u_wallace._1494_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7206_  (.A(\u_cpu.ALU.u_wallace._4007_ ),
    .B(\u_cpu.ALU.u_wallace._4291_ ),
    .C(\u_cpu.ALU.u_wallace._4900_ ),
    .D(\u_cpu.ALU.u_wallace._4909_ ),
    .Y(\u_cpu.ALU.u_wallace._1495_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7207_  (.A1(\u_cpu.ALU.u_wallace._4291_ ),
    .A2(\u_cpu.ALU.u_wallace._4790_ ),
    .B1(\u_cpu.ALU.u_wallace._4909_ ),
    .B2(\u_cpu.ALU.u_wallace._4007_ ),
    .X(\u_cpu.ALU.u_wallace._1496_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._7208_  (.A1_N(\u_cpu.ALU.u_wallace._4601_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0169_ ),
    .B1(\u_cpu.ALU.u_wallace._1495_ ),
    .B2(\u_cpu.ALU.u_wallace._1496_ ),
    .Y(\u_cpu.ALU.u_wallace._1498_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7209_  (.A1(\u_cpu.ALU.u_wallace._4598_ ),
    .A2(\u_cpu.ALU.u_wallace._4900_ ),
    .B1(\u_cpu.ALU.u_wallace._4907_ ),
    .B2(\u_cpu.ALU.u_wallace._4716_ ),
    .Y(\u_cpu.ALU.u_wallace._1499_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7210_  (.A(\u_cpu.ALU.u_wallace._1495_ ),
    .B(\u_cpu.ALU.u_wallace._4794_ ),
    .C(\u_cpu.ALU.u_wallace._4604_ ),
    .Y(\u_cpu.ALU.u_wallace._1500_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7211_  (.A(\u_cpu.ALU.u_wallace._1499_ ),
    .B(\u_cpu.ALU.u_wallace._1500_ ),
    .Y(\u_cpu.ALU.u_wallace._1501_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7212_  (.A(\u_cpu.ALU.u_wallace._4551_ ),
    .B(\u_cpu.ALU.u_wallace._0041_ ),
    .Y(\u_cpu.ALU.u_wallace._1502_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7213_  (.A1(\u_cpu.ALU.u_wallace._1502_ ),
    .A2(\u_cpu.ALU.u_wallace._1334_ ),
    .B1(\u_cpu.ALU.u_wallace._1331_ ),
    .Y(\u_cpu.ALU.u_wallace._1503_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._7214_  (.A1(\u_cpu.ALU.u_wallace._1498_ ),
    .A2(\u_cpu.ALU.u_wallace._1501_ ),
    .B1_N(\u_cpu.ALU.u_wallace._1503_ ),
    .Y(\u_cpu.ALU.u_wallace._1504_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7215_  (.A1(\u_cpu.ALU.u_wallace._4604_ ),
    .A2(\u_cpu.ALU.u_wallace._4798_ ),
    .B1(\u_cpu.ALU.u_wallace._1495_ ),
    .B2(\u_cpu.ALU.u_wallace._1496_ ),
    .X(\u_cpu.ALU.u_wallace._1505_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7216_  (.A1(\u_cpu.ALU.u_wallace._1499_ ),
    .A2(\u_cpu.ALU.u_wallace._1500_ ),
    .B1(\u_cpu.ALU.u_wallace._1503_ ),
    .C1(\u_cpu.ALU.u_wallace._1505_ ),
    .Y(\u_cpu.ALU.u_wallace._1506_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7217_  (.A(\u_cpu.ALU.u_wallace._1494_ ),
    .B(\u_cpu.ALU.u_wallace._1504_ ),
    .C(\u_cpu.ALU.u_wallace._1506_ ),
    .Y(\u_cpu.ALU.u_wallace._1507_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._7218_  (.A1(\u_cpu.ALU.u_wallace._4677_ ),
    .A2(\u_cpu.ALU.u_wallace._0037_ ),
    .B1(\u_cpu.ALU.u_wallace._1490_ ),
    .B2(\u_cpu.ALU.u_wallace._1491_ ),
    .X(\u_cpu.ALU.u_wallace._1509_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7219_  (.A(\u_cpu.ALU.u_wallace._4444_ ),
    .B(\u_cpu.ALU.u_wallace._4550_ ),
    .C(\u_cpu.ALU.u_wallace._4836_ ),
    .D(\u_cpu.ALU.SrcB[12] ),
    .Y(\u_cpu.ALU.u_wallace._1510_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.ALU.u_wallace._7220_  (.A_N(\u_cpu.ALU.u_wallace._1490_ ),
    .B(\u_cpu.ALU.u_wallace._1510_ ),
    .C(\u_cpu.ALU.u_wallace._4669_ ),
    .D(\u_cpu.ALU.u_wallace._0057_ ),
    .X(\u_cpu.ALU.u_wallace._1511_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7221_  (.A1_N(\u_cpu.ALU.u_wallace._1506_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1504_ ),
    .B1(\u_cpu.ALU.u_wallace._1509_ ),
    .B2(\u_cpu.ALU.u_wallace._1511_ ),
    .Y(\u_cpu.ALU.u_wallace._1512_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7222_  (.A1(\u_cpu.ALU.u_wallace._1316_ ),
    .A2(\u_cpu.ALU.u_wallace._1489_ ),
    .B1(\u_cpu.ALU.u_wallace._1507_ ),
    .C1(\u_cpu.ALU.u_wallace._1512_ ),
    .X(\u_cpu.ALU.u_wallace._1513_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7223_  (.A1(\u_cpu.ALU.u_wallace._1325_ ),
    .A2(\u_cpu.ALU.u_wallace._1317_ ),
    .B1(\u_cpu.ALU.u_wallace._1312_ ),
    .Y(\u_cpu.ALU.u_wallace._1514_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7224_  (.A1(\u_cpu.ALU.u_wallace._1507_ ),
    .A2(\u_cpu.ALU.u_wallace._1512_ ),
    .B1(\u_cpu.ALU.u_wallace._1514_ ),
    .Y(\u_cpu.ALU.u_wallace._1515_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._7225_  (.A1(\u_cpu.ALU.u_wallace._1339_ ),
    .A2(\u_cpu.ALU.u_wallace._1485_ ),
    .B1(\u_cpu.ALU.u_wallace._1513_ ),
    .B2(\u_cpu.ALU.u_wallace._1515_ ),
    .X(\u_cpu.ALU.u_wallace._1516_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7226_  (.A1(\u_cpu.ALU.u_wallace._1507_ ),
    .A2(\u_cpu.ALU.u_wallace._1512_ ),
    .B1(\u_cpu.ALU.u_wallace._1514_ ),
    .X(\u_cpu.ALU.u_wallace._1517_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._7227_  (.A1(\u_cpu.ALU.u_wallace._1342_ ),
    .A2(\u_cpu.ALU.u_wallace._1340_ ),
    .A3(\u_cpu.ALU.u_wallace._1341_ ),
    .B1(\u_cpu.ALU.u_wallace._1351_ ),
    .X(\u_cpu.ALU.u_wallace._1518_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7228_  (.A1(\u_cpu.ALU.u_wallace._1316_ ),
    .A2(\u_cpu.ALU.u_wallace._1489_ ),
    .B1(\u_cpu.ALU.u_wallace._1507_ ),
    .C1(\u_cpu.ALU.u_wallace._1512_ ),
    .Y(\u_cpu.ALU.u_wallace._1520_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7229_  (.A(\u_cpu.ALU.u_wallace._1517_ ),
    .B(\u_cpu.ALU.u_wallace._1518_ ),
    .C(\u_cpu.ALU.u_wallace._1520_ ),
    .X(\u_cpu.ALU.u_wallace._1521_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7230_  (.A(\u_cpu.ALU.SrcA[21] ),
    .Y(\u_cpu.ALU.u_wallace._1522_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7231_  (.A1(\u_cpu.ALU.u_wallace._4649_ ),
    .A2(\u_cpu.ALU.u_wallace._0324_ ),
    .B1(\u_cpu.ALU.u_wallace._0813_ ),
    .B2(\u_cpu.ALU.u_wallace._0895_ ),
    .Y(\u_cpu.ALU.u_wallace._1523_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7232_  (.A(\u_cpu.ALU.u_wallace._1815_ ),
    .B(\u_cpu.ALU.SrcA[4] ),
    .C(\u_cpu.ALU.SrcA[15] ),
    .D(\u_cpu.ALU.u_wallace._0628_ ),
    .X(\u_cpu.ALU.u_wallace._1524_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7233_  (.A1(\u_cpu.ALU.u_wallace._0634_ ),
    .A2(\u_cpu.ALU.u_wallace._1522_ ),
    .B1(\u_cpu.ALU.u_wallace._1523_ ),
    .B2(\u_cpu.ALU.u_wallace._1524_ ),
    .Y(\u_cpu.ALU.u_wallace._1525_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7234_  (.A(\u_cpu.ALU.u_wallace._1815_ ),
    .B(\u_cpu.ALU.SrcA[15] ),
    .Y(\u_cpu.ALU.u_wallace._1526_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7235_  (.A(\u_cpu.ALU.SrcA[4] ),
    .B(\u_cpu.ALU.SrcB[17] ),
    .Y(\u_cpu.ALU.u_wallace._1527_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7236_  (.A(\u_cpu.ALU.u_wallace._1526_ ),
    .B(\u_cpu.ALU.u_wallace._1527_ ),
    .Y(\u_cpu.ALU.u_wallace._1528_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7237_  (.A(\u_cpu.ALU.u_wallace._4649_ ),
    .B(\u_cpu.ALU.SrcA[4] ),
    .C(\u_cpu.ALU.u_wallace._0324_ ),
    .D(\u_cpu.ALU.u_wallace._0813_ ),
    .Y(\u_cpu.ALU.u_wallace._1529_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7238_  (.A(\u_cpu.ALU.SrcA[21] ),
    .X(\u_cpu.ALU.u_wallace._1531_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7239_  (.A(\u_cpu.ALU.u_wallace._1528_ ),
    .B(\u_cpu.ALU.u_wallace._1529_ ),
    .C(\u_cpu.ALU.u_wallace._0873_ ),
    .D(\u_cpu.ALU.u_wallace._1531_ ),
    .Y(\u_cpu.ALU.u_wallace._1532_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7240_  (.A1(\u_cpu.ALU.u_wallace._1265_ ),
    .A2(\u_cpu.ALU.u_wallace._1264_ ),
    .B1(\u_cpu.ALU.u_wallace._1277_ ),
    .Y(\u_cpu.ALU.u_wallace._1533_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7241_  (.A1(\u_cpu.ALU.u_wallace._1525_ ),
    .A2(\u_cpu.ALU.u_wallace._1532_ ),
    .B1(\u_cpu.ALU.u_wallace._1533_ ),
    .Y(\u_cpu.ALU.u_wallace._1534_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7242_  (.A(\u_cpu.ALU.SrcA[21] ),
    .X(\u_cpu.ALU.u_wallace._1535_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7243_  (.A1(\u_cpu.ALU.u_wallace._1859_ ),
    .A2(\u_cpu.ALU.u_wallace._1535_ ),
    .B1(\u_cpu.ALU.u_wallace._1528_ ),
    .B2(\u_cpu.ALU.u_wallace._1529_ ),
    .Y(\u_cpu.ALU.u_wallace._1536_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7244_  (.A(\u_cpu.ALU.u_wallace._1771_ ),
    .B(\u_cpu.ALU.u_wallace._0177_ ),
    .Y(\u_cpu.ALU.u_wallace._1537_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7245_  (.A(\u_cpu.ALU.u_wallace._0600_ ),
    .B(\u_cpu.ALU.u_wallace._0639_ ),
    .Y(\u_cpu.ALU.u_wallace._1538_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7246_  (.A1(\u_cpu.ALU.u_wallace._1537_ ),
    .A2(\u_cpu.ALU.u_wallace._1538_ ),
    .B1(\u_cpu.ALU.u_wallace._1265_ ),
    .Y(\u_cpu.ALU.u_wallace._1539_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7247_  (.A1(\u_cpu.ALU.u_wallace._1272_ ),
    .A2(\u_cpu.ALU.u_wallace._1539_ ),
    .B1(\u_cpu.ALU.u_wallace._1532_ ),
    .Y(\u_cpu.ALU.u_wallace._1540_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7248_  (.A1(\u_cpu.ALU.u_wallace._0534_ ),
    .A2(\u_cpu.ALU.SrcA[19] ),
    .B1(\u_cpu.ALU.u_wallace._1270_ ),
    .B2(\u_cpu.ALU.u_wallace._0775_ ),
    .X(\u_cpu.ALU.u_wallace._1542_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7249_  (.A(\u_cpu.ALU.SrcA[20] ),
    .X(\u_cpu.ALU.u_wallace._1543_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7250_  (.A(\u_cpu.ALU.u_wallace._0742_ ),
    .B(\u_cpu.ALU.u_wallace._0808_ ),
    .Y(\u_cpu.ALU.u_wallace._1544_ ));
 sky130_fd_sc_hd__a41oi_2 \u_cpu.ALU.u_wallace._7251_  (.A1(\u_cpu.ALU.u_wallace._0187_ ),
    .A2(\u_cpu.ALU.u_wallace._0304_ ),
    .A3(\u_cpu.ALU.u_wallace._1090_ ),
    .A4(\u_cpu.ALU.u_wallace._1543_ ),
    .B1(\u_cpu.ALU.u_wallace._1544_ ),
    .Y(\u_cpu.ALU.u_wallace._1545_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7252_  (.A(\u_cpu.ALU.u_wallace._0775_ ),
    .B(\u_cpu.ALU.u_wallace._0534_ ),
    .C(\u_cpu.ALU.SrcA[19] ),
    .D(\u_cpu.ALU.SrcA[20] ),
    .Y(\u_cpu.ALU.u_wallace._1546_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7253_  (.A1(\u_cpu.ALU.u_wallace._0753_ ),
    .A2(\u_cpu.ALU.u_wallace._0815_ ),
    .B1(\u_cpu.ALU.u_wallace._1542_ ),
    .B2(\u_cpu.ALU.u_wallace._1546_ ),
    .Y(\u_cpu.ALU.u_wallace._1547_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7254_  (.A1(\u_cpu.ALU.u_wallace._1542_ ),
    .A2(\u_cpu.ALU.u_wallace._1545_ ),
    .B1(\u_cpu.ALU.u_wallace._1547_ ),
    .Y(\u_cpu.ALU.u_wallace._1548_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7255_  (.A1(\u_cpu.ALU.u_wallace._1536_ ),
    .A2(\u_cpu.ALU.u_wallace._1540_ ),
    .B1(\u_cpu.ALU.u_wallace._1548_ ),
    .Y(\u_cpu.ALU.u_wallace._1549_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7256_  (.A1(\u_cpu.ALU.u_wallace._1264_ ),
    .A2(\u_cpu.ALU.u_wallace._1266_ ),
    .B1(\u_cpu.ALU.u_wallace._1273_ ),
    .Y(\u_cpu.ALU.u_wallace._1550_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7257_  (.A1(\u_cpu.ALU.u_wallace._1261_ ),
    .A2(\u_cpu.ALU.u_wallace._1260_ ),
    .B1(\u_cpu.ALU.u_wallace._1263_ ),
    .Y(\u_cpu.ALU.u_wallace._1551_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7258_  (.A1(\u_cpu.ALU.u_wallace._1550_ ),
    .A2(\u_cpu.ALU.u_wallace._1281_ ),
    .B1(\u_cpu.ALU.u_wallace._1551_ ),
    .Y(\u_cpu.ALU.u_wallace._1553_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7259_  (.A(\u_cpu.ALU.u_wallace._1542_ ),
    .B(\u_cpu.ALU.u_wallace._1546_ ),
    .C(\u_cpu.ALU.u_wallace._4662_ ),
    .D(\u_cpu.ALU.u_wallace._0815_ ),
    .X(\u_cpu.ALU.u_wallace._1554_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7260_  (.A(\u_cpu.ALU.u_wallace._1529_ ),
    .B(\u_cpu.ALU.u_wallace._1535_ ),
    .C(\u_cpu.ALU.u_wallace._1859_ ),
    .Y(\u_cpu.ALU.u_wallace._1555_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._7261_  (.A1(\u_cpu.ALU.u_wallace._1523_ ),
    .A2(\u_cpu.ALU.u_wallace._1555_ ),
    .B1(\u_cpu.ALU.u_wallace._1539_ ),
    .B2(\u_cpu.ALU.u_wallace._1272_ ),
    .C1(\u_cpu.ALU.u_wallace._1525_ ),
    .X(\u_cpu.ALU.u_wallace._1556_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7262_  (.A1(\u_cpu.ALU.u_wallace._1547_ ),
    .A2(\u_cpu.ALU.u_wallace._1554_ ),
    .B1(\u_cpu.ALU.u_wallace._1556_ ),
    .B2(\u_cpu.ALU.u_wallace._1534_ ),
    .Y(\u_cpu.ALU.u_wallace._1557_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._7263_  (.A1(\u_cpu.ALU.u_wallace._1534_ ),
    .A2(\u_cpu.ALU.u_wallace._1549_ ),
    .B1(\u_cpu.ALU.u_wallace._1288_ ),
    .B2(\u_cpu.ALU.u_wallace._1553_ ),
    .C1(\u_cpu.ALU.u_wallace._1557_ ),
    .X(\u_cpu.ALU.u_wallace._1558_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7264_  (.A1(\u_cpu.ALU.u_wallace._1556_ ),
    .A2(\u_cpu.ALU.u_wallace._1534_ ),
    .B1(\u_cpu.ALU.u_wallace._1548_ ),
    .Y(\u_cpu.ALU.u_wallace._1559_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7265_  (.A1(\u_cpu.ALU.u_wallace._1526_ ),
    .A2(\u_cpu.ALU.u_wallace._1527_ ),
    .B1(\u_cpu.ALU.u_wallace._1555_ ),
    .Y(\u_cpu.ALU.u_wallace._1560_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._7266_  (.A1(\u_cpu.ALU.u_wallace._1536_ ),
    .A2(\u_cpu.ALU.u_wallace._1560_ ),
    .B1_N(\u_cpu.ALU.u_wallace._1533_ ),
    .Y(\u_cpu.ALU.u_wallace._1561_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._7267_  (.A1(\u_cpu.ALU.u_wallace._1547_ ),
    .A2(\u_cpu.ALU.u_wallace._1554_ ),
    .B1(\u_cpu.ALU.u_wallace._1536_ ),
    .B2(\u_cpu.ALU.u_wallace._1540_ ),
    .C1(\u_cpu.ALU.u_wallace._1561_ ),
    .Y(\u_cpu.ALU.u_wallace._1562_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._7268_  (.A1(\u_cpu.ALU.u_wallace._1265_ ),
    .A2(\u_cpu.ALU.u_wallace._1264_ ),
    .A3(\u_cpu.ALU.u_wallace._1272_ ),
    .B1(\u_cpu.ALU.u_wallace._1269_ ),
    .X(\u_cpu.ALU.u_wallace._1564_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7269_  (.A1(\u_cpu.ALU.u_wallace._1273_ ),
    .A2(\u_cpu.ALU.u_wallace._1564_ ),
    .B1(\u_cpu.ALU.u_wallace._1282_ ),
    .B2(\u_cpu.ALU.u_wallace._1294_ ),
    .Y(\u_cpu.ALU.u_wallace._1565_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7270_  (.A(\u_cpu.ALU.u_wallace._1559_ ),
    .B(\u_cpu.ALU.u_wallace._1562_ ),
    .C(\u_cpu.ALU.u_wallace._1565_ ),
    .Y(\u_cpu.ALU.u_wallace._1566_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7271_  (.A1(\u_cpu.ALU.u_wallace._1486_ ),
    .A2(\u_cpu.ALU.u_wallace._0447_ ),
    .B1(\u_cpu.ALU.SrcA[17] ),
    .B2(\u_cpu.ALU.u_wallace._1026_ ),
    .X(\u_cpu.ALU.u_wallace._1567_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7272_  (.A(\u_cpu.ALU.u_wallace._4467_ ),
    .B(\u_cpu.ALU.u_wallace._1497_ ),
    .C(\u_cpu.ALU.u_wallace._0448_ ),
    .D(\u_cpu.ALU.u_wallace._1073_ ),
    .Y(\u_cpu.ALU.u_wallace._1568_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7273_  (.A1(\u_cpu.ALU.u_wallace._3404_ ),
    .A2(\u_cpu.ALU.u_wallace._0179_ ),
    .B1(\u_cpu.ALU.u_wallace._1567_ ),
    .B2(\u_cpu.ALU.u_wallace._1568_ ),
    .Y(\u_cpu.ALU.u_wallace._1569_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7274_  (.A1(\u_cpu.ALU.u_wallace._1259_ ),
    .A2(\u_cpu.ALU.u_wallace._1261_ ),
    .B1(\u_cpu.ALU.u_wallace._1285_ ),
    .Y(\u_cpu.ALU.u_wallace._1570_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7275_  (.A(\u_cpu.ALU.u_wallace._2144_ ),
    .B(\u_cpu.ALU.u_wallace._1541_ ),
    .C(\u_cpu.ALU.u_wallace._0441_ ),
    .Y(\u_cpu.ALU.u_wallace._1571_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._7276_  (.A1(\u_cpu.ALU.u_wallace._0635_ ),
    .A2(\u_cpu.ALU.u_wallace._1571_ ),
    .B1(\u_cpu.ALU.u_wallace._2604_ ),
    .C1(\u_cpu.ALU.u_wallace._0652_ ),
    .D1(\u_cpu.ALU.u_wallace._1567_ ),
    .Y(\u_cpu.ALU.u_wallace._1572_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7277_  (.A(\u_cpu.ALU.u_wallace._1570_ ),
    .B(\u_cpu.ALU.u_wallace._1572_ ),
    .Y(\u_cpu.ALU.u_wallace._1573_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._7278_  (.A(\u_cpu.ALU.SrcB[7] ),
    .B(\u_cpu.ALU.SrcA[14] ),
    .X(\u_cpu.ALU.u_wallace._1575_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7279_  (.A1(\u_cpu.ALU.u_wallace._0635_ ),
    .A2(\u_cpu.ALU.u_wallace._1571_ ),
    .B1(\u_cpu.ALU.u_wallace._1575_ ),
    .C1(\u_cpu.ALU.u_wallace._1567_ ),
    .X(\u_cpu.ALU.u_wallace._1576_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._7280_  (.A1(\u_cpu.ALU.u_wallace._1569_ ),
    .A2(\u_cpu.ALU.u_wallace._1576_ ),
    .B1_N(\u_cpu.ALU.u_wallace._1570_ ),
    .Y(\u_cpu.ALU.u_wallace._1577_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7281_  (.A(\u_cpu.ALU.u_wallace._0188_ ),
    .X(\u_cpu.ALU.u_wallace._1578_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7282_  (.A1(\u_cpu.ALU.u_wallace._1305_ ),
    .A2(\u_cpu.ALU.u_wallace._1578_ ),
    .A3(\u_cpu.ALU.u_wallace._2604_ ),
    .B1(\u_cpu.ALU.u_wallace._1309_ ),
    .X(\u_cpu.ALU.u_wallace._1579_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7283_  (.A1(\u_cpu.ALU.u_wallace._1569_ ),
    .A2(\u_cpu.ALU.u_wallace._1573_ ),
    .B1(\u_cpu.ALU.u_wallace._1577_ ),
    .C1(\u_cpu.ALU.u_wallace._1579_ ),
    .Y(\u_cpu.ALU.u_wallace._1580_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7284_  (.A1(\u_cpu.ALU.u_wallace._2626_ ),
    .A2(\u_cpu.ALU.u_wallace._0320_ ),
    .B1(\u_cpu.ALU.u_wallace._1567_ ),
    .B2(\u_cpu.ALU.u_wallace._1568_ ),
    .X(\u_cpu.ALU.u_wallace._1581_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7285_  (.A(\u_cpu.ALU.u_wallace._1570_ ),
    .B(\u_cpu.ALU.u_wallace._1581_ ),
    .C(\u_cpu.ALU.u_wallace._1572_ ),
    .Y(\u_cpu.ALU.u_wallace._1582_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7286_  (.A1(\u_cpu.ALU.u_wallace._1582_ ),
    .A2(\u_cpu.ALU.u_wallace._1577_ ),
    .B1(\u_cpu.ALU.u_wallace._1579_ ),
    .X(\u_cpu.ALU.u_wallace._1583_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7287_  (.A(\u_cpu.ALU.u_wallace._1566_ ),
    .B(\u_cpu.ALU.u_wallace._1580_ ),
    .C(\u_cpu.ALU.u_wallace._1583_ ),
    .Y(\u_cpu.ALU.u_wallace._1584_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._7288_  (.A1(\u_cpu.ALU.u_wallace._1534_ ),
    .A2(\u_cpu.ALU.u_wallace._1549_ ),
    .B1(\u_cpu.ALU.u_wallace._1288_ ),
    .B2(\u_cpu.ALU.u_wallace._1553_ ),
    .C1(\u_cpu.ALU.u_wallace._1557_ ),
    .Y(\u_cpu.ALU.u_wallace._1586_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7289_  (.A(\u_cpu.ALU.u_wallace._1579_ ),
    .B(\u_cpu.ALU.u_wallace._1582_ ),
    .C(\u_cpu.ALU.u_wallace._1577_ ),
    .X(\u_cpu.ALU.u_wallace._1587_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7290_  (.A1(\u_cpu.ALU.u_wallace._1582_ ),
    .A2(\u_cpu.ALU.u_wallace._1577_ ),
    .B1(\u_cpu.ALU.u_wallace._1579_ ),
    .Y(\u_cpu.ALU.u_wallace._1588_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7291_  (.A1_N(\u_cpu.ALU.u_wallace._1586_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1566_ ),
    .B1(\u_cpu.ALU.u_wallace._1587_ ),
    .B2(\u_cpu.ALU.u_wallace._1588_ ),
    .Y(\u_cpu.ALU.u_wallace._1589_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7292_  (.A(\u_cpu.ALU.u_wallace._1283_ ),
    .Y(\u_cpu.ALU.u_wallace._1590_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7293_  (.A(\u_cpu.ALU.u_wallace._1258_ ),
    .B(\u_cpu.ALU.u_wallace._1292_ ),
    .Y(\u_cpu.ALU.u_wallace._1591_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7294_  (.A1_N(\u_cpu.ALU.u_wallace._1299_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1327_ ),
    .B1(\u_cpu.ALU.u_wallace._1590_ ),
    .B2(\u_cpu.ALU.u_wallace._1591_ ),
    .Y(\u_cpu.ALU.u_wallace._1592_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7295_  (.A1(\u_cpu.ALU.u_wallace._1558_ ),
    .A2(\u_cpu.ALU.u_wallace._1584_ ),
    .B1(\u_cpu.ALU.u_wallace._1589_ ),
    .C1(\u_cpu.ALU.u_wallace._1592_ ),
    .Y(\u_cpu.ALU.u_wallace._1593_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7296_  (.A(\u_cpu.ALU.u_wallace._1586_ ),
    .B(\u_cpu.ALU.u_wallace._1566_ ),
    .C(\u_cpu.ALU.u_wallace._1580_ ),
    .D(\u_cpu.ALU.u_wallace._1583_ ),
    .Y(\u_cpu.ALU.u_wallace._1594_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7297_  (.A1(\u_cpu.ALU.u_wallace._1589_ ),
    .A2(\u_cpu.ALU.u_wallace._1594_ ),
    .B1(\u_cpu.ALU.u_wallace._1592_ ),
    .X(\u_cpu.ALU.u_wallace._1595_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7298_  (.A1(\u_cpu.ALU.u_wallace._1516_ ),
    .A2(\u_cpu.ALU.u_wallace._1521_ ),
    .B1(\u_cpu.ALU.u_wallace._1593_ ),
    .C1(\u_cpu.ALU.u_wallace._1595_ ),
    .Y(\u_cpu.ALU.u_wallace._1597_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7299_  (.A1(\u_cpu.ALU.u_wallace._1339_ ),
    .A2(\u_cpu.ALU.u_wallace._1485_ ),
    .B1(\u_cpu.ALU.u_wallace._1520_ ),
    .C1(\u_cpu.ALU.u_wallace._1517_ ),
    .Y(\u_cpu.ALU.u_wallace._1598_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7300_  (.A1(\u_cpu.ALU.u_wallace._1513_ ),
    .A2(\u_cpu.ALU.u_wallace._1515_ ),
    .B1(\u_cpu.ALU.u_wallace._1518_ ),
    .Y(\u_cpu.ALU.u_wallace._1599_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7301_  (.A1(\u_cpu.ALU.u_wallace._1558_ ),
    .A2(\u_cpu.ALU.u_wallace._1584_ ),
    .B1(\u_cpu.ALU.u_wallace._1589_ ),
    .C1(\u_cpu.ALU.u_wallace._1592_ ),
    .X(\u_cpu.ALU.u_wallace._1600_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7302_  (.A1(\u_cpu.ALU.u_wallace._1589_ ),
    .A2(\u_cpu.ALU.u_wallace._1594_ ),
    .B1(\u_cpu.ALU.u_wallace._1592_ ),
    .Y(\u_cpu.ALU.u_wallace._1601_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7303_  (.A1_N(\u_cpu.ALU.u_wallace._1598_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1599_ ),
    .B1(\u_cpu.ALU.u_wallace._1600_ ),
    .B2(\u_cpu.ALU.u_wallace._1601_ ),
    .Y(\u_cpu.ALU.u_wallace._1602_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7304_  (.A(\u_cpu.ALU.u_wallace._1484_ ),
    .B(\u_cpu.ALU.u_wallace._1597_ ),
    .C(\u_cpu.ALU.u_wallace._1602_ ),
    .X(\u_cpu.ALU.u_wallace._1603_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7305_  (.A1(\u_cpu.ALU.u_wallace._1516_ ),
    .A2(\u_cpu.ALU.u_wallace._1521_ ),
    .B1(\u_cpu.ALU.u_wallace._1600_ ),
    .B2(\u_cpu.ALU.u_wallace._1601_ ),
    .Y(\u_cpu.ALU.u_wallace._1604_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7306_  (.A1(\u_cpu.ALU.u_wallace._1352_ ),
    .A2(\u_cpu.ALU.u_wallace._1351_ ),
    .B1(\u_cpu.ALU.u_wallace._1520_ ),
    .B2(\u_cpu.ALU.u_wallace._1517_ ),
    .X(\u_cpu.ALU.u_wallace._1605_ ));
 sky130_fd_sc_hd__or3b_2 \u_cpu.ALU.u_wallace._7307_  (.A(\u_cpu.ALU.u_wallace._1513_ ),
    .B(\u_cpu.ALU.u_wallace._1515_ ),
    .C_N(\u_cpu.ALU.u_wallace._1518_ ),
    .X(\u_cpu.ALU.u_wallace._1606_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7308_  (.A(\u_cpu.ALU.u_wallace._1605_ ),
    .B(\u_cpu.ALU.u_wallace._1606_ ),
    .C(\u_cpu.ALU.u_wallace._1593_ ),
    .D(\u_cpu.ALU.u_wallace._1595_ ),
    .Y(\u_cpu.ALU.u_wallace._1608_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._7309_  (.A1(\u_cpu.ALU.u_wallace._1483_ ),
    .A2(\u_cpu.ALU.u_wallace._1330_ ),
    .B1(\u_cpu.ALU.u_wallace._1372_ ),
    .C1(\u_cpu.ALU.u_wallace._1604_ ),
    .D1(\u_cpu.ALU.u_wallace._1608_ ),
    .Y(\u_cpu.ALU.u_wallace._1609_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7310_  (.A(\u_cpu.ALU.SrcB[21] ),
    .X(\u_cpu.ALU.u_wallace._1610_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7311_  (.A(\u_cpu.ALU.u_wallace._1610_ ),
    .X(\u_cpu.ALU.u_wallace._1611_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7312_  (.A1(\u_cpu.ALU.u_wallace._0764_ ),
    .A2(\u_cpu.ALU.u_wallace._0957_ ),
    .B1(\u_cpu.ALU.SrcB[19] ),
    .B2(\u_cpu.ALU.u_wallace._0392_ ),
    .X(\u_cpu.ALU.u_wallace._1612_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7313_  (.A(\u_cpu.ALU.u_wallace._4597_ ),
    .B(\u_cpu.ALU.u_wallace._1421_ ),
    .C(\u_cpu.ALU.u_wallace._0958_ ),
    .D(\u_cpu.ALU.u_wallace._1208_ ),
    .Y(\u_cpu.ALU.u_wallace._1613_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7314_  (.A1(\u_cpu.ALU.u_wallace._0162_ ),
    .A2(\u_cpu.ALU.u_wallace._1392_ ),
    .B1(\u_cpu.ALU.u_wallace._1612_ ),
    .B2(\u_cpu.ALU.u_wallace._1613_ ),
    .X(\u_cpu.ALU.u_wallace._1614_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7315_  (.A(\u_cpu.ALU.u_wallace._1386_ ),
    .X(\u_cpu.ALU.u_wallace._1615_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7316_  (.A(\u_cpu.ALU.u_wallace._1612_ ),
    .B(\u_cpu.ALU.u_wallace._1613_ ),
    .C(\u_cpu.ALU.u_wallace._0272_ ),
    .D(\u_cpu.ALU.u_wallace._1615_ ),
    .Y(\u_cpu.ALU.u_wallace._1616_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7317_  (.A(\u_cpu.ALU.u_wallace._1410_ ),
    .B(\u_cpu.ALU.u_wallace._0731_ ),
    .C(\u_cpu.ALU.u_wallace._1387_ ),
    .D(\u_cpu.ALU.u_wallace._1175_ ),
    .X(\u_cpu.ALU.u_wallace._1617_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7318_  (.A1(\u_cpu.ALU.u_wallace._1390_ ),
    .A2(\u_cpu.ALU.u_wallace._1392_ ),
    .A3(\u_cpu.ALU.u_wallace._0108_ ),
    .B1(\u_cpu.ALU.u_wallace._1617_ ),
    .X(\u_cpu.ALU.u_wallace._1619_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7319_  (.A1(\u_cpu.ALU.u_wallace._1614_ ),
    .A2(\u_cpu.ALU.u_wallace._1616_ ),
    .B1(\u_cpu.ALU.u_wallace._1619_ ),
    .X(\u_cpu.ALU.u_wallace._1620_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7320_  (.A(\u_cpu.ALU.u_wallace._1619_ ),
    .B(\u_cpu.ALU.u_wallace._1614_ ),
    .C(\u_cpu.ALU.u_wallace._1616_ ),
    .Y(\u_cpu.ALU.u_wallace._1621_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7321_  (.A1(\u_cpu.ALU.u_wallace._3996_ ),
    .A2(\u_cpu.ALU.u_wallace._1611_ ),
    .B1(\u_cpu.ALU.u_wallace._1620_ ),
    .B2(\u_cpu.ALU.u_wallace._1621_ ),
    .X(\u_cpu.ALU.u_wallace._1622_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7322_  (.A(\u_cpu.ALU.u_wallace._1620_ ),
    .B(\u_cpu.ALU.u_wallace._1621_ ),
    .C(\u_cpu.ALU.u_wallace._0129_ ),
    .D(\u_cpu.ALU.u_wallace._1611_ ),
    .Y(\u_cpu.ALU.u_wallace._1623_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7323_  (.A1(\u_cpu.ALU.u_wallace._2790_ ),
    .A2(\u_cpu.ALU.u_wallace._0727_ ),
    .B1(\u_cpu.ALU.u_wallace._0728_ ),
    .B2(\u_cpu.ALU.u_wallace._2834_ ),
    .Y(\u_cpu.ALU.u_wallace._1624_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7324_  (.A(\u_cpu.ALU.u_wallace._2878_ ),
    .B(\u_cpu.ALU.u_wallace._1782_ ),
    .C(\u_cpu.ALU.SrcB[14] ),
    .D(\u_cpu.ALU.u_wallace._0278_ ),
    .X(\u_cpu.ALU.u_wallace._1625_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7325_  (.A1(\u_cpu.ALU.u_wallace._4812_ ),
    .A2(\u_cpu.ALU.u_wallace._0553_ ),
    .B1(\u_cpu.ALU.u_wallace._1624_ ),
    .B2(\u_cpu.ALU.u_wallace._1625_ ),
    .Y(\u_cpu.ALU.u_wallace._1626_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7326_  (.A1(\u_cpu.ALU.u_wallace._2878_ ),
    .A2(\u_cpu.ALU.u_wallace._0727_ ),
    .B1(\u_cpu.ALU.u_wallace._0278_ ),
    .B2(\u_cpu.ALU.u_wallace._1837_ ),
    .X(\u_cpu.ALU.u_wallace._1627_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7327_  (.A(\u_cpu.ALU.u_wallace._4447_ ),
    .B(\u_cpu.ALU.u_wallace._2834_ ),
    .C(\u_cpu.ALU.u_wallace._0120_ ),
    .D(\u_cpu.ALU.u_wallace._0728_ ),
    .Y(\u_cpu.ALU.u_wallace._1628_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7328_  (.A(\u_cpu.ALU.u_wallace._1627_ ),
    .B(\u_cpu.ALU.u_wallace._1628_ ),
    .C(\u_cpu.ALU.u_wallace._4529_ ),
    .D(\u_cpu.ALU.u_wallace._0550_ ),
    .Y(\u_cpu.ALU.u_wallace._1630_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7329_  (.A1(\u_cpu.ALU.u_wallace._4412_ ),
    .A2(\u_cpu.ALU.u_wallace._0364_ ),
    .B1(\u_cpu.ALU.u_wallace._0144_ ),
    .B2(\u_cpu.ALU.u_wallace._4561_ ),
    .Y(\u_cpu.ALU.u_wallace._1631_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7330_  (.A1(\u_cpu.ALU.u_wallace._1347_ ),
    .A2(\u_cpu.ALU.u_wallace._1631_ ),
    .B1(\u_cpu.ALU.u_wallace._1346_ ),
    .Y(\u_cpu.ALU.u_wallace._1632_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7331_  (.A1(\u_cpu.ALU.u_wallace._1626_ ),
    .A2(\u_cpu.ALU.u_wallace._1630_ ),
    .B1(\u_cpu.ALU.u_wallace._1632_ ),
    .Y(\u_cpu.ALU.u_wallace._1633_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7332_  (.A(\u_cpu.ALU.u_wallace._1626_ ),
    .B(\u_cpu.ALU.u_wallace._1630_ ),
    .C(\u_cpu.ALU.u_wallace._1632_ ),
    .X(\u_cpu.ALU.u_wallace._1634_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._7333_  (.A1(\u_cpu.ALU.u_wallace._0939_ ),
    .A2(\u_cpu.ALU.u_wallace._0941_ ),
    .A3(\u_cpu.ALU.u_wallace._1400_ ),
    .B1(\u_cpu.ALU.u_wallace._1401_ ),
    .X(\u_cpu.ALU.u_wallace._1635_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7334_  (.A1(\u_cpu.ALU.u_wallace._1633_ ),
    .A2(\u_cpu.ALU.u_wallace._1634_ ),
    .B1(\u_cpu.ALU.u_wallace._1635_ ),
    .Y(\u_cpu.ALU.u_wallace._1636_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7335_  (.A1(\u_cpu.ALU.u_wallace._1626_ ),
    .A2(\u_cpu.ALU.u_wallace._1630_ ),
    .B1(\u_cpu.ALU.u_wallace._1632_ ),
    .X(\u_cpu.ALU.u_wallace._1637_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7336_  (.A(\u_cpu.ALU.u_wallace._1626_ ),
    .B(\u_cpu.ALU.u_wallace._1630_ ),
    .C(\u_cpu.ALU.u_wallace._1632_ ),
    .Y(\u_cpu.ALU.u_wallace._1638_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._7337_  (.A_N(\u_cpu.ALU.u_wallace._1635_ ),
    .B(\u_cpu.ALU.u_wallace._1637_ ),
    .C(\u_cpu.ALU.u_wallace._1638_ ),
    .Y(\u_cpu.ALU.u_wallace._1639_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7338_  (.A1(\u_cpu.ALU.u_wallace._1413_ ),
    .A2(\u_cpu.ALU.u_wallace._1412_ ),
    .B1(\u_cpu.ALU.u_wallace._1416_ ),
    .Y(\u_cpu.ALU.u_wallace._1641_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7339_  (.A1(\u_cpu.ALU.u_wallace._1636_ ),
    .A2(\u_cpu.ALU.u_wallace._1639_ ),
    .B1(\u_cpu.ALU.u_wallace._1641_ ),
    .Y(\u_cpu.ALU.u_wallace._1642_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7340_  (.A(\u_cpu.ALU.u_wallace._1641_ ),
    .B(\u_cpu.ALU.u_wallace._1636_ ),
    .C(\u_cpu.ALU.u_wallace._1639_ ),
    .X(\u_cpu.ALU.u_wallace._1643_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7341_  (.A1_N(\u_cpu.ALU.u_wallace._1622_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1623_ ),
    .B1(\u_cpu.ALU.u_wallace._1642_ ),
    .B2(\u_cpu.ALU.u_wallace._1643_ ),
    .Y(\u_cpu.ALU.u_wallace._1644_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7342_  (.A1(\u_cpu.ALU.u_wallace._1636_ ),
    .A2(\u_cpu.ALU.u_wallace._1639_ ),
    .B1(\u_cpu.ALU.u_wallace._1641_ ),
    .X(\u_cpu.ALU.u_wallace._1645_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7343_  (.A(\u_cpu.ALU.u_wallace._1641_ ),
    .B(\u_cpu.ALU.u_wallace._1636_ ),
    .C(\u_cpu.ALU.u_wallace._1639_ ),
    .Y(\u_cpu.ALU.u_wallace._1646_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7344_  (.A(\u_cpu.ALU.u_wallace._1622_ ),
    .B(\u_cpu.ALU.u_wallace._1623_ ),
    .C(\u_cpu.ALU.u_wallace._1645_ ),
    .D(\u_cpu.ALU.u_wallace._1646_ ),
    .Y(\u_cpu.ALU.u_wallace._1647_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.ALU.u_wallace._7345_  (.A1_N(\u_cpu.ALU.u_wallace._1365_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1361_ ),
    .B1(\u_cpu.ALU.u_wallace._1374_ ),
    .B2(\u_cpu.ALU.u_wallace._1367_ ),
    .X(\u_cpu.ALU.u_wallace._1648_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7346_  (.A1(\u_cpu.ALU.u_wallace._1644_ ),
    .A2(\u_cpu.ALU.u_wallace._1647_ ),
    .B1(\u_cpu.ALU.u_wallace._1648_ ),
    .X(\u_cpu.ALU.u_wallace._1649_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7347_  (.A(\u_cpu.ALU.u_wallace._1648_ ),
    .B(\u_cpu.ALU.u_wallace._1644_ ),
    .C(\u_cpu.ALU.u_wallace._1647_ ),
    .Y(\u_cpu.ALU.u_wallace._1650_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7348_  (.A(\u_cpu.ALU.u_wallace._1435_ ),
    .B(\u_cpu.ALU.u_wallace._1649_ ),
    .C(\u_cpu.ALU.u_wallace._1650_ ),
    .Y(\u_cpu.ALU.u_wallace._1652_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7349_  (.A1(\u_cpu.ALU.u_wallace._1644_ ),
    .A2(\u_cpu.ALU.u_wallace._1647_ ),
    .B1(\u_cpu.ALU.u_wallace._1648_ ),
    .Y(\u_cpu.ALU.u_wallace._1653_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7350_  (.A(\u_cpu.ALU.u_wallace._1648_ ),
    .B(\u_cpu.ALU.u_wallace._1644_ ),
    .C(\u_cpu.ALU.u_wallace._1647_ ),
    .X(\u_cpu.ALU.u_wallace._1654_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._7351_  (.A1(\u_cpu.ALU.u_wallace._1394_ ),
    .A2(\u_cpu.ALU.u_wallace._1423_ ),
    .A3(\u_cpu.ALU.u_wallace._1425_ ),
    .B1(\u_cpu.ALU.u_wallace._1415_ ),
    .X(\u_cpu.ALU.u_wallace._1655_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7352_  (.A1(\u_cpu.ALU.u_wallace._1653_ ),
    .A2(\u_cpu.ALU.u_wallace._1654_ ),
    .B1(\u_cpu.ALU.u_wallace._1655_ ),
    .Y(\u_cpu.ALU.u_wallace._1656_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7353_  (.A(\u_cpu.ALU.u_wallace._1609_ ),
    .B(\u_cpu.ALU.u_wallace._1652_ ),
    .C(\u_cpu.ALU.u_wallace._1656_ ),
    .Y(\u_cpu.ALU.u_wallace._1657_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7354_  (.A(\u_cpu.ALU.u_wallace._1484_ ),
    .B(\u_cpu.ALU.u_wallace._1597_ ),
    .C(\u_cpu.ALU.u_wallace._1602_ ),
    .Y(\u_cpu.ALU.u_wallace._1658_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7355_  (.A(\u_cpu.ALU.u_wallace._1658_ ),
    .B(\u_cpu.ALU.u_wallace._1609_ ),
    .Y(\u_cpu.ALU.u_wallace._1659_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7356_  (.A(\u_cpu.ALU.u_wallace._1652_ ),
    .B(\u_cpu.ALU.u_wallace._1656_ ),
    .Y(\u_cpu.ALU.u_wallace._1660_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._7357_  (.A1_N(\u_cpu.ALU.u_wallace._1603_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1657_ ),
    .B1(\u_cpu.ALU.u_wallace._1659_ ),
    .B2(\u_cpu.ALU.u_wallace._1660_ ),
    .Y(\u_cpu.ALU.u_wallace._1661_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7358_  (.A1(\u_cpu.ALU.u_wallace._1480_ ),
    .A2(\u_cpu.ALU.u_wallace._1481_ ),
    .B1(\u_cpu.ALU.u_wallace._1482_ ),
    .B2(\u_cpu.ALU.u_wallace._1661_ ),
    .Y(\u_cpu.ALU.u_wallace._1663_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7359_  (.A(\u_cpu.ALU.u_wallace._1435_ ),
    .B(\u_cpu.ALU.u_wallace._1649_ ),
    .C(\u_cpu.ALU.u_wallace._1650_ ),
    .X(\u_cpu.ALU.u_wallace._1664_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._7360_  (.A1(\u_cpu.ALU.u_wallace._1396_ ),
    .A2(\u_cpu.ALU.u_wallace._1425_ ),
    .B1(\u_cpu.ALU.u_wallace._1653_ ),
    .B2(\u_cpu.ALU.u_wallace._1654_ ),
    .C1(\u_cpu.ALU.u_wallace._1415_ ),
    .X(\u_cpu.ALU.u_wallace._1665_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7361_  (.A1_N(\u_cpu.ALU.u_wallace._1658_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1609_ ),
    .B1(\u_cpu.ALU.u_wallace._1664_ ),
    .B2(\u_cpu.ALU.u_wallace._1665_ ),
    .Y(\u_cpu.ALU.u_wallace._1666_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7362_  (.A1(\u_cpu.ALU.u_wallace._1603_ ),
    .A2(\u_cpu.ALU.u_wallace._1657_ ),
    .B1(\u_cpu.ALU.u_wallace._1666_ ),
    .C1(\u_cpu.ALU.u_wallace._1482_ ),
    .X(\u_cpu.ALU.u_wallace._1667_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU.u_wallace._7363_  (.A(\u_cpu.ALU.u_wallace._1480_ ),
    .B(\u_cpu.ALU.u_wallace._1481_ ),
    .X(\u_cpu.ALU.u_wallace._1668_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7364_  (.A(\u_cpu.ALU.u_wallace._1658_ ),
    .B(\u_cpu.ALU.u_wallace._1609_ ),
    .C(\u_cpu.ALU.u_wallace._1652_ ),
    .D(\u_cpu.ALU.u_wallace._1656_ ),
    .Y(\u_cpu.ALU.u_wallace._1669_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7365_  (.A1(\u_cpu.ALU.u_wallace._1669_ ),
    .A2(\u_cpu.ALU.u_wallace._1666_ ),
    .B1(\u_cpu.ALU.u_wallace._1482_ ),
    .Y(\u_cpu.ALU.u_wallace._1670_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7366_  (.A(\u_cpu.ALU.u_wallace._1667_ ),
    .B(\u_cpu.ALU.u_wallace._1670_ ),
    .Y(\u_cpu.ALU.u_wallace._1671_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7367_  (.A(\u_cpu.ALU.u_wallace._1446_ ),
    .B(\u_cpu.ALU.u_wallace._1453_ ),
    .Y(\u_cpu.ALU.u_wallace._1672_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._7368_  (.A1(\u_cpu.ALU.u_wallace._1663_ ),
    .A2(\u_cpu.ALU.u_wallace._1667_ ),
    .B1(\u_cpu.ALU.u_wallace._1668_ ),
    .B2(\u_cpu.ALU.u_wallace._1671_ ),
    .C1(\u_cpu.ALU.u_wallace._1672_ ),
    .Y(\u_cpu.ALU.u_wallace._1674_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7369_  (.A1(\u_cpu.ALU.u_wallace._1482_ ),
    .A2(\u_cpu.ALU.u_wallace._1669_ ),
    .A3(\u_cpu.ALU.u_wallace._1666_ ),
    .B1(\u_cpu.ALU.u_wallace._1663_ ),
    .X(\u_cpu.ALU.u_wallace._1675_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7370_  (.A(\u_cpu.ALU.u_wallace._1480_ ),
    .B(\u_cpu.ALU.u_wallace._1481_ ),
    .Y(\u_cpu.ALU.u_wallace._1676_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7371_  (.A1(\u_cpu.ALU.u_wallace._1667_ ),
    .A2(\u_cpu.ALU.u_wallace._1670_ ),
    .B1(\u_cpu.ALU.u_wallace._1676_ ),
    .Y(\u_cpu.ALU.u_wallace._1677_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7372_  (.A1(\u_cpu.ALU.u_wallace._1675_ ),
    .A2(\u_cpu.ALU.u_wallace._1677_ ),
    .B1(\u_cpu.ALU.u_wallace._1672_ ),
    .X(\u_cpu.ALU.u_wallace._1678_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7373_  (.A(\u_cpu.ALU.u_wallace._1478_ ),
    .B(\u_cpu.ALU.u_wallace._1674_ ),
    .C(\u_cpu.ALU.u_wallace._1678_ ),
    .Y(\u_cpu.ALU.u_wallace._1679_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._7374_  (.A1(\u_cpu.ALU.u_wallace._1663_ ),
    .A2(\u_cpu.ALU.u_wallace._1667_ ),
    .B1(\u_cpu.ALU.u_wallace._1668_ ),
    .B2(\u_cpu.ALU.u_wallace._1671_ ),
    .C1(\u_cpu.ALU.u_wallace._1672_ ),
    .X(\u_cpu.ALU.u_wallace._1680_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7375_  (.A1(\u_cpu.ALU.u_wallace._1675_ ),
    .A2(\u_cpu.ALU.u_wallace._1677_ ),
    .B1(\u_cpu.ALU.u_wallace._1672_ ),
    .Y(\u_cpu.ALU.u_wallace._1681_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7376_  (.A1_N(\u_cpu.ALU.u_wallace._1457_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1478_ ),
    .B1(\u_cpu.ALU.u_wallace._1680_ ),
    .B2(\u_cpu.ALU.u_wallace._1681_ ),
    .Y(\u_cpu.ALU.u_wallace._1682_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7377_  (.A1(\u_cpu.ALU.u_wallace._1477_ ),
    .A2(\u_cpu.ALU.u_wallace._1679_ ),
    .B1(\u_cpu.ALU.u_wallace._1682_ ),
    .Y(\u_cpu.ALU.u_wallace._1683_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7378_  (.A(\u_cpu.ALU.u_wallace._1463_ ),
    .B(\u_cpu.ALU.u_wallace._1457_ ),
    .C(\u_cpu.ALU.u_wallace._1460_ ),
    .D(\u_cpu.ALU.u_wallace._1240_ ),
    .X(\u_cpu.ALU.u_wallace._1685_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._7379_  (.A1(\u_cpu.ALU.u_wallace._1467_ ),
    .A2(\u_cpu.ALU.u_wallace._1475_ ),
    .B1_N(\u_cpu.ALU.u_wallace._1685_ ),
    .Y(\u_cpu.ALU.u_wallace._1686_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._7380_  (.A(\u_cpu.ALU.u_wallace._1683_ ),
    .B(\u_cpu.ALU.u_wallace._1686_ ),
    .X(\u_cpu.ALU.Product_Wallace[21] ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7381_  (.A1(\u_cpu.ALU.u_wallace._1667_ ),
    .A2(\u_cpu.ALU.u_wallace._1663_ ),
    .B1(\u_cpu.ALU.u_wallace._1677_ ),
    .Y(\u_cpu.ALU.u_wallace._1687_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._7382_  (.A1(\u_cpu.ALU.u_wallace._1451_ ),
    .A2(\u_cpu.ALU.u_wallace._1449_ ),
    .A3(\u_cpu.ALU.u_wallace._1450_ ),
    .B1(\u_cpu.ALU.u_wallace._1453_ ),
    .X(\u_cpu.ALU.u_wallace._1688_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7383_  (.A1(\u_cpu.ALU.u_wallace._1687_ ),
    .A2(\u_cpu.ALU.u_wallace._1688_ ),
    .B1(\u_cpu.ALU.u_wallace._1457_ ),
    .Y(\u_cpu.ALU.u_wallace._1689_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.ALU.u_wallace._7384_  (.A1_N(\u_cpu.ALU.u_wallace._1573_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1569_ ),
    .B1(\u_cpu.ALU.u_wallace._1579_ ),
    .B2(\u_cpu.ALU.u_wallace._1577_ ),
    .X(\u_cpu.ALU.u_wallace._1690_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7385_  (.A1(\u_cpu.ALU.u_wallace._4797_ ),
    .A2(\u_cpu.ALU.u_wallace._4836_ ),
    .B1(\u_cpu.ALU.u_wallace._4841_ ),
    .B2(\u_cpu.ALU.u_wallace._4557_ ),
    .X(\u_cpu.ALU.u_wallace._1691_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7386_  (.A(\u_cpu.ALU.u_wallace._4551_ ),
    .B(\u_cpu.ALU.u_wallace._4653_ ),
    .C(\u_cpu.ALU.u_wallace._4731_ ),
    .D(\u_cpu.ALU.u_wallace._0144_ ),
    .Y(\u_cpu.ALU.u_wallace._1692_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7387_  (.A(\u_cpu.ALU.u_wallace._4567_ ),
    .B(\u_cpu.ALU.u_wallace._0033_ ),
    .Y(\u_cpu.ALU.u_wallace._1693_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7388_  (.A1(\u_cpu.ALU.u_wallace._1691_ ),
    .A2(\u_cpu.ALU.u_wallace._1692_ ),
    .B1(\u_cpu.ALU.u_wallace._1693_ ),
    .Y(\u_cpu.ALU.u_wallace._1695_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7389_  (.A(\u_cpu.ALU.u_wallace._1693_ ),
    .B(\u_cpu.ALU.u_wallace._1691_ ),
    .C(\u_cpu.ALU.u_wallace._1692_ ),
    .X(\u_cpu.ALU.u_wallace._1696_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7390_  (.A1(\u_cpu.ALU.u_wallace._4291_ ),
    .A2(\u_cpu.ALU.u_wallace._4920_ ),
    .B1(\u_cpu.ALU.u_wallace._0182_ ),
    .B2(\u_cpu.ALU.u_wallace._4007_ ),
    .Y(\u_cpu.ALU.u_wallace._1697_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7391_  (.A(\u_cpu.ALU.u_wallace._0041_ ),
    .B(\u_cpu.ALU.u_wallace._4900_ ),
    .Y(\u_cpu.ALU.u_wallace._1698_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._7392_  (.A1(\u_cpu.ALU.u_wallace._4594_ ),
    .A2(\u_cpu.ALU.u_wallace._4595_ ),
    .A3(\u_cpu.ALU.u_wallace._4921_ ),
    .A4(\u_cpu.ALU.u_wallace._0179_ ),
    .B1(\u_cpu.ALU.u_wallace._1698_ ),
    .X(\u_cpu.ALU.u_wallace._1699_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7393_  (.A(\u_cpu.ALU.u_wallace._0041_ ),
    .B(\u_cpu.ALU.u_wallace._4653_ ),
    .Y(\u_cpu.ALU.u_wallace._1700_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7394_  (.A1(\u_cpu.ALU.u_wallace._1700_ ),
    .A2(\u_cpu.ALU.u_wallace._1499_ ),
    .B1(\u_cpu.ALU.u_wallace._1495_ ),
    .Y(\u_cpu.ALU.u_wallace._1701_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7395_  (.A(\u_cpu.ALU.u_wallace._4716_ ),
    .B(\u_cpu.ALU.u_wallace._4598_ ),
    .C(\u_cpu.ALU.u_wallace._4909_ ),
    .D(\u_cpu.ALU.u_wallace._0177_ ),
    .Y(\u_cpu.ALU.u_wallace._1702_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7396_  (.A1(\u_cpu.ALU.u_wallace._4598_ ),
    .A2(\u_cpu.ALU.u_wallace._4909_ ),
    .B1(\u_cpu.ALU.u_wallace._0177_ ),
    .B2(\u_cpu.ALU.u_wallace._4716_ ),
    .X(\u_cpu.ALU.u_wallace._1703_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7397_  (.A1_N(\u_cpu.ALU.u_wallace._1702_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1703_ ),
    .B1(\u_cpu.ALU.u_wallace._4601_ ),
    .B2(\u_cpu.ALU.u_wallace._4913_ ),
    .Y(\u_cpu.ALU.u_wallace._1704_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7398_  (.A1(\u_cpu.ALU.u_wallace._1697_ ),
    .A2(\u_cpu.ALU.u_wallace._1699_ ),
    .B1(\u_cpu.ALU.u_wallace._1701_ ),
    .C1(\u_cpu.ALU.u_wallace._1704_ ),
    .Y(\u_cpu.ALU.u_wallace._1706_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7399_  (.A(\u_cpu.ALU.u_wallace._1703_ ),
    .B(\u_cpu.ALU.u_wallace._0475_ ),
    .C(\u_cpu.ALU.u_wallace._0052_ ),
    .D(\u_cpu.ALU.u_wallace._1702_ ),
    .Y(\u_cpu.ALU.u_wallace._1707_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7400_  (.A1(\u_cpu.ALU.u_wallace._1704_ ),
    .A2(\u_cpu.ALU.u_wallace._1707_ ),
    .B1(\u_cpu.ALU.u_wallace._1701_ ),
    .X(\u_cpu.ALU.u_wallace._1708_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7401_  (.A1(\u_cpu.ALU.u_wallace._1695_ ),
    .A2(\u_cpu.ALU.u_wallace._1696_ ),
    .B1(\u_cpu.ALU.u_wallace._1706_ ),
    .C1(\u_cpu.ALU.u_wallace._1708_ ),
    .Y(\u_cpu.ALU.u_wallace._1709_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7402_  (.A1(\u_cpu.ALU.u_wallace._1697_ ),
    .A2(\u_cpu.ALU.u_wallace._1699_ ),
    .B1(\u_cpu.ALU.u_wallace._1701_ ),
    .C1(\u_cpu.ALU.u_wallace._1704_ ),
    .X(\u_cpu.ALU.u_wallace._1710_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7403_  (.A1(\u_cpu.ALU.u_wallace._1704_ ),
    .A2(\u_cpu.ALU.u_wallace._1707_ ),
    .B1(\u_cpu.ALU.u_wallace._1701_ ),
    .Y(\u_cpu.ALU.u_wallace._1711_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7404_  (.A(\u_cpu.ALU.u_wallace._1695_ ),
    .B(\u_cpu.ALU.u_wallace._1696_ ),
    .Y(\u_cpu.ALU.u_wallace._1712_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7405_  (.A1(\u_cpu.ALU.u_wallace._1710_ ),
    .A2(\u_cpu.ALU.u_wallace._1711_ ),
    .B1(\u_cpu.ALU.u_wallace._1712_ ),
    .Y(\u_cpu.ALU.u_wallace._1713_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7406_  (.A(\u_cpu.ALU.u_wallace._1690_ ),
    .B(\u_cpu.ALU.u_wallace._1709_ ),
    .C(\u_cpu.ALU.u_wallace._1713_ ),
    .Y(\u_cpu.ALU.u_wallace._1714_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._7407_  (.A1(\u_cpu.ALU.u_wallace._1579_ ),
    .A2(\u_cpu.ALU.u_wallace._1577_ ),
    .B1_N(\u_cpu.ALU.u_wallace._1582_ ),
    .Y(\u_cpu.ALU.u_wallace._1715_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7408_  (.A1(\u_cpu.ALU.u_wallace._1695_ ),
    .A2(\u_cpu.ALU.u_wallace._1696_ ),
    .B1(\u_cpu.ALU.u_wallace._1710_ ),
    .B2(\u_cpu.ALU.u_wallace._1711_ ),
    .Y(\u_cpu.ALU.u_wallace._1717_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7409_  (.A(\u_cpu.ALU.u_wallace._1708_ ),
    .B(\u_cpu.ALU.u_wallace._1712_ ),
    .C(\u_cpu.ALU.u_wallace._1706_ ),
    .Y(\u_cpu.ALU.u_wallace._1718_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7410_  (.A(\u_cpu.ALU.u_wallace._1715_ ),
    .B(\u_cpu.ALU.u_wallace._1717_ ),
    .C(\u_cpu.ALU.u_wallace._1718_ ),
    .Y(\u_cpu.ALU.u_wallace._1719_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._7411_  (.A1(\u_cpu.ALU.u_wallace._1494_ ),
    .A2(\u_cpu.ALU.u_wallace._1504_ ),
    .B1_N(\u_cpu.ALU.u_wallace._1506_ ),
    .Y(\u_cpu.ALU.u_wallace._1720_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7412_  (.A1(\u_cpu.ALU.u_wallace._1714_ ),
    .A2(\u_cpu.ALU.u_wallace._1719_ ),
    .B1(\u_cpu.ALU.u_wallace._1720_ ),
    .Y(\u_cpu.ALU.u_wallace._1721_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7413_  (.A(\u_cpu.ALU.u_wallace._1714_ ),
    .B(\u_cpu.ALU.u_wallace._1719_ ),
    .C(\u_cpu.ALU.u_wallace._1720_ ),
    .X(\u_cpu.ALU.u_wallace._1722_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7414_  (.A1_N(\u_cpu.ALU.u_wallace._1548_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1561_ ),
    .B1(\u_cpu.ALU.u_wallace._1540_ ),
    .B2(\u_cpu.ALU.u_wallace._1536_ ),
    .Y(\u_cpu.ALU.u_wallace._1723_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7415_  (.A(\u_cpu.ALU.u_wallace._0742_ ),
    .B(\u_cpu.ALU.u_wallace._1100_ ),
    .Y(\u_cpu.ALU.u_wallace._1724_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._7416_  (.A1(\u_cpu.ALU.u_wallace._1158_ ),
    .A2(\u_cpu.ALU.u_wallace._0545_ ),
    .A3(\u_cpu.ALU.u_wallace._1543_ ),
    .A4(\u_cpu.ALU.u_wallace._1535_ ),
    .B1(\u_cpu.ALU.u_wallace._1724_ ),
    .X(\u_cpu.ALU.u_wallace._1725_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7417_  (.A1(\u_cpu.ALU.u_wallace._0293_ ),
    .A2(\u_cpu.ALU.SrcA[20] ),
    .B1(\u_cpu.ALU.SrcA[21] ),
    .B2(\u_cpu.ALU.u_wallace._0797_ ),
    .Y(\u_cpu.ALU.u_wallace._1726_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7418_  (.A(\u_cpu.ALU.u_wallace._0775_ ),
    .B(\u_cpu.ALU.u_wallace._0534_ ),
    .C(\u_cpu.ALU.SrcA[20] ),
    .D(\u_cpu.ALU.SrcA[21] ),
    .X(\u_cpu.ALU.u_wallace._1728_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7419_  (.A1(\u_cpu.ALU.u_wallace._1726_ ),
    .A2(\u_cpu.ALU.u_wallace._1728_ ),
    .B1(\u_cpu.ALU.u_wallace._1724_ ),
    .Y(\u_cpu.ALU.u_wallace._1729_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7420_  (.A(\u_cpu.ALU.SrcA[21] ),
    .X(\u_cpu.ALU.u_wallace._1730_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7421_  (.A(\u_cpu.ALU.u_wallace._0075_ ),
    .B(\u_cpu.ALU.u_wallace._1730_ ),
    .Y(\u_cpu.ALU.u_wallace._1731_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7422_  (.A1(\u_cpu.ALU.u_wallace._1526_ ),
    .A2(\u_cpu.ALU.u_wallace._1527_ ),
    .B1(\u_cpu.ALU.u_wallace._1731_ ),
    .Y(\u_cpu.ALU.u_wallace._1732_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7423_  (.A(\u_cpu.ALU.u_wallace._1815_ ),
    .B(\u_cpu.ALU.u_wallace._1114_ ),
    .C(\u_cpu.ALU.u_wallace._0447_ ),
    .D(\u_cpu.ALU.u_wallace._0628_ ),
    .Y(\u_cpu.ALU.u_wallace._1733_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7424_  (.A(\u_cpu.ALU.SrcA[22] ),
    .X(\u_cpu.ALU.u_wallace._1734_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7425_  (.A(\u_cpu.ALU.u_wallace._1733_ ),
    .B(\u_cpu.ALU.u_wallace._1734_ ),
    .C(\u_cpu.ALU.u_wallace._1749_ ),
    .Y(\u_cpu.ALU.u_wallace._1735_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7426_  (.A1(\u_cpu.ALU.u_wallace._1760_ ),
    .A2(\u_cpu.ALU.u_wallace._0447_ ),
    .B1(\u_cpu.ALU.u_wallace._0628_ ),
    .B2(\u_cpu.ALU.u_wallace._1114_ ),
    .Y(\u_cpu.ALU.u_wallace._1736_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7427_  (.A(\u_cpu.ALU.SrcA[22] ),
    .Y(\u_cpu.ALU.u_wallace._1737_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7428_  (.A(\u_cpu.ALU.u_wallace._1815_ ),
    .B(\u_cpu.ALU.u_wallace._1114_ ),
    .C(\u_cpu.ALU.u_wallace._0447_ ),
    .D(\u_cpu.ALU.u_wallace._0628_ ),
    .X(\u_cpu.ALU.u_wallace._1739_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7429_  (.A1(\u_cpu.ALU.u_wallace._0634_ ),
    .A2(\u_cpu.ALU.u_wallace._1737_ ),
    .B1(\u_cpu.ALU.u_wallace._1736_ ),
    .B2(\u_cpu.ALU.u_wallace._1739_ ),
    .Y(\u_cpu.ALU.u_wallace._1740_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._7430_  (.A1(\u_cpu.ALU.u_wallace._1524_ ),
    .A2(\u_cpu.ALU.u_wallace._1732_ ),
    .B1(\u_cpu.ALU.u_wallace._1735_ ),
    .B2(\u_cpu.ALU.u_wallace._1736_ ),
    .C1(\u_cpu.ALU.u_wallace._1740_ ),
    .Y(\u_cpu.ALU.u_wallace._1741_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7431_  (.A(\u_cpu.ALU.SrcA[22] ),
    .X(\u_cpu.ALU.u_wallace._1742_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7432_  (.A1(\u_cpu.ALU.u_wallace._3678_ ),
    .A2(\u_cpu.ALU.u_wallace._0441_ ),
    .B1(\u_cpu.ALU.u_wallace._0639_ ),
    .B2(\u_cpu.ALU.u_wallace._1311_ ),
    .X(\u_cpu.ALU.u_wallace._1743_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7433_  (.A1(\u_cpu.ALU.u_wallace._2757_ ),
    .A2(\u_cpu.ALU.u_wallace._1742_ ),
    .B1(\u_cpu.ALU.u_wallace._1743_ ),
    .B2(\u_cpu.ALU.u_wallace._1733_ ),
    .Y(\u_cpu.ALU.u_wallace._1744_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7434_  (.A(\u_cpu.ALU.u_wallace._1736_ ),
    .B(\u_cpu.ALU.u_wallace._1735_ ),
    .Y(\u_cpu.ALU.u_wallace._1745_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._7435_  (.A1(\u_cpu.ALU.u_wallace._0634_ ),
    .A2(\u_cpu.ALU.u_wallace._1522_ ),
    .A3(\u_cpu.ALU.u_wallace._1523_ ),
    .B1(\u_cpu.ALU.u_wallace._1529_ ),
    .X(\u_cpu.ALU.u_wallace._1746_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7436_  (.A1(\u_cpu.ALU.u_wallace._1744_ ),
    .A2(\u_cpu.ALU.u_wallace._1745_ ),
    .B1(\u_cpu.ALU.u_wallace._1746_ ),
    .Y(\u_cpu.ALU.u_wallace._1747_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._7437_  (.A1(\u_cpu.ALU.u_wallace._1725_ ),
    .A2(\u_cpu.ALU.u_wallace._1726_ ),
    .B1(\u_cpu.ALU.u_wallace._1729_ ),
    .C1(\u_cpu.ALU.u_wallace._1741_ ),
    .D1(\u_cpu.ALU.u_wallace._1747_ ),
    .Y(\u_cpu.ALU.u_wallace._1748_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._7438_  (.A1(\u_cpu.ALU.u_wallace._4678_ ),
    .A2(\u_cpu.ALU.u_wallace._1096_ ),
    .B1(\u_cpu.ALU.u_wallace._1726_ ),
    .B2(\u_cpu.ALU.u_wallace._1728_ ),
    .X(\u_cpu.ALU.u_wallace._1750_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7439_  (.A1(\u_cpu.ALU.u_wallace._0545_ ),
    .A2(\u_cpu.ALU.u_wallace._1270_ ),
    .B1(\u_cpu.ALU.u_wallace._1535_ ),
    .B2(\u_cpu.ALU.u_wallace._1957_ ),
    .X(\u_cpu.ALU.u_wallace._1751_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7440_  (.A(\u_cpu.ALU.u_wallace._0187_ ),
    .B(\u_cpu.ALU.u_wallace._0304_ ),
    .C(\u_cpu.ALU.u_wallace._1543_ ),
    .D(\u_cpu.ALU.u_wallace._1535_ ),
    .Y(\u_cpu.ALU.u_wallace._1752_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7441_  (.A(\u_cpu.ALU.u_wallace._1751_ ),
    .B(\u_cpu.ALU.u_wallace._1752_ ),
    .C(\u_cpu.ALU.u_wallace._0578_ ),
    .D(\u_cpu.ALU.u_wallace._1101_ ),
    .X(\u_cpu.ALU.u_wallace._1753_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._7442_  (.A1(\u_cpu.ALU.u_wallace._1736_ ),
    .A2(\u_cpu.ALU.u_wallace._1735_ ),
    .B1(\u_cpu.ALU.u_wallace._1732_ ),
    .B2(\u_cpu.ALU.u_wallace._1524_ ),
    .C1(\u_cpu.ALU.u_wallace._1740_ ),
    .X(\u_cpu.ALU.u_wallace._1754_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7443_  (.A(\u_cpu.ALU.u_wallace._1743_ ),
    .B(\u_cpu.ALU.u_wallace._1733_ ),
    .C(\u_cpu.ALU.u_wallace._2757_ ),
    .D(\u_cpu.ALU.u_wallace._1742_ ),
    .Y(\u_cpu.ALU.u_wallace._1755_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7444_  (.A1(\u_cpu.ALU.u_wallace._1731_ ),
    .A2(\u_cpu.ALU.u_wallace._1523_ ),
    .B1(\u_cpu.ALU.u_wallace._1529_ ),
    .Y(\u_cpu.ALU.u_wallace._1756_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7445_  (.A1(\u_cpu.ALU.u_wallace._1740_ ),
    .A2(\u_cpu.ALU.u_wallace._1755_ ),
    .B1(\u_cpu.ALU.u_wallace._1756_ ),
    .Y(\u_cpu.ALU.u_wallace._1757_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7446_  (.A1(\u_cpu.ALU.u_wallace._1750_ ),
    .A2(\u_cpu.ALU.u_wallace._1753_ ),
    .B1(\u_cpu.ALU.u_wallace._1754_ ),
    .B2(\u_cpu.ALU.u_wallace._1757_ ),
    .Y(\u_cpu.ALU.u_wallace._1758_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7447_  (.A(\u_cpu.ALU.u_wallace._1723_ ),
    .B(\u_cpu.ALU.u_wallace._1748_ ),
    .C(\u_cpu.ALU.u_wallace._1758_ ),
    .Y(\u_cpu.ALU.u_wallace._1759_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._7448_  (.A1(\u_cpu.ALU.u_wallace._1726_ ),
    .A2(\u_cpu.ALU.u_wallace._1725_ ),
    .B1(\u_cpu.ALU.u_wallace._1729_ ),
    .X(\u_cpu.ALU.u_wallace._1761_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7449_  (.A1(\u_cpu.ALU.u_wallace._1754_ ),
    .A2(\u_cpu.ALU.u_wallace._1757_ ),
    .B1(\u_cpu.ALU.u_wallace._1761_ ),
    .Y(\u_cpu.ALU.u_wallace._1762_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7450_  (.A1(\u_cpu.ALU.u_wallace._1750_ ),
    .A2(\u_cpu.ALU.u_wallace._1753_ ),
    .B1(\u_cpu.ALU.u_wallace._1741_ ),
    .C1(\u_cpu.ALU.u_wallace._1747_ ),
    .Y(\u_cpu.ALU.u_wallace._1763_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.ALU.u_wallace._7451_  (.A1(\u_cpu.ALU.u_wallace._1731_ ),
    .A2(\u_cpu.ALU.u_wallace._1523_ ),
    .A3(\u_cpu.ALU.u_wallace._1524_ ),
    .B1(\u_cpu.ALU.u_wallace._1539_ ),
    .B2(\u_cpu.ALU.u_wallace._1272_ ),
    .X(\u_cpu.ALU.u_wallace._1764_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7452_  (.A1(\u_cpu.ALU.u_wallace._1525_ ),
    .A2(\u_cpu.ALU.u_wallace._1764_ ),
    .B1(\u_cpu.ALU.u_wallace._1561_ ),
    .B2(\u_cpu.ALU.u_wallace._1548_ ),
    .Y(\u_cpu.ALU.u_wallace._1765_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7453_  (.A(\u_cpu.ALU.u_wallace._1762_ ),
    .B(\u_cpu.ALU.u_wallace._1763_ ),
    .C(\u_cpu.ALU.u_wallace._1765_ ),
    .Y(\u_cpu.ALU.u_wallace._1766_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7454_  (.A(\u_cpu.ALU.SrcB[4] ),
    .B(\u_cpu.ALU.u_wallace._1486_ ),
    .C(\u_cpu.ALU.SrcA[17] ),
    .D(\u_cpu.ALU.SrcA[18] ),
    .Y(\u_cpu.ALU.u_wallace._1767_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7455_  (.A1(\u_cpu.ALU.u_wallace._1486_ ),
    .A2(\u_cpu.ALU.SrcA[17] ),
    .B1(\u_cpu.ALU.SrcA[18] ),
    .B2(\u_cpu.ALU.SrcB[4] ),
    .X(\u_cpu.ALU.u_wallace._1768_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7456_  (.A1_N(\u_cpu.ALU.u_wallace._1767_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1768_ ),
    .B1(\u_cpu.ALU.u_wallace._4470_ ),
    .B2(\u_cpu.ALU.u_wallace._1324_ ),
    .Y(\u_cpu.ALU.u_wallace._1769_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7457_  (.A(\u_cpu.ALU.u_wallace._1768_ ),
    .B(\u_cpu.ALU.u_wallace._0332_ ),
    .C(\u_cpu.ALU.SrcB[7] ),
    .D(\u_cpu.ALU.u_wallace._1767_ ),
    .Y(\u_cpu.ALU.u_wallace._1770_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7458_  (.A1(\u_cpu.ALU.u_wallace._0282_ ),
    .A2(\u_cpu.ALU.SrcA[19] ),
    .B1(\u_cpu.ALU.SrcA[20] ),
    .B2(\u_cpu.ALU.u_wallace._0195_ ),
    .Y(\u_cpu.ALU.u_wallace._1772_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7459_  (.A1(\u_cpu.ALU.u_wallace._1544_ ),
    .A2(\u_cpu.ALU.u_wallace._1772_ ),
    .B1(\u_cpu.ALU.u_wallace._1546_ ),
    .Y(\u_cpu.ALU.u_wallace._1773_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7460_  (.A(\u_cpu.ALU.u_wallace._1769_ ),
    .B(\u_cpu.ALU.u_wallace._1770_ ),
    .C(\u_cpu.ALU.u_wallace._1773_ ),
    .X(\u_cpu.ALU.u_wallace._1774_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7461_  (.A(\u_cpu.ALU.u_wallace._1774_ ),
    .X(\u_cpu.ALU.u_wallace._1775_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7462_  (.A1(\u_cpu.ALU.u_wallace._1769_ ),
    .A2(\u_cpu.ALU.u_wallace._1770_ ),
    .B1(\u_cpu.ALU.u_wallace._1773_ ),
    .X(\u_cpu.ALU.u_wallace._1776_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.ALU.u_wallace._7463_  (.A1_N(\u_cpu.ALU.u_wallace._0635_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1571_ ),
    .B1(\u_cpu.ALU.u_wallace._1575_ ),
    .B2(\u_cpu.ALU.u_wallace._1567_ ),
    .X(\u_cpu.ALU.u_wallace._1777_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7464_  (.A(\u_cpu.ALU.u_wallace._1776_ ),
    .B(\u_cpu.ALU.u_wallace._1777_ ),
    .Y(\u_cpu.ALU.u_wallace._1778_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7465_  (.A1(\u_cpu.ALU.u_wallace._1769_ ),
    .A2(\u_cpu.ALU.u_wallace._1770_ ),
    .B1(\u_cpu.ALU.u_wallace._1773_ ),
    .Y(\u_cpu.ALU.u_wallace._1779_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._7466_  (.A1(\u_cpu.ALU.u_wallace._1779_ ),
    .A2(\u_cpu.ALU.u_wallace._1775_ ),
    .B1_N(\u_cpu.ALU.u_wallace._1777_ ),
    .Y(\u_cpu.ALU.u_wallace._1780_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7467_  (.A1(\u_cpu.ALU.u_wallace._1775_ ),
    .A2(\u_cpu.ALU.u_wallace._1778_ ),
    .B1(\u_cpu.ALU.u_wallace._1780_ ),
    .Y(\u_cpu.ALU.u_wallace._1781_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7468_  (.A1(\u_cpu.ALU.u_wallace._1759_ ),
    .A2(\u_cpu.ALU.u_wallace._1766_ ),
    .B1(\u_cpu.ALU.u_wallace._1781_ ),
    .X(\u_cpu.ALU.u_wallace._1783_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7469_  (.A(\u_cpu.ALU.u_wallace._1769_ ),
    .B(\u_cpu.ALU.u_wallace._1770_ ),
    .C(\u_cpu.ALU.u_wallace._1773_ ),
    .Y(\u_cpu.ALU.u_wallace._1784_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7470_  (.A1(\u_cpu.ALU.u_wallace._1776_ ),
    .A2(\u_cpu.ALU.u_wallace._1784_ ),
    .B1(\u_cpu.ALU.u_wallace._1777_ ),
    .Y(\u_cpu.ALU.u_wallace._1785_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7471_  (.A(\u_cpu.ALU.u_wallace._1776_ ),
    .B(\u_cpu.ALU.u_wallace._1784_ ),
    .C(\u_cpu.ALU.u_wallace._1777_ ),
    .X(\u_cpu.ALU.u_wallace._1786_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7472_  (.A1(\u_cpu.ALU.u_wallace._1785_ ),
    .A2(\u_cpu.ALU.u_wallace._1786_ ),
    .B1(\u_cpu.ALU.u_wallace._1759_ ),
    .C1(\u_cpu.ALU.u_wallace._1766_ ),
    .Y(\u_cpu.ALU.u_wallace._1787_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._7473_  (.A1(\u_cpu.ALU.u_wallace._1566_ ),
    .A2(\u_cpu.ALU.u_wallace._1580_ ),
    .A3(\u_cpu.ALU.u_wallace._1583_ ),
    .B1(\u_cpu.ALU.u_wallace._1558_ ),
    .Y(\u_cpu.ALU.u_wallace._1788_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7474_  (.A(\u_cpu.ALU.u_wallace._1783_ ),
    .B(\u_cpu.ALU.u_wallace._1787_ ),
    .C(\u_cpu.ALU.u_wallace._1788_ ),
    .Y(\u_cpu.ALU.u_wallace._1789_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7475_  (.A1(\u_cpu.ALU.u_wallace._1721_ ),
    .A2(\u_cpu.ALU.u_wallace._1722_ ),
    .B1(\u_cpu.ALU.u_wallace._1789_ ),
    .Y(\u_cpu.ALU.u_wallace._1790_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7476_  (.A1(\u_cpu.ALU.u_wallace._1586_ ),
    .A2(\u_cpu.ALU.u_wallace._1584_ ),
    .B1(\u_cpu.ALU.u_wallace._1783_ ),
    .B2(\u_cpu.ALU.u_wallace._1787_ ),
    .Y(\u_cpu.ALU.u_wallace._1791_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7477_  (.A1(\u_cpu.ALU.u_wallace._1299_ ),
    .A2(\u_cpu.ALU.u_wallace._1327_ ),
    .B1(\u_cpu.ALU.u_wallace._1370_ ),
    .Y(\u_cpu.ALU.u_wallace._1792_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU.u_wallace._7478_  (.A1_N(\u_cpu.ALU.u_wallace._1586_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1566_ ),
    .B1(\u_cpu.ALU.u_wallace._1587_ ),
    .B2(\u_cpu.ALU.u_wallace._1588_ ),
    .X(\u_cpu.ALU.u_wallace._1794_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7479_  (.A(\u_cpu.ALU.u_wallace._1586_ ),
    .B(\u_cpu.ALU.u_wallace._1566_ ),
    .C(\u_cpu.ALU.u_wallace._1580_ ),
    .D(\u_cpu.ALU.u_wallace._1583_ ),
    .X(\u_cpu.ALU.u_wallace._1795_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7480_  (.A(\u_cpu.ALU.u_wallace._1598_ ),
    .B(\u_cpu.ALU.u_wallace._1599_ ),
    .Y(\u_cpu.ALU.u_wallace._1796_ ));
 sky130_fd_sc_hd__o32ai_2 \u_cpu.ALU.u_wallace._7481_  (.A1(\u_cpu.ALU.u_wallace._1792_ ),
    .A2(\u_cpu.ALU.u_wallace._1794_ ),
    .A3(\u_cpu.ALU.u_wallace._1795_ ),
    .B1(\u_cpu.ALU.u_wallace._1601_ ),
    .B2(\u_cpu.ALU.u_wallace._1796_ ),
    .Y(\u_cpu.ALU.u_wallace._1797_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7482_  (.A1(\u_cpu.ALU.u_wallace._1566_ ),
    .A2(\u_cpu.ALU.u_wallace._1580_ ),
    .A3(\u_cpu.ALU.u_wallace._1583_ ),
    .B1(\u_cpu.ALU.u_wallace._1558_ ),
    .X(\u_cpu.ALU.u_wallace._1798_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._7483_  (.A1(\u_cpu.ALU.u_wallace._1778_ ),
    .A2(\u_cpu.ALU.u_wallace._1775_ ),
    .B1(\u_cpu.ALU.u_wallace._1780_ ),
    .C1(\u_cpu.ALU.u_wallace._1759_ ),
    .D1(\u_cpu.ALU.u_wallace._1766_ ),
    .Y(\u_cpu.ALU.u_wallace._1799_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7484_  (.A(\u_cpu.ALU.u_wallace._1764_ ),
    .B(\u_cpu.ALU.u_wallace._1525_ ),
    .Y(\u_cpu.ALU.u_wallace._1800_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7485_  (.A(\u_cpu.ALU.u_wallace._1561_ ),
    .B(\u_cpu.ALU.u_wallace._1548_ ),
    .Y(\u_cpu.ALU.u_wallace._1801_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7486_  (.A1(\u_cpu.ALU.u_wallace._1800_ ),
    .A2(\u_cpu.ALU.u_wallace._1801_ ),
    .B1(\u_cpu.ALU.u_wallace._1762_ ),
    .B2(\u_cpu.ALU.u_wallace._1763_ ),
    .Y(\u_cpu.ALU.u_wallace._1802_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7487_  (.A1(\u_cpu.ALU.u_wallace._1748_ ),
    .A2(\u_cpu.ALU.u_wallace._1758_ ),
    .B1(\u_cpu.ALU.u_wallace._1723_ ),
    .Y(\u_cpu.ALU.u_wallace._1803_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7488_  (.A1(\u_cpu.ALU.u_wallace._1785_ ),
    .A2(\u_cpu.ALU.u_wallace._1786_ ),
    .B1(\u_cpu.ALU.u_wallace._1802_ ),
    .B2(\u_cpu.ALU.u_wallace._1803_ ),
    .Y(\u_cpu.ALU.u_wallace._1805_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7489_  (.A(\u_cpu.ALU.u_wallace._1798_ ),
    .B(\u_cpu.ALU.u_wallace._1799_ ),
    .C(\u_cpu.ALU.u_wallace._1805_ ),
    .Y(\u_cpu.ALU.u_wallace._1806_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._7490_  (.A1(\u_cpu.ALU.u_wallace._1715_ ),
    .A2(\u_cpu.ALU.u_wallace._1717_ ),
    .A3(\u_cpu.ALU.u_wallace._1718_ ),
    .B1(\u_cpu.ALU.u_wallace._1720_ ),
    .Y(\u_cpu.ALU.u_wallace._1807_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7491_  (.A(\u_cpu.ALU.u_wallace._1714_ ),
    .B(\u_cpu.ALU.u_wallace._1719_ ),
    .Y(\u_cpu.ALU.u_wallace._1808_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7492_  (.A1(\u_cpu.ALU.u_wallace._1714_ ),
    .A2(\u_cpu.ALU.u_wallace._1807_ ),
    .B1(\u_cpu.ALU.u_wallace._1808_ ),
    .B2(\u_cpu.ALU.u_wallace._1720_ ),
    .Y(\u_cpu.ALU.u_wallace._1809_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7493_  (.A1(\u_cpu.ALU.u_wallace._1806_ ),
    .A2(\u_cpu.ALU.u_wallace._1789_ ),
    .B1(\u_cpu.ALU.u_wallace._1809_ ),
    .X(\u_cpu.ALU.u_wallace._1810_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7494_  (.A1(\u_cpu.ALU.u_wallace._1790_ ),
    .A2(\u_cpu.ALU.u_wallace._1791_ ),
    .B1(\u_cpu.ALU.u_wallace._1797_ ),
    .C1(\u_cpu.ALU.u_wallace._1810_ ),
    .X(\u_cpu.ALU.u_wallace._1811_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7495_  (.A1(\u_cpu.ALU.u_wallace._1518_ ),
    .A2(\u_cpu.ALU.u_wallace._1515_ ),
    .B1(\u_cpu.ALU.u_wallace._1520_ ),
    .Y(\u_cpu.ALU.u_wallace._1812_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7496_  (.A(\u_cpu.ALU.SrcB[20] ),
    .Y(\u_cpu.ALU.u_wallace._1813_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7497_  (.A1(\u_cpu.ALU.u_wallace._4556_ ),
    .A2(\u_cpu.ALU.u_wallace._0957_ ),
    .B1(\u_cpu.ALU.SrcB[19] ),
    .B2(\u_cpu.ALU.u_wallace._2549_ ),
    .Y(\u_cpu.ALU.u_wallace._1814_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7498_  (.A(\u_cpu.ALU.u_wallace._4556_ ),
    .B(\u_cpu.ALU.u_wallace._2549_ ),
    .C(\u_cpu.ALU.u_wallace._0957_ ),
    .D(\u_cpu.ALU.SrcB[19] ),
    .X(\u_cpu.ALU.u_wallace._1816_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7499_  (.A1(\u_cpu.ALU.u_wallace._0403_ ),
    .A2(\u_cpu.ALU.u_wallace._1813_ ),
    .B1(\u_cpu.ALU.u_wallace._1814_ ),
    .B2(\u_cpu.ALU.u_wallace._1816_ ),
    .Y(\u_cpu.ALU.u_wallace._1817_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7500_  (.A(\u_cpu.ALU.u_wallace._1267_ ),
    .B(\u_cpu.ALU.u_wallace._1278_ ),
    .C(\u_cpu.ALU.u_wallace._1387_ ),
    .D(\u_cpu.ALU.u_wallace._1210_ ),
    .Y(\u_cpu.ALU.u_wallace._1818_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._7501_  (.A_N(\u_cpu.ALU.u_wallace._1814_ ),
    .B(\u_cpu.ALU.u_wallace._1818_ ),
    .C(\u_cpu.ALU.u_wallace._4597_ ),
    .D(\u_cpu.ALU.u_wallace._1386_ ),
    .Y(\u_cpu.ALU.u_wallace._1819_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7502_  (.A(\u_cpu.ALU.u_wallace._0392_ ),
    .B(\u_cpu.ALU.u_wallace._0764_ ),
    .C(\u_cpu.ALU.u_wallace._0957_ ),
    .D(\u_cpu.ALU.SrcB[19] ),
    .X(\u_cpu.ALU.u_wallace._1820_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7503_  (.A1(\u_cpu.ALU.u_wallace._1612_ ),
    .A2(\u_cpu.ALU.u_wallace._1386_ ),
    .A3(\u_cpu.ALU.u_wallace._0151_ ),
    .B1(\u_cpu.ALU.u_wallace._1820_ ),
    .X(\u_cpu.ALU.u_wallace._1821_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7504_  (.A1(\u_cpu.ALU.u_wallace._1817_ ),
    .A2(\u_cpu.ALU.u_wallace._1819_ ),
    .B1(\u_cpu.ALU.u_wallace._1821_ ),
    .X(\u_cpu.ALU.u_wallace._1822_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7505_  (.A(\u_cpu.ALU.u_wallace._1821_ ),
    .B(\u_cpu.ALU.u_wallace._1817_ ),
    .C(\u_cpu.ALU.u_wallace._1819_ ),
    .Y(\u_cpu.ALU.u_wallace._1823_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7506_  (.A(\u_cpu.ALU.SrcB[22] ),
    .X(\u_cpu.ALU.u_wallace._1824_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7507_  (.A(\u_cpu.ALU.u_wallace._0446_ ),
    .B(\u_cpu.ALU.u_wallace._1454_ ),
    .C(\u_cpu.ALU.SrcB[21] ),
    .X(\u_cpu.ALU.u_wallace._1825_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7508_  (.A1(\u_cpu.ALU.u_wallace._4463_ ),
    .A2(\u_cpu.ALU.SrcB[21] ),
    .B1(\u_cpu.ALU.SrcB[22] ),
    .B2(\u_cpu.ALU.u_wallace._0994_ ),
    .Y(\u_cpu.ALU.u_wallace._1827_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7509_  (.A1(\u_cpu.ALU.u_wallace._1824_ ),
    .A2(\u_cpu.ALU.u_wallace._1825_ ),
    .B1(\u_cpu.ALU.u_wallace._1827_ ),
    .Y(\u_cpu.ALU.u_wallace._1828_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7510_  (.A1(\u_cpu.ALU.u_wallace._1822_ ),
    .A2(\u_cpu.ALU.u_wallace._1823_ ),
    .B1(\u_cpu.ALU.u_wallace._1828_ ),
    .Y(\u_cpu.ALU.u_wallace._1829_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7511_  (.A(\u_cpu.ALU.u_wallace._1822_ ),
    .B(\u_cpu.ALU.u_wallace._1823_ ),
    .C(\u_cpu.ALU.u_wallace._1828_ ),
    .X(\u_cpu.ALU.u_wallace._1830_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7512_  (.A1(\u_cpu.ALU.u_wallace._3645_ ),
    .A2(\u_cpu.ALU.SrcB[14] ),
    .B1(\u_cpu.ALU.u_wallace._0278_ ),
    .B2(\u_cpu.ALU.u_wallace._2878_ ),
    .Y(\u_cpu.ALU.u_wallace._1831_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7513_  (.A(\u_cpu.ALU.SrcA[8] ),
    .B(\u_cpu.ALU.SrcA[7] ),
    .C(\u_cpu.ALU.SrcB[14] ),
    .D(\u_cpu.ALU.SrcB[15] ),
    .X(\u_cpu.ALU.u_wallace._1832_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7514_  (.A1(\u_cpu.ALU.u_wallace._4454_ ),
    .A2(\u_cpu.ALU.u_wallace._0553_ ),
    .B1(\u_cpu.ALU.u_wallace._1831_ ),
    .B2(\u_cpu.ALU.u_wallace._1832_ ),
    .Y(\u_cpu.ALU.u_wallace._1833_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7515_  (.A1(\u_cpu.ALU.SrcA[8] ),
    .A2(\u_cpu.ALU.SrcB[14] ),
    .B1(\u_cpu.ALU.SrcB[15] ),
    .B2(\u_cpu.ALU.SrcA[7] ),
    .X(\u_cpu.ALU.u_wallace._1834_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7516_  (.A(\u_cpu.ALU.u_wallace._3645_ ),
    .B(\u_cpu.ALU.u_wallace._2878_ ),
    .C(\u_cpu.ALU.SrcB[14] ),
    .D(\u_cpu.ALU.u_wallace._0278_ ),
    .Y(\u_cpu.ALU.u_wallace._1835_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7517_  (.A(\u_cpu.ALU.u_wallace._1834_ ),
    .B(\u_cpu.ALU.u_wallace._1835_ ),
    .C(\u_cpu.ALU.u_wallace._3777_ ),
    .D(\u_cpu.ALU.u_wallace._0550_ ),
    .Y(\u_cpu.ALU.u_wallace._1836_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7518_  (.A(\u_cpu.ALU.u_wallace._3645_ ),
    .B(\u_cpu.ALU.SrcB[13] ),
    .Y(\u_cpu.ALU.u_wallace._1838_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7519_  (.A1(\u_cpu.ALU.u_wallace._1838_ ),
    .A2(\u_cpu.ALU.u_wallace._1490_ ),
    .B1(\u_cpu.ALU.u_wallace._1510_ ),
    .Y(\u_cpu.ALU.u_wallace._1839_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7520_  (.A1(\u_cpu.ALU.u_wallace._1833_ ),
    .A2(\u_cpu.ALU.u_wallace._1836_ ),
    .B1(\u_cpu.ALU.u_wallace._1839_ ),
    .Y(\u_cpu.ALU.u_wallace._1840_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7521_  (.A(\u_cpu.ALU.u_wallace._1833_ ),
    .B(\u_cpu.ALU.u_wallace._1836_ ),
    .C(\u_cpu.ALU.u_wallace._1839_ ),
    .X(\u_cpu.ALU.u_wallace._1841_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._7522_  (.A1(\u_cpu.ALU.u_wallace._4813_ ),
    .A2(\u_cpu.ALU.u_wallace._0941_ ),
    .A3(\u_cpu.ALU.u_wallace._1624_ ),
    .B1(\u_cpu.ALU.u_wallace._1628_ ),
    .X(\u_cpu.ALU.u_wallace._1842_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7523_  (.A1(\u_cpu.ALU.u_wallace._1840_ ),
    .A2(\u_cpu.ALU.u_wallace._1841_ ),
    .B1(\u_cpu.ALU.u_wallace._1842_ ),
    .Y(\u_cpu.ALU.u_wallace._1843_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7524_  (.A(\u_cpu.ALU.u_wallace._1833_ ),
    .B(\u_cpu.ALU.u_wallace._1836_ ),
    .C(\u_cpu.ALU.u_wallace._1839_ ),
    .Y(\u_cpu.ALU.u_wallace._1844_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7525_  (.A1(\u_cpu.ALU.u_wallace._1627_ ),
    .A2(\u_cpu.ALU.u_wallace._0735_ ),
    .A3(\u_cpu.ALU.u_wallace._1136_ ),
    .B1(\u_cpu.ALU.u_wallace._1625_ ),
    .X(\u_cpu.ALU.u_wallace._1845_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._7526_  (.A_N(\u_cpu.ALU.u_wallace._1840_ ),
    .B(\u_cpu.ALU.u_wallace._1844_ ),
    .C(\u_cpu.ALU.u_wallace._1845_ ),
    .Y(\u_cpu.ALU.u_wallace._1846_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7527_  (.A1(\u_cpu.ALU.u_wallace._1635_ ),
    .A2(\u_cpu.ALU.u_wallace._1633_ ),
    .B1(\u_cpu.ALU.u_wallace._1638_ ),
    .Y(\u_cpu.ALU.u_wallace._1847_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7528_  (.A1(\u_cpu.ALU.u_wallace._1843_ ),
    .A2(\u_cpu.ALU.u_wallace._1846_ ),
    .B1(\u_cpu.ALU.u_wallace._1847_ ),
    .Y(\u_cpu.ALU.u_wallace._1849_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7529_  (.A(\u_cpu.ALU.u_wallace._1635_ ),
    .B(\u_cpu.ALU.u_wallace._1633_ ),
    .Y(\u_cpu.ALU.u_wallace._1850_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7530_  (.A1(\u_cpu.ALU.u_wallace._1634_ ),
    .A2(\u_cpu.ALU.u_wallace._1850_ ),
    .B1(\u_cpu.ALU.u_wallace._1843_ ),
    .C1(\u_cpu.ALU.u_wallace._1846_ ),
    .X(\u_cpu.ALU.u_wallace._1851_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7531_  (.A1(\u_cpu.ALU.u_wallace._1829_ ),
    .A2(\u_cpu.ALU.u_wallace._1830_ ),
    .B1(\u_cpu.ALU.u_wallace._1849_ ),
    .B2(\u_cpu.ALU.u_wallace._1851_ ),
    .Y(\u_cpu.ALU.u_wallace._1852_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7532_  (.A1(\u_cpu.ALU.u_wallace._1843_ ),
    .A2(\u_cpu.ALU.u_wallace._1846_ ),
    .B1(\u_cpu.ALU.u_wallace._1847_ ),
    .X(\u_cpu.ALU.u_wallace._1853_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7533_  (.A1(\u_cpu.ALU.u_wallace._1634_ ),
    .A2(\u_cpu.ALU.u_wallace._1850_ ),
    .B1(\u_cpu.ALU.u_wallace._1843_ ),
    .C1(\u_cpu.ALU.u_wallace._1846_ ),
    .Y(\u_cpu.ALU.u_wallace._1854_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7534_  (.A(\u_cpu.ALU.u_wallace._1824_ ),
    .X(\u_cpu.ALU.u_wallace._1855_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7535_  (.A1(\u_cpu.ALU.u_wallace._1817_ ),
    .A2(\u_cpu.ALU.u_wallace._1819_ ),
    .B1(\u_cpu.ALU.u_wallace._1821_ ),
    .Y(\u_cpu.ALU.u_wallace._1856_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU.u_wallace._7536_  (.A1(\u_cpu.ALU.u_wallace._1855_ ),
    .A2(\u_cpu.ALU.u_wallace._1825_ ),
    .B1(\u_cpu.ALU.u_wallace._1827_ ),
    .C1(\u_cpu.ALU.u_wallace._1856_ ),
    .Y(\u_cpu.ALU.u_wallace._1857_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7537_  (.A1(\u_cpu.ALU.u_wallace._1857_ ),
    .A2(\u_cpu.ALU.u_wallace._1823_ ),
    .B1(\u_cpu.ALU.u_wallace._1829_ ),
    .Y(\u_cpu.ALU.u_wallace._1858_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7538_  (.A(\u_cpu.ALU.u_wallace._1853_ ),
    .B(\u_cpu.ALU.u_wallace._1854_ ),
    .C(\u_cpu.ALU.u_wallace._1858_ ),
    .Y(\u_cpu.ALU.u_wallace._1860_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7539_  (.A(\u_cpu.ALU.u_wallace._1812_ ),
    .B(\u_cpu.ALU.u_wallace._1852_ ),
    .C(\u_cpu.ALU.u_wallace._1860_ ),
    .Y(\u_cpu.ALU.u_wallace._1861_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7540_  (.A(\u_cpu.ALU.u_wallace._1861_ ),
    .Y(\u_cpu.ALU.u_wallace._1862_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7541_  (.A1(\u_cpu.ALU.u_wallace._1852_ ),
    .A2(\u_cpu.ALU.u_wallace._1860_ ),
    .B1(\u_cpu.ALU.u_wallace._1812_ ),
    .X(\u_cpu.ALU.u_wallace._1863_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7542_  (.A1(\u_cpu.ALU.u_wallace._1622_ ),
    .A2(\u_cpu.ALU.u_wallace._1623_ ),
    .A3(\u_cpu.ALU.u_wallace._1645_ ),
    .B1(\u_cpu.ALU.u_wallace._1643_ ),
    .X(\u_cpu.ALU.u_wallace._1864_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7543_  (.A(\u_cpu.ALU.u_wallace._1863_ ),
    .B(\u_cpu.ALU.u_wallace._1864_ ),
    .Y(\u_cpu.ALU.u_wallace._1865_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7544_  (.A1(\u_cpu.ALU.u_wallace._1863_ ),
    .A2(\u_cpu.ALU.u_wallace._1861_ ),
    .B1(\u_cpu.ALU.u_wallace._1864_ ),
    .X(\u_cpu.ALU.u_wallace._1866_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.ALU.u_wallace._7545_  (.A1(\u_cpu.ALU.u_wallace._1792_ ),
    .A2(\u_cpu.ALU.u_wallace._1794_ ),
    .A3(\u_cpu.ALU.u_wallace._1795_ ),
    .B1(\u_cpu.ALU.u_wallace._1601_ ),
    .B2(\u_cpu.ALU.u_wallace._1796_ ),
    .X(\u_cpu.ALU.u_wallace._1867_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7546_  (.A1(\u_cpu.ALU.u_wallace._1799_ ),
    .A2(\u_cpu.ALU.u_wallace._1805_ ),
    .B1(\u_cpu.ALU.u_wallace._1798_ ),
    .Y(\u_cpu.ALU.u_wallace._1868_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7547_  (.A1(\u_cpu.ALU.u_wallace._1721_ ),
    .A2(\u_cpu.ALU.u_wallace._1722_ ),
    .B1(\u_cpu.ALU.u_wallace._1791_ ),
    .B2(\u_cpu.ALU.u_wallace._1868_ ),
    .Y(\u_cpu.ALU.u_wallace._1869_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._7548_  (.A_N(\u_cpu.ALU.u_wallace._1809_ ),
    .B(\u_cpu.ALU.u_wallace._1806_ ),
    .C(\u_cpu.ALU.u_wallace._1789_ ),
    .Y(\u_cpu.ALU.u_wallace._1871_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7549_  (.A(\u_cpu.ALU.u_wallace._1867_ ),
    .B(\u_cpu.ALU.u_wallace._1869_ ),
    .C(\u_cpu.ALU.u_wallace._1871_ ),
    .Y(\u_cpu.ALU.u_wallace._1872_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7550_  (.A1(\u_cpu.ALU.u_wallace._1862_ ),
    .A2(\u_cpu.ALU.u_wallace._1865_ ),
    .B1(\u_cpu.ALU.u_wallace._1866_ ),
    .C1(\u_cpu.ALU.u_wallace._1872_ ),
    .Y(\u_cpu.ALU.u_wallace._1873_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7551_  (.A1(\u_cpu.ALU.u_wallace._1790_ ),
    .A2(\u_cpu.ALU.u_wallace._1791_ ),
    .B1(\u_cpu.ALU.u_wallace._1797_ ),
    .C1(\u_cpu.ALU.u_wallace._1810_ ),
    .Y(\u_cpu.ALU.u_wallace._1874_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7552_  (.A1(\u_cpu.ALU.u_wallace._1863_ ),
    .A2(\u_cpu.ALU.u_wallace._1861_ ),
    .B1(\u_cpu.ALU.u_wallace._1864_ ),
    .Y(\u_cpu.ALU.u_wallace._1875_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7553_  (.A(\u_cpu.ALU.u_wallace._1863_ ),
    .B(\u_cpu.ALU.u_wallace._1861_ ),
    .C(\u_cpu.ALU.u_wallace._1864_ ),
    .Y(\u_cpu.ALU.u_wallace._1876_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7554_  (.A(\u_cpu.ALU.u_wallace._1876_ ),
    .Y(\u_cpu.ALU.u_wallace._1877_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7555_  (.A1_N(\u_cpu.ALU.u_wallace._1874_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1872_ ),
    .B1(\u_cpu.ALU.u_wallace._1875_ ),
    .B2(\u_cpu.ALU.u_wallace._1877_ ),
    .Y(\u_cpu.ALU.u_wallace._1878_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7556_  (.A(\u_cpu.ALU.u_wallace._1658_ ),
    .B(\u_cpu.ALU.u_wallace._1657_ ),
    .Y(\u_cpu.ALU.u_wallace._1879_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7557_  (.A1(\u_cpu.ALU.u_wallace._1811_ ),
    .A2(\u_cpu.ALU.u_wallace._1873_ ),
    .B1(\u_cpu.ALU.u_wallace._1878_ ),
    .C1(\u_cpu.ALU.u_wallace._1879_ ),
    .Y(\u_cpu.ALU.u_wallace._1880_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._7558_  (.A1(\u_cpu.ALU.u_wallace._1862_ ),
    .A2(\u_cpu.ALU.u_wallace._1865_ ),
    .B1(\u_cpu.ALU.u_wallace._1866_ ),
    .C1(\u_cpu.ALU.u_wallace._1874_ ),
    .D1(\u_cpu.ALU.u_wallace._1872_ ),
    .X(\u_cpu.ALU.u_wallace._1882_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7559_  (.A1(\u_cpu.ALU.u_wallace._1874_ ),
    .A2(\u_cpu.ALU.u_wallace._1872_ ),
    .B1(\u_cpu.ALU.u_wallace._1866_ ),
    .B2(\u_cpu.ALU.u_wallace._1876_ ),
    .Y(\u_cpu.ALU.u_wallace._1883_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._7560_  (.A1(\u_cpu.ALU.u_wallace._1609_ ),
    .A2(\u_cpu.ALU.u_wallace._1652_ ),
    .A3(\u_cpu.ALU.u_wallace._1656_ ),
    .B1(\u_cpu.ALU.u_wallace._1603_ ),
    .Y(\u_cpu.ALU.u_wallace._1884_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7561_  (.A1(\u_cpu.ALU.u_wallace._1882_ ),
    .A2(\u_cpu.ALU.u_wallace._1883_ ),
    .B1(\u_cpu.ALU.u_wallace._1884_ ),
    .Y(\u_cpu.ALU.u_wallace._1885_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7562_  (.A(\u_cpu.ALU.u_wallace._0129_ ),
    .X(\u_cpu.ALU.u_wallace._1886_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7563_  (.A(\u_cpu.ALU.u_wallace._1619_ ),
    .B(\u_cpu.ALU.u_wallace._1614_ ),
    .C(\u_cpu.ALU.u_wallace._1616_ ),
    .X(\u_cpu.ALU.u_wallace._1887_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7564_  (.A1(\u_cpu.ALU.u_wallace._1620_ ),
    .A2(\u_cpu.ALU.u_wallace._1611_ ),
    .A3(\u_cpu.ALU.u_wallace._1886_ ),
    .B1(\u_cpu.ALU.u_wallace._1887_ ),
    .X(\u_cpu.ALU.u_wallace._1888_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7565_  (.A(\u_cpu.ALU.u_wallace._1888_ ),
    .Y(\u_cpu.ALU.u_wallace._1889_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7566_  (.A1(\u_cpu.ALU.u_wallace._1650_ ),
    .A2(\u_cpu.ALU.u_wallace._1652_ ),
    .B1(\u_cpu.ALU.u_wallace._1889_ ),
    .X(\u_cpu.ALU.u_wallace._1890_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7567_  (.A(\u_cpu.ALU.u_wallace._1890_ ),
    .Y(\u_cpu.ALU.u_wallace._1891_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7568_  (.A(\u_cpu.ALU.u_wallace._1650_ ),
    .B(\u_cpu.ALU.u_wallace._1652_ ),
    .C(\u_cpu.ALU.u_wallace._1889_ ),
    .X(\u_cpu.ALU.u_wallace._1893_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7569_  (.A1_N(\u_cpu.ALU.u_wallace._1880_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1885_ ),
    .B1(\u_cpu.ALU.u_wallace._1891_ ),
    .B2(\u_cpu.ALU.u_wallace._1893_ ),
    .Y(\u_cpu.ALU.u_wallace._1894_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7570_  (.A1(\u_cpu.ALU.u_wallace._1650_ ),
    .A2(\u_cpu.ALU.u_wallace._1652_ ),
    .B1(\u_cpu.ALU.u_wallace._1888_ ),
    .Y(\u_cpu.ALU.u_wallace._1895_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7571_  (.A(\u_cpu.ALU.u_wallace._1650_ ),
    .B(\u_cpu.ALU.u_wallace._1652_ ),
    .C(\u_cpu.ALU.u_wallace._1888_ ),
    .X(\u_cpu.ALU.u_wallace._1896_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7572_  (.A1(\u_cpu.ALU.u_wallace._1895_ ),
    .A2(\u_cpu.ALU.u_wallace._1896_ ),
    .B1(\u_cpu.ALU.u_wallace._1880_ ),
    .C1(\u_cpu.ALU.u_wallace._1885_ ),
    .Y(\u_cpu.ALU.u_wallace._1897_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7573_  (.A(\u_cpu.ALU.u_wallace._1661_ ),
    .B(\u_cpu.ALU.u_wallace._1482_ ),
    .Y(\u_cpu.ALU.u_wallace._1898_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7574_  (.A1(\u_cpu.ALU.u_wallace._1676_ ),
    .A2(\u_cpu.ALU.u_wallace._1670_ ),
    .B1(\u_cpu.ALU.u_wallace._1898_ ),
    .Y(\u_cpu.ALU.u_wallace._1899_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7575_  (.A1(\u_cpu.ALU.u_wallace._1894_ ),
    .A2(\u_cpu.ALU.u_wallace._1897_ ),
    .B1(\u_cpu.ALU.u_wallace._1899_ ),
    .X(\u_cpu.ALU.u_wallace._1900_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7576_  (.A1(\u_cpu.ALU.u_wallace._1811_ ),
    .A2(\u_cpu.ALU.u_wallace._1873_ ),
    .B1(\u_cpu.ALU.u_wallace._1878_ ),
    .C1(\u_cpu.ALU.u_wallace._1879_ ),
    .X(\u_cpu.ALU.u_wallace._1901_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7577_  (.A1(\u_cpu.ALU.u_wallace._1811_ ),
    .A2(\u_cpu.ALU.u_wallace._1873_ ),
    .B1(\u_cpu.ALU.u_wallace._1878_ ),
    .Y(\u_cpu.ALU.u_wallace._1902_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.ALU.u_wallace._7578_  (.A1_N(\u_cpu.ALU.u_wallace._1895_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1896_ ),
    .B1(\u_cpu.ALU.u_wallace._1884_ ),
    .B2(\u_cpu.ALU.u_wallace._1902_ ),
    .X(\u_cpu.ALU.u_wallace._1904_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7579_  (.A1(\u_cpu.ALU.u_wallace._1901_ ),
    .A2(\u_cpu.ALU.u_wallace._1904_ ),
    .B1(\u_cpu.ALU.u_wallace._1894_ ),
    .C1(\u_cpu.ALU.u_wallace._1899_ ),
    .Y(\u_cpu.ALU.u_wallace._1905_ ));
 sky130_fd_sc_hd__a2111o_2 \u_cpu.ALU.u_wallace._7580_  (.A1(\u_cpu.ALU.u_wallace._1427_ ),
    .A2(\u_cpu.ALU.u_wallace._1434_ ),
    .B1(\u_cpu.ALU.u_wallace._1179_ ),
    .C1(\u_cpu.ALU.u_wallace._1177_ ),
    .D1(\u_cpu.ALU.u_wallace._1422_ ),
    .X(\u_cpu.ALU.u_wallace._1906_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7581_  (.A(\u_cpu.ALU.u_wallace._1906_ ),
    .Y(\u_cpu.ALU.u_wallace._1907_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7582_  (.A1(\u_cpu.ALU.u_wallace._1900_ ),
    .A2(\u_cpu.ALU.u_wallace._1905_ ),
    .B1(\u_cpu.ALU.u_wallace._1907_ ),
    .Y(\u_cpu.ALU.u_wallace._1908_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._7583_  (.A1(\u_cpu.ALU.u_wallace._1428_ ),
    .A2(\u_cpu.ALU.u_wallace._1448_ ),
    .B1(\u_cpu.ALU.u_wallace._1905_ ),
    .C1(\u_cpu.ALU.u_wallace._1394_ ),
    .D1(\u_cpu.ALU.u_wallace._1900_ ),
    .X(\u_cpu.ALU.u_wallace._1909_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7584_  (.A1(\u_cpu.ALU.u_wallace._1680_ ),
    .A2(\u_cpu.ALU.u_wallace._1689_ ),
    .B1(\u_cpu.ALU.u_wallace._1908_ ),
    .B2(\u_cpu.ALU.u_wallace._1909_ ),
    .Y(\u_cpu.ALU.u_wallace._1910_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7585_  (.A1(\u_cpu.ALU.u_wallace._1894_ ),
    .A2(\u_cpu.ALU.u_wallace._1897_ ),
    .B1(\u_cpu.ALU.u_wallace._1899_ ),
    .Y(\u_cpu.ALU.u_wallace._1911_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7586_  (.A1(\u_cpu.ALU.u_wallace._1901_ ),
    .A2(\u_cpu.ALU.u_wallace._1904_ ),
    .B1(\u_cpu.ALU.u_wallace._1894_ ),
    .C1(\u_cpu.ALU.u_wallace._1899_ ),
    .X(\u_cpu.ALU.u_wallace._1912_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7587_  (.A1(\u_cpu.ALU.u_wallace._1911_ ),
    .A2(\u_cpu.ALU.u_wallace._1912_ ),
    .B1(\u_cpu.ALU.u_wallace._1906_ ),
    .Y(\u_cpu.ALU.u_wallace._1913_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._7588_  (.A1(\u_cpu.ALU.u_wallace._1428_ ),
    .A2(\u_cpu.ALU.u_wallace._1448_ ),
    .B1(\u_cpu.ALU.u_wallace._1905_ ),
    .C1(\u_cpu.ALU.u_wallace._1394_ ),
    .D1(\u_cpu.ALU.u_wallace._1900_ ),
    .Y(\u_cpu.ALU.u_wallace._1915_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._7589_  (.A1(\u_cpu.ALU.u_wallace._1457_ ),
    .A2(\u_cpu.ALU.u_wallace._1681_ ),
    .B1(\u_cpu.ALU.u_wallace._1913_ ),
    .C1(\u_cpu.ALU.u_wallace._1915_ ),
    .D1(\u_cpu.ALU.u_wallace._1674_ ),
    .Y(\u_cpu.ALU.u_wallace._1916_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7590_  (.A(\u_cpu.ALU.u_wallace._1910_ ),
    .B(\u_cpu.ALU.u_wallace._1916_ ),
    .Y(\u_cpu.ALU.u_wallace._1917_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7591_  (.A1(\u_cpu.ALU.u_wallace._1254_ ),
    .A2(\u_cpu.ALU.u_wallace._1453_ ),
    .A3(\u_cpu.ALU.u_wallace._1456_ ),
    .B1(\u_cpu.ALU.u_wallace._1478_ ),
    .X(\u_cpu.ALU.u_wallace._1918_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7592_  (.A(\u_cpu.ALU.u_wallace._1674_ ),
    .B(\u_cpu.ALU.u_wallace._1678_ ),
    .Y(\u_cpu.ALU.u_wallace._1919_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7593_  (.A1_N(\u_cpu.ALU.u_wallace._1683_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1686_ ),
    .B1(\u_cpu.ALU.u_wallace._1918_ ),
    .B2(\u_cpu.ALU.u_wallace._1919_ ),
    .Y(\u_cpu.ALU.u_wallace._1920_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._7594_  (.A(\u_cpu.ALU.u_wallace._1917_ ),
    .B(\u_cpu.ALU.u_wallace._1920_ ),
    .X(\u_cpu.ALU.Product_Wallace[22] ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._7595_  (.A1_N(\u_cpu.ALU.u_wallace._1895_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1896_ ),
    .B1(\u_cpu.ALU.u_wallace._1884_ ),
    .B2(\u_cpu.ALU.u_wallace._1902_ ),
    .Y(\u_cpu.ALU.u_wallace._1921_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._7596_  (.A1(\u_cpu.ALU.u_wallace._1712_ ),
    .A2(\u_cpu.ALU.u_wallace._1711_ ),
    .B1(\u_cpu.ALU.u_wallace._1706_ ),
    .X(\u_cpu.ALU.u_wallace._1922_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7597_  (.A(\u_cpu.ALU.SrcB[8] ),
    .B(\u_cpu.ALU.SrcB[9] ),
    .C(\u_cpu.ALU.SrcA[14] ),
    .D(\u_cpu.ALU.SrcA[15] ),
    .Y(\u_cpu.ALU.u_wallace._1923_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7598_  (.A1(\u_cpu.ALU.SrcB[9] ),
    .A2(\u_cpu.ALU.SrcA[14] ),
    .B1(\u_cpu.ALU.SrcA[15] ),
    .B2(\u_cpu.ALU.SrcB[8] ),
    .X(\u_cpu.ALU.u_wallace._1925_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7599_  (.A1_N(\u_cpu.ALU.u_wallace._1923_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1925_ ),
    .B1(\u_cpu.ALU.u_wallace._4601_ ),
    .B2(\u_cpu.ALU.u_wallace._0458_ ),
    .Y(\u_cpu.ALU.u_wallace._1926_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7600_  (.A(\u_cpu.ALU.u_wallace._1925_ ),
    .B(\u_cpu.ALU.u_wallace._4921_ ),
    .C(\u_cpu.ALU.u_wallace._0041_ ),
    .D(\u_cpu.ALU.u_wallace._1923_ ),
    .Y(\u_cpu.ALU.u_wallace._1927_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7601_  (.A1(\u_cpu.ALU.u_wallace._1698_ ),
    .A2(\u_cpu.ALU.u_wallace._1697_ ),
    .B1(\u_cpu.ALU.u_wallace._1702_ ),
    .Y(\u_cpu.ALU.u_wallace._1928_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7602_  (.A1(\u_cpu.ALU.u_wallace._1926_ ),
    .A2(\u_cpu.ALU.u_wallace._1927_ ),
    .B1(\u_cpu.ALU.u_wallace._1928_ ),
    .Y(\u_cpu.ALU.u_wallace._1929_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7603_  (.A1(\u_cpu.ALU.u_wallace._4836_ ),
    .A2(\u_cpu.ALU.u_wallace._4790_ ),
    .B1(\u_cpu.ALU.u_wallace._4841_ ),
    .B2(\u_cpu.ALU.u_wallace._4650_ ),
    .X(\u_cpu.ALU.u_wallace._1930_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7604_  (.A(\u_cpu.ALU.u_wallace._4647_ ),
    .B(\u_cpu.ALU.u_wallace._0364_ ),
    .C(\u_cpu.ALU.u_wallace._4900_ ),
    .D(\u_cpu.ALU.u_wallace._4841_ ),
    .Y(\u_cpu.ALU.u_wallace._1931_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7605_  (.A(\u_cpu.ALU.u_wallace._4551_ ),
    .B(\u_cpu.ALU.SrcB[13] ),
    .Y(\u_cpu.ALU.u_wallace._1932_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7606_  (.A1(\u_cpu.ALU.u_wallace._1930_ ),
    .A2(\u_cpu.ALU.u_wallace._1931_ ),
    .B1(\u_cpu.ALU.u_wallace._1932_ ),
    .Y(\u_cpu.ALU.u_wallace._1933_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7607_  (.A(\u_cpu.ALU.u_wallace._1932_ ),
    .B(\u_cpu.ALU.u_wallace._1930_ ),
    .C(\u_cpu.ALU.u_wallace._1931_ ),
    .X(\u_cpu.ALU.u_wallace._1934_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7608_  (.A(\u_cpu.ALU.u_wallace._4716_ ),
    .B(\u_cpu.ALU.u_wallace._4598_ ),
    .C(\u_cpu.ALU.u_wallace._4909_ ),
    .D(\u_cpu.ALU.u_wallace._0177_ ),
    .X(\u_cpu.ALU.u_wallace._1936_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7609_  (.A(\u_cpu.ALU.u_wallace._1698_ ),
    .B(\u_cpu.ALU.u_wallace._1697_ ),
    .Y(\u_cpu.ALU.u_wallace._1937_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7610_  (.A1(\u_cpu.ALU.u_wallace._1936_ ),
    .A2(\u_cpu.ALU.u_wallace._1937_ ),
    .B1(\u_cpu.ALU.u_wallace._1926_ ),
    .C1(\u_cpu.ALU.u_wallace._1927_ ),
    .Y(\u_cpu.ALU.u_wallace._1938_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7611_  (.A1(\u_cpu.ALU.u_wallace._1933_ ),
    .A2(\u_cpu.ALU.u_wallace._1934_ ),
    .B1(\u_cpu.ALU.u_wallace._1938_ ),
    .Y(\u_cpu.ALU.u_wallace._1939_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7612_  (.A(\u_cpu.ALU.u_wallace._1769_ ),
    .B(\u_cpu.ALU.u_wallace._1770_ ),
    .Y(\u_cpu.ALU.u_wallace._1940_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._7613_  (.A1(\u_cpu.ALU.u_wallace._1892_ ),
    .A2(\u_cpu.ALU.u_wallace._0809_ ),
    .A3(\u_cpu.ALU.u_wallace._1772_ ),
    .B1(\u_cpu.ALU.u_wallace._1546_ ),
    .X(\u_cpu.ALU.u_wallace._1941_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._7614_  (.A1(\u_cpu.ALU.u_wallace._1940_ ),
    .A2(\u_cpu.ALU.u_wallace._1941_ ),
    .B1_N(\u_cpu.ALU.u_wallace._1777_ ),
    .Y(\u_cpu.ALU.u_wallace._1942_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7615_  (.A1(\u_cpu.ALU.u_wallace._0364_ ),
    .A2(\u_cpu.ALU.u_wallace._4785_ ),
    .B1(\u_cpu.ALU.u_wallace._0365_ ),
    .B2(\u_cpu.ALU.u_wallace._4647_ ),
    .Y(\u_cpu.ALU.u_wallace._1943_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7616_  (.A(\u_cpu.ALU.u_wallace._4650_ ),
    .B(\u_cpu.ALU.u_wallace._4836_ ),
    .C(\u_cpu.ALU.u_wallace._4790_ ),
    .D(\u_cpu.ALU.SrcB[12] ),
    .X(\u_cpu.ALU.u_wallace._1944_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._7617_  (.A1(\u_cpu.ALU.u_wallace._4904_ ),
    .A2(\u_cpu.ALU.u_wallace._0036_ ),
    .B1(\u_cpu.ALU.u_wallace._1943_ ),
    .B2(\u_cpu.ALU.u_wallace._1944_ ),
    .X(\u_cpu.ALU.u_wallace._1945_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7618_  (.A(\u_cpu.ALU.u_wallace._1930_ ),
    .B(\u_cpu.ALU.u_wallace._1931_ ),
    .C(\u_cpu.ALU.u_wallace._4554_ ),
    .D(\u_cpu.ALU.u_wallace._0033_ ),
    .X(\u_cpu.ALU.u_wallace._1947_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7619_  (.A1(\u_cpu.ALU.u_wallace._1936_ ),
    .A2(\u_cpu.ALU.u_wallace._1937_ ),
    .B1(\u_cpu.ALU.u_wallace._1926_ ),
    .C1(\u_cpu.ALU.u_wallace._1927_ ),
    .X(\u_cpu.ALU.u_wallace._1948_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7620_  (.A1(\u_cpu.ALU.u_wallace._1945_ ),
    .A2(\u_cpu.ALU.u_wallace._1947_ ),
    .B1(\u_cpu.ALU.u_wallace._1929_ ),
    .B2(\u_cpu.ALU.u_wallace._1948_ ),
    .Y(\u_cpu.ALU.u_wallace._1949_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._7621_  (.A1(\u_cpu.ALU.u_wallace._1929_ ),
    .A2(\u_cpu.ALU.u_wallace._1939_ ),
    .B1(\u_cpu.ALU.u_wallace._1775_ ),
    .B2(\u_cpu.ALU.u_wallace._1942_ ),
    .C1(\u_cpu.ALU.u_wallace._1949_ ),
    .X(\u_cpu.ALU.u_wallace._1950_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7622_  (.A(\u_cpu.ALU.u_wallace._1950_ ),
    .X(\u_cpu.ALU.u_wallace._1951_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7623_  (.A1(\u_cpu.ALU.u_wallace._1926_ ),
    .A2(\u_cpu.ALU.u_wallace._1927_ ),
    .B1(\u_cpu.ALU.u_wallace._1928_ ),
    .X(\u_cpu.ALU.u_wallace._1952_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7624_  (.A1(\u_cpu.ALU.u_wallace._1933_ ),
    .A2(\u_cpu.ALU.u_wallace._1934_ ),
    .B1(\u_cpu.ALU.u_wallace._1952_ ),
    .C1(\u_cpu.ALU.u_wallace._1938_ ),
    .Y(\u_cpu.ALU.u_wallace._1953_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7625_  (.A1(\u_cpu.ALU.u_wallace._1776_ ),
    .A2(\u_cpu.ALU.u_wallace._1777_ ),
    .B1(\u_cpu.ALU.u_wallace._1775_ ),
    .X(\u_cpu.ALU.u_wallace._1954_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7626_  (.A1(\u_cpu.ALU.u_wallace._1953_ ),
    .A2(\u_cpu.ALU.u_wallace._1949_ ),
    .B1(\u_cpu.ALU.u_wallace._1954_ ),
    .Y(\u_cpu.ALU.u_wallace._1955_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._7627_  (.A(\u_cpu.ALU.u_wallace._1922_ ),
    .B(\u_cpu.ALU.u_wallace._1951_ ),
    .C(\u_cpu.ALU.u_wallace._1955_ ),
    .Y(\u_cpu.ALU.u_wallace._1956_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._7628_  (.A1(\u_cpu.ALU.u_wallace._1951_ ),
    .A2(\u_cpu.ALU.u_wallace._1955_ ),
    .B1(\u_cpu.ALU.u_wallace._1922_ ),
    .X(\u_cpu.ALU.u_wallace._1958_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7629_  (.A1(\u_cpu.ALU.u_wallace._2538_ ),
    .A2(\u_cpu.ALU.u_wallace._1084_ ),
    .B1(\u_cpu.ALU.u_wallace._1100_ ),
    .B2(\u_cpu.ALU.u_wallace._1465_ ),
    .Y(\u_cpu.ALU.u_wallace._1959_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7630_  (.A(\u_cpu.ALU.u_wallace._1026_ ),
    .B(\u_cpu.ALU.u_wallace._1486_ ),
    .C(\u_cpu.ALU.u_wallace._0808_ ),
    .D(\u_cpu.ALU.SrcA[19] ),
    .X(\u_cpu.ALU.u_wallace._1960_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7631_  (.A1(\u_cpu.ALU.u_wallace._4470_ ),
    .A2(\u_cpu.ALU.u_wallace._0442_ ),
    .B1(\u_cpu.ALU.u_wallace._1959_ ),
    .B2(\u_cpu.ALU.u_wallace._1960_ ),
    .Y(\u_cpu.ALU.u_wallace._1961_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7632_  (.A1(\u_cpu.ALU.u_wallace._2538_ ),
    .A2(\u_cpu.ALU.u_wallace._0808_ ),
    .B1(\u_cpu.ALU.u_wallace._1100_ ),
    .B2(\u_cpu.ALU.u_wallace._2144_ ),
    .X(\u_cpu.ALU.u_wallace._1962_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7633_  (.A(\u_cpu.ALU.u_wallace._4467_ ),
    .B(\u_cpu.ALU.u_wallace._1497_ ),
    .C(\u_cpu.ALU.u_wallace._1084_ ),
    .D(\u_cpu.ALU.u_wallace._1100_ ),
    .Y(\u_cpu.ALU.u_wallace._1963_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7634_  (.A(\u_cpu.ALU.u_wallace._1962_ ),
    .B(\u_cpu.ALU.u_wallace._1963_ ),
    .C(\u_cpu.ALU.u_wallace._3404_ ),
    .D(\u_cpu.ALU.u_wallace._0850_ ),
    .Y(\u_cpu.ALU.u_wallace._1964_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7635_  (.A1(\u_cpu.ALU.u_wallace._1724_ ),
    .A2(\u_cpu.ALU.u_wallace._1726_ ),
    .B1(\u_cpu.ALU.u_wallace._1752_ ),
    .Y(\u_cpu.ALU.u_wallace._1965_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7636_  (.A1(\u_cpu.ALU.u_wallace._1961_ ),
    .A2(\u_cpu.ALU.u_wallace._1964_ ),
    .B1(\u_cpu.ALU.u_wallace._1965_ ),
    .X(\u_cpu.ALU.u_wallace._1966_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7637_  (.A(\u_cpu.ALU.u_wallace._1530_ ),
    .B(\u_cpu.ALU.u_wallace._1552_ ),
    .C(\u_cpu.ALU.u_wallace._0642_ ),
    .D(\u_cpu.ALU.u_wallace._0802_ ),
    .X(\u_cpu.ALU.u_wallace._1967_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7638_  (.A1(\u_cpu.ALU.u_wallace._1768_ ),
    .A2(\u_cpu.ALU.u_wallace._0826_ ),
    .A3(\u_cpu.ALU.u_wallace._3481_ ),
    .B1(\u_cpu.ALU.u_wallace._1967_ ),
    .X(\u_cpu.ALU.u_wallace._1969_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7639_  (.A(\u_cpu.ALU.u_wallace._1966_ ),
    .B(\u_cpu.ALU.u_wallace._1969_ ),
    .Y(\u_cpu.ALU.u_wallace._1970_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7640_  (.A(\u_cpu.ALU.u_wallace._1724_ ),
    .B(\u_cpu.ALU.u_wallace._1726_ ),
    .Y(\u_cpu.ALU.u_wallace._1971_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7641_  (.A1(\u_cpu.ALU.u_wallace._1728_ ),
    .A2(\u_cpu.ALU.u_wallace._1971_ ),
    .B1(\u_cpu.ALU.u_wallace._1961_ ),
    .C1(\u_cpu.ALU.u_wallace._1964_ ),
    .X(\u_cpu.ALU.u_wallace._1972_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7642_  (.A1(\u_cpu.ALU.u_wallace._1961_ ),
    .A2(\u_cpu.ALU.u_wallace._1964_ ),
    .B1(\u_cpu.ALU.u_wallace._1965_ ),
    .Y(\u_cpu.ALU.u_wallace._1973_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7643_  (.A(\u_cpu.ALU.u_wallace._0325_ ),
    .X(\u_cpu.ALU.u_wallace._1974_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._7644_  (.A1(\u_cpu.ALU.u_wallace._1768_ ),
    .A2(\u_cpu.ALU.u_wallace._1974_ ),
    .A3(\u_cpu.ALU.u_wallace._4542_ ),
    .B1(\u_cpu.ALU.u_wallace._1967_ ),
    .Y(\u_cpu.ALU.u_wallace._1975_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7645_  (.A1(\u_cpu.ALU.u_wallace._1973_ ),
    .A2(\u_cpu.ALU.u_wallace._1972_ ),
    .B1(\u_cpu.ALU.u_wallace._1975_ ),
    .Y(\u_cpu.ALU.u_wallace._1976_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7646_  (.A1(\u_cpu.ALU.u_wallace._1736_ ),
    .A2(\u_cpu.ALU.u_wallace._1735_ ),
    .B1(\u_cpu.ALU.u_wallace._1740_ ),
    .Y(\u_cpu.ALU.u_wallace._1977_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7647_  (.A1(\u_cpu.ALU.u_wallace._1726_ ),
    .A2(\u_cpu.ALU.u_wallace._1725_ ),
    .B1(\u_cpu.ALU.u_wallace._1729_ ),
    .Y(\u_cpu.ALU.u_wallace._1978_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7648_  (.A1(\u_cpu.ALU.u_wallace._1977_ ),
    .A2(\u_cpu.ALU.u_wallace._1746_ ),
    .B1(\u_cpu.ALU.u_wallace._1978_ ),
    .Y(\u_cpu.ALU.u_wallace._1980_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7649_  (.A1(\u_cpu.ALU.u_wallace._1837_ ),
    .A2(\u_cpu.ALU.u_wallace._0626_ ),
    .B1(\u_cpu.ALU.u_wallace._0630_ ),
    .B2(\u_cpu.ALU.u_wallace._2768_ ),
    .Y(\u_cpu.ALU.u_wallace._1981_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7650_  (.A(\u_cpu.ALU.u_wallace._0064_ ),
    .B(\u_cpu.ALU.SrcA[23] ),
    .Y(\u_cpu.ALU.u_wallace._1982_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._7651_  (.A1(\u_cpu.ALU.u_wallace._4431_ ),
    .A2(\u_cpu.ALU.u_wallace._1793_ ),
    .A3(\u_cpu.ALU.u_wallace._1102_ ),
    .A4(\u_cpu.ALU.u_wallace._1073_ ),
    .B1(\u_cpu.ALU.u_wallace._1982_ ),
    .X(\u_cpu.ALU.u_wallace._1983_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7652_  (.A(\u_cpu.ALU.u_wallace._0075_ ),
    .B(\u_cpu.ALU.u_wallace._1734_ ),
    .Y(\u_cpu.ALU.u_wallace._1984_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7653_  (.A1(\u_cpu.ALU.u_wallace._1984_ ),
    .A2(\u_cpu.ALU.u_wallace._1736_ ),
    .B1(\u_cpu.ALU.u_wallace._1733_ ),
    .Y(\u_cpu.ALU.u_wallace._1985_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7654_  (.A1(\u_cpu.ALU.u_wallace._1981_ ),
    .A2(\u_cpu.ALU.u_wallace._1983_ ),
    .B1(\u_cpu.ALU.u_wallace._1985_ ),
    .Y(\u_cpu.ALU.u_wallace._1986_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7655_  (.A(\u_cpu.ALU.SrcA[23] ),
    .Y(\u_cpu.ALU.u_wallace._1987_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7656_  (.A(\u_cpu.ALU.u_wallace._4649_ ),
    .B(\u_cpu.ALU.u_wallace._1782_ ),
    .C(\u_cpu.ALU.u_wallace._0626_ ),
    .D(\u_cpu.ALU.SrcA[17] ),
    .X(\u_cpu.ALU.u_wallace._1988_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._7657_  (.A1(\u_cpu.ALU.u_wallace._4923_ ),
    .A2(\u_cpu.ALU.u_wallace._1987_ ),
    .B1(\u_cpu.ALU.u_wallace._1981_ ),
    .B2(\u_cpu.ALU.u_wallace._1988_ ),
    .X(\u_cpu.ALU.u_wallace._1989_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7658_  (.A(\u_cpu.ALU.u_wallace._0479_ ),
    .B(\u_cpu.ALU.u_wallace._1914_ ),
    .C(\u_cpu.ALU.u_wallace._1730_ ),
    .D(\u_cpu.ALU.SrcA[22] ),
    .X(\u_cpu.ALU.u_wallace._1991_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7659_  (.A1(\u_cpu.ALU.u_wallace._4658_ ),
    .A2(\u_cpu.ALU.u_wallace._1730_ ),
    .B1(\u_cpu.ALU.u_wallace._1734_ ),
    .B2(\u_cpu.ALU.u_wallace._4657_ ),
    .Y(\u_cpu.ALU.u_wallace._1992_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7660_  (.A1(\u_cpu.ALU.u_wallace._1892_ ),
    .A2(\u_cpu.ALU.u_wallace._1271_ ),
    .B1(\u_cpu.ALU.u_wallace._1991_ ),
    .B2(\u_cpu.ALU.u_wallace._1992_ ),
    .Y(\u_cpu.ALU.u_wallace._1993_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7661_  (.A1(\u_cpu.ALU.u_wallace._4658_ ),
    .A2(\u_cpu.ALU.u_wallace._1730_ ),
    .B1(\u_cpu.ALU.u_wallace._1734_ ),
    .B2(\u_cpu.ALU.u_wallace._0206_ ),
    .X(\u_cpu.ALU.u_wallace._1994_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7662_  (.A(\u_cpu.ALU.u_wallace._1957_ ),
    .B(\u_cpu.ALU.u_wallace._1968_ ),
    .C(\u_cpu.ALU.u_wallace._1730_ ),
    .D(\u_cpu.ALU.u_wallace._1734_ ),
    .Y(\u_cpu.ALU.u_wallace._1995_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7663_  (.A(\u_cpu.ALU.u_wallace._1994_ ),
    .B(\u_cpu.ALU.u_wallace._1275_ ),
    .C(\u_cpu.ALU.u_wallace._4662_ ),
    .D(\u_cpu.ALU.u_wallace._1995_ ),
    .Y(\u_cpu.ALU.u_wallace._1996_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7664_  (.A1(\u_cpu.ALU.u_wallace._0634_ ),
    .A2(\u_cpu.ALU.u_wallace._1987_ ),
    .B1(\u_cpu.ALU.u_wallace._1981_ ),
    .B2(\u_cpu.ALU.u_wallace._1988_ ),
    .Y(\u_cpu.ALU.u_wallace._1997_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7665_  (.A1(\u_cpu.ALU.u_wallace._1837_ ),
    .A2(\u_cpu.ALU.u_wallace._0813_ ),
    .B1(\u_cpu.ALU.u_wallace._0630_ ),
    .B2(\u_cpu.ALU.u_wallace._3678_ ),
    .X(\u_cpu.ALU.u_wallace._1998_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7666_  (.A(\u_cpu.ALU.u_wallace._4645_ ),
    .B(\u_cpu.ALU.u_wallace._2834_ ),
    .C(\u_cpu.ALU.u_wallace._0639_ ),
    .D(\u_cpu.ALU.u_wallace._1073_ ),
    .Y(\u_cpu.ALU.u_wallace._1999_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7667_  (.A(\u_cpu.ALU.SrcA[23] ),
    .X(\u_cpu.ALU.u_wallace._2000_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7668_  (.A(\u_cpu.ALU.u_wallace._2000_ ),
    .X(\u_cpu.ALU.u_wallace._2002_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7669_  (.A(\u_cpu.ALU.u_wallace._1998_ ),
    .B(\u_cpu.ALU.u_wallace._1999_ ),
    .C(\u_cpu.ALU.u_wallace._0873_ ),
    .D(\u_cpu.ALU.u_wallace._2002_ ),
    .Y(\u_cpu.ALU.u_wallace._2003_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7670_  (.A1(\u_cpu.ALU.u_wallace._1997_ ),
    .A2(\u_cpu.ALU.u_wallace._2003_ ),
    .B1(\u_cpu.ALU.u_wallace._1985_ ),
    .X(\u_cpu.ALU.u_wallace._2004_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._7671_  (.A1(\u_cpu.ALU.u_wallace._1986_ ),
    .A2(\u_cpu.ALU.u_wallace._1989_ ),
    .B1(\u_cpu.ALU.u_wallace._1993_ ),
    .C1(\u_cpu.ALU.u_wallace._1996_ ),
    .D1(\u_cpu.ALU.u_wallace._2004_ ),
    .Y(\u_cpu.ALU.u_wallace._2005_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7672_  (.A(\u_cpu.ALU.u_wallace._1994_ ),
    .B(\u_cpu.ALU.u_wallace._1275_ ),
    .C(\u_cpu.ALU.u_wallace._4662_ ),
    .D(\u_cpu.ALU.u_wallace._1995_ ),
    .X(\u_cpu.ALU.u_wallace._2006_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._7673_  (.A1(\u_cpu.ALU.u_wallace._1892_ ),
    .A2(\u_cpu.ALU.u_wallace._1271_ ),
    .B1(\u_cpu.ALU.u_wallace._1991_ ),
    .B2(\u_cpu.ALU.u_wallace._1992_ ),
    .X(\u_cpu.ALU.u_wallace._2007_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7674_  (.A1(\u_cpu.ALU.u_wallace._1983_ ),
    .A2(\u_cpu.ALU.u_wallace._1981_ ),
    .B1(\u_cpu.ALU.u_wallace._1985_ ),
    .C1(\u_cpu.ALU.u_wallace._1997_ ),
    .X(\u_cpu.ALU.u_wallace._2008_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7675_  (.A1(\u_cpu.ALU.u_wallace._1997_ ),
    .A2(\u_cpu.ALU.u_wallace._2003_ ),
    .B1(\u_cpu.ALU.u_wallace._1985_ ),
    .Y(\u_cpu.ALU.u_wallace._2009_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7676_  (.A1(\u_cpu.ALU.u_wallace._2006_ ),
    .A2(\u_cpu.ALU.u_wallace._2007_ ),
    .B1(\u_cpu.ALU.u_wallace._2008_ ),
    .B2(\u_cpu.ALU.u_wallace._2009_ ),
    .Y(\u_cpu.ALU.u_wallace._2010_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7677_  (.A1(\u_cpu.ALU.u_wallace._1754_ ),
    .A2(\u_cpu.ALU.u_wallace._1980_ ),
    .B1(\u_cpu.ALU.u_wallace._2005_ ),
    .C1(\u_cpu.ALU.u_wallace._2010_ ),
    .Y(\u_cpu.ALU.u_wallace._2011_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7678_  (.A1(\u_cpu.ALU.u_wallace._1970_ ),
    .A2(\u_cpu.ALU.u_wallace._1972_ ),
    .B1(\u_cpu.ALU.u_wallace._1976_ ),
    .C1(\u_cpu.ALU.u_wallace._2011_ ),
    .Y(\u_cpu.ALU.u_wallace._2013_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._7679_  (.A1(\u_cpu.ALU.u_wallace._1740_ ),
    .A2(\u_cpu.ALU.u_wallace._1755_ ),
    .A3(\u_cpu.ALU.u_wallace._1756_ ),
    .B1(\u_cpu.ALU.u_wallace._1747_ ),
    .B2(\u_cpu.ALU.u_wallace._1761_ ),
    .X(\u_cpu.ALU.u_wallace._2014_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7680_  (.A1(\u_cpu.ALU.u_wallace._2005_ ),
    .A2(\u_cpu.ALU.u_wallace._2010_ ),
    .B1(\u_cpu.ALU.u_wallace._2014_ ),
    .Y(\u_cpu.ALU.u_wallace._2015_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7681_  (.A(\u_cpu.ALU.u_wallace._1748_ ),
    .Y(\u_cpu.ALU.u_wallace._2016_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7682_  (.A(\u_cpu.ALU.u_wallace._1723_ ),
    .B(\u_cpu.ALU.u_wallace._1758_ ),
    .Y(\u_cpu.ALU.u_wallace._2017_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7683_  (.A1(\u_cpu.ALU.u_wallace._2016_ ),
    .A2(\u_cpu.ALU.u_wallace._2017_ ),
    .B1(\u_cpu.ALU.u_wallace._1781_ ),
    .B2(\u_cpu.ALU.u_wallace._1803_ ),
    .Y(\u_cpu.ALU.u_wallace._2018_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7684_  (.A1(\u_cpu.ALU.u_wallace._1728_ ),
    .A2(\u_cpu.ALU.u_wallace._1971_ ),
    .B1(\u_cpu.ALU.u_wallace._1961_ ),
    .C1(\u_cpu.ALU.u_wallace._1964_ ),
    .Y(\u_cpu.ALU.u_wallace._2019_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7685_  (.A1(\u_cpu.ALU.u_wallace._1966_ ),
    .A2(\u_cpu.ALU.u_wallace._2019_ ),
    .B1(\u_cpu.ALU.u_wallace._1969_ ),
    .Y(\u_cpu.ALU.u_wallace._2020_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7686_  (.A(\u_cpu.ALU.u_wallace._1966_ ),
    .B(\u_cpu.ALU.u_wallace._2019_ ),
    .C(\u_cpu.ALU.u_wallace._1969_ ),
    .X(\u_cpu.ALU.u_wallace._2021_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7687_  (.A1(\u_cpu.ALU.u_wallace._1754_ ),
    .A2(\u_cpu.ALU.u_wallace._1980_ ),
    .B1(\u_cpu.ALU.u_wallace._2005_ ),
    .C1(\u_cpu.ALU.u_wallace._2010_ ),
    .X(\u_cpu.ALU.u_wallace._2022_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7688_  (.A1(\u_cpu.ALU.u_wallace._2020_ ),
    .A2(\u_cpu.ALU.u_wallace._2021_ ),
    .B1(\u_cpu.ALU.u_wallace._2022_ ),
    .B2(\u_cpu.ALU.u_wallace._2015_ ),
    .Y(\u_cpu.ALU.u_wallace._2024_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7689_  (.A1(\u_cpu.ALU.u_wallace._2013_ ),
    .A2(\u_cpu.ALU.u_wallace._2015_ ),
    .B1(\u_cpu.ALU.u_wallace._2018_ ),
    .C1(\u_cpu.ALU.u_wallace._2024_ ),
    .Y(\u_cpu.ALU.u_wallace._2025_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7690_  (.A(\u_cpu.ALU.u_wallace._1996_ ),
    .B(\u_cpu.ALU.u_wallace._1993_ ),
    .Y(\u_cpu.ALU.u_wallace._2026_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._7691_  (.A1(\u_cpu.ALU.u_wallace._2008_ ),
    .A2(\u_cpu.ALU.u_wallace._2009_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2026_ ),
    .Y(\u_cpu.ALU.u_wallace._2027_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._7692_  (.A1(\u_cpu.ALU.u_wallace._2006_ ),
    .A2(\u_cpu.ALU.u_wallace._2007_ ),
    .B1(\u_cpu.ALU.u_wallace._1989_ ),
    .B2(\u_cpu.ALU.u_wallace._1986_ ),
    .C1(\u_cpu.ALU.u_wallace._2004_ ),
    .Y(\u_cpu.ALU.u_wallace._2028_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.ALU.u_wallace._7693_  (.A1(\u_cpu.ALU.u_wallace._1744_ ),
    .A2(\u_cpu.ALU.u_wallace._1745_ ),
    .A3(\u_cpu.ALU.u_wallace._1746_ ),
    .B1(\u_cpu.ALU.u_wallace._1978_ ),
    .B2(\u_cpu.ALU.u_wallace._1757_ ),
    .X(\u_cpu.ALU.u_wallace._2029_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7694_  (.A(\u_cpu.ALU.u_wallace._2027_ ),
    .B(\u_cpu.ALU.u_wallace._2028_ ),
    .C(\u_cpu.ALU.u_wallace._2029_ ),
    .Y(\u_cpu.ALU.u_wallace._2030_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7695_  (.A(\u_cpu.ALU.u_wallace._1966_ ),
    .B(\u_cpu.ALU.u_wallace._2019_ ),
    .C(\u_cpu.ALU.u_wallace._1969_ ),
    .Y(\u_cpu.ALU.u_wallace._2031_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7696_  (.A(\u_cpu.ALU.u_wallace._1976_ ),
    .B(\u_cpu.ALU.u_wallace._2031_ ),
    .Y(\u_cpu.ALU.u_wallace._2032_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7697_  (.A1(\u_cpu.ALU.u_wallace._2011_ ),
    .A2(\u_cpu.ALU.u_wallace._2030_ ),
    .B1(\u_cpu.ALU.u_wallace._2032_ ),
    .X(\u_cpu.ALU.u_wallace._2033_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7698_  (.A1(\u_cpu.ALU.u_wallace._2020_ ),
    .A2(\u_cpu.ALU.u_wallace._2021_ ),
    .B1(\u_cpu.ALU.u_wallace._2011_ ),
    .C1(\u_cpu.ALU.u_wallace._2030_ ),
    .Y(\u_cpu.ALU.u_wallace._2035_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7699_  (.A1(\u_cpu.ALU.u_wallace._1784_ ),
    .A2(\u_cpu.ALU.u_wallace._1942_ ),
    .B1(\u_cpu.ALU.u_wallace._1785_ ),
    .Y(\u_cpu.ALU.u_wallace._2036_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7700_  (.A1(\u_cpu.ALU.u_wallace._2036_ ),
    .A2(\u_cpu.ALU.u_wallace._1766_ ),
    .B1(\u_cpu.ALU.u_wallace._1802_ ),
    .Y(\u_cpu.ALU.u_wallace._2037_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7701_  (.A(\u_cpu.ALU.u_wallace._2033_ ),
    .B(\u_cpu.ALU.u_wallace._2035_ ),
    .C(\u_cpu.ALU.u_wallace._2037_ ),
    .Y(\u_cpu.ALU.u_wallace._2038_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._7702_  (.A1_N(\u_cpu.ALU.u_wallace._1956_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1958_ ),
    .B1(\u_cpu.ALU.u_wallace._2025_ ),
    .B2(\u_cpu.ALU.u_wallace._2038_ ),
    .Y(\u_cpu.ALU.u_wallace._2039_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7703_  (.A1(\u_cpu.ALU.u_wallace._1776_ ),
    .A2(\u_cpu.ALU.u_wallace._1777_ ),
    .B1(\u_cpu.ALU.u_wallace._1775_ ),
    .Y(\u_cpu.ALU.u_wallace._2040_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7704_  (.A1(\u_cpu.ALU.u_wallace._1929_ ),
    .A2(\u_cpu.ALU.u_wallace._1939_ ),
    .B1(\u_cpu.ALU.u_wallace._1949_ ),
    .Y(\u_cpu.ALU.u_wallace._2041_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._7705_  (.A1(\u_cpu.ALU.u_wallace._1695_ ),
    .A2(\u_cpu.ALU.u_wallace._1696_ ),
    .B1(\u_cpu.ALU.u_wallace._1708_ ),
    .X(\u_cpu.ALU.u_wallace._2042_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7706_  (.A1_N(\u_cpu.ALU.u_wallace._2040_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2041_ ),
    .B1(\u_cpu.ALU.u_wallace._1710_ ),
    .B2(\u_cpu.ALU.u_wallace._2042_ ),
    .Y(\u_cpu.ALU.u_wallace._2043_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7707_  (.A1(\u_cpu.ALU.u_wallace._1951_ ),
    .A2(\u_cpu.ALU.u_wallace._1955_ ),
    .B1(\u_cpu.ALU.u_wallace._1922_ ),
    .Y(\u_cpu.ALU.u_wallace._2044_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._7708_  (.A1(\u_cpu.ALU.u_wallace._1951_ ),
    .A2(\u_cpu.ALU.u_wallace._2043_ ),
    .B1(\u_cpu.ALU.u_wallace._2044_ ),
    .C1(\u_cpu.ALU.u_wallace._2025_ ),
    .D1(\u_cpu.ALU.u_wallace._2038_ ),
    .X(\u_cpu.ALU.u_wallace._2046_ ));
 sky130_fd_sc_hd__a32oi_2 \u_cpu.ALU.u_wallace._7709_  (.A1(\u_cpu.ALU.u_wallace._1798_ ),
    .A2(\u_cpu.ALU.u_wallace._1799_ ),
    .A3(\u_cpu.ALU.u_wallace._1805_ ),
    .B1(\u_cpu.ALU.u_wallace._1789_ ),
    .B2(\u_cpu.ALU.u_wallace._1809_ ),
    .Y(\u_cpu.ALU.u_wallace._2047_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._7710_  (.A1(\u_cpu.ALU.u_wallace._2039_ ),
    .A2(\u_cpu.ALU.u_wallace._2046_ ),
    .B1(\u_cpu.ALU.u_wallace._2047_ ),
    .X(\u_cpu.ALU.u_wallace._2048_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7711_  (.A1(\u_cpu.ALU.u_wallace._1979_ ),
    .A2(\u_cpu.ALU.u_wallace._1387_ ),
    .B1(\u_cpu.ALU.u_wallace._1210_ ),
    .B2(\u_cpu.ALU.u_wallace._1267_ ),
    .X(\u_cpu.ALU.u_wallace._2049_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7712_  (.A(\u_cpu.ALU.u_wallace._0957_ ),
    .X(\u_cpu.ALU.u_wallace._2050_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7713_  (.A(\u_cpu.ALU.u_wallace._1322_ ),
    .B(\u_cpu.ALU.u_wallace._0906_ ),
    .C(\u_cpu.ALU.u_wallace._2050_ ),
    .D(\u_cpu.ALU.u_wallace._1208_ ),
    .Y(\u_cpu.ALU.u_wallace._2051_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7714_  (.A(\u_cpu.ALU.u_wallace._2049_ ),
    .B(\u_cpu.ALU.u_wallace._2051_ ),
    .C(\u_cpu.ALU.u_wallace._4541_ ),
    .D(\u_cpu.ALU.u_wallace._1392_ ),
    .Y(\u_cpu.ALU.u_wallace._2052_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7715_  (.A(\u_cpu.ALU.u_wallace._1813_ ),
    .X(\u_cpu.ALU.u_wallace._2053_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7716_  (.A1(\u_cpu.ALU.u_wallace._1322_ ),
    .A2(\u_cpu.ALU.u_wallace._2050_ ),
    .B1(\u_cpu.ALU.u_wallace._1208_ ),
    .B2(\u_cpu.ALU.u_wallace._0906_ ),
    .Y(\u_cpu.ALU.u_wallace._2054_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7717_  (.A(\u_cpu.ALU.u_wallace._1979_ ),
    .B(\u_cpu.ALU.u_wallace._2922_ ),
    .C(\u_cpu.ALU.u_wallace._0957_ ),
    .D(\u_cpu.ALU.SrcB[19] ),
    .X(\u_cpu.ALU.u_wallace._2055_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7718_  (.A1(\u_cpu.ALU.u_wallace._0610_ ),
    .A2(\u_cpu.ALU.u_wallace._2053_ ),
    .B1(\u_cpu.ALU.u_wallace._2054_ ),
    .B2(\u_cpu.ALU.u_wallace._2055_ ),
    .Y(\u_cpu.ALU.u_wallace._2057_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.ALU.u_wallace._7719_  (.A1(\u_cpu.ALU.u_wallace._0414_ ),
    .A2(\u_cpu.ALU.u_wallace._2053_ ),
    .A3(\u_cpu.ALU.u_wallace._1814_ ),
    .B1(\u_cpu.ALU.u_wallace._1818_ ),
    .Y(\u_cpu.ALU.u_wallace._2058_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7720_  (.A1(\u_cpu.ALU.u_wallace._2052_ ),
    .A2(\u_cpu.ALU.u_wallace._2057_ ),
    .B1(\u_cpu.ALU.u_wallace._2058_ ),
    .X(\u_cpu.ALU.u_wallace._2059_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7721_  (.A(\u_cpu.ALU.u_wallace._2058_ ),
    .B(\u_cpu.ALU.u_wallace._2052_ ),
    .C(\u_cpu.ALU.u_wallace._2057_ ),
    .Y(\u_cpu.ALU.u_wallace._2060_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7722_  (.A(\u_cpu.ALU.u_wallace._4545_ ),
    .B(\u_cpu.ALU.u_wallace._4463_ ),
    .C(\u_cpu.ALU.u_wallace._1610_ ),
    .D(\u_cpu.ALU.u_wallace._1824_ ),
    .Y(\u_cpu.ALU.u_wallace._2061_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7723_  (.A1(\u_cpu.ALU.u_wallace._4545_ ),
    .A2(\u_cpu.ALU.SrcB[21] ),
    .B1(\u_cpu.ALU.SrcB[22] ),
    .B2(\u_cpu.ALU.u_wallace._0261_ ),
    .X(\u_cpu.ALU.u_wallace._2062_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._7724_  (.A(\u_cpu.ALU.u_wallace._2061_ ),
    .B(\u_cpu.ALU.u_wallace._2062_ ),
    .X(\u_cpu.ALU.u_wallace._2063_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7725_  (.A1(\u_cpu.ALU.u_wallace._2059_ ),
    .A2(\u_cpu.ALU.u_wallace._2060_ ),
    .B1(\u_cpu.ALU.u_wallace._2063_ ),
    .Y(\u_cpu.ALU.u_wallace._2064_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7726_  (.A(\u_cpu.ALU.u_wallace._2059_ ),
    .B(\u_cpu.ALU.u_wallace._2060_ ),
    .C(\u_cpu.ALU.u_wallace._2063_ ),
    .X(\u_cpu.ALU.u_wallace._2065_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7727_  (.A1(\u_cpu.ALU.u_wallace._4444_ ),
    .A2(\u_cpu.ALU.u_wallace._0727_ ),
    .B1(\u_cpu.ALU.u_wallace._0278_ ),
    .B2(\u_cpu.ALU.u_wallace._3689_ ),
    .X(\u_cpu.ALU.u_wallace._2066_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7728_  (.A(\u_cpu.ALU.u_wallace._3623_ ),
    .B(\u_cpu.ALU.u_wallace._4412_ ),
    .C(\u_cpu.ALU.u_wallace._0730_ ),
    .D(\u_cpu.ALU.u_wallace._0732_ ),
    .Y(\u_cpu.ALU.u_wallace._2068_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7729_  (.A(\u_cpu.ALU.u_wallace._2066_ ),
    .B(\u_cpu.ALU.u_wallace._0550_ ),
    .C(\u_cpu.ALU.u_wallace._2801_ ),
    .D(\u_cpu.ALU.u_wallace._2068_ ),
    .Y(\u_cpu.ALU.u_wallace._2069_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7730_  (.A1_N(\u_cpu.ALU.u_wallace._2068_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2066_ ),
    .B1(\u_cpu.ALU.u_wallace._0203_ ),
    .B2(\u_cpu.ALU.u_wallace._0941_ ),
    .Y(\u_cpu.ALU.u_wallace._2070_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7731_  (.A(\u_cpu.ALU.u_wallace._4553_ ),
    .B(\u_cpu.ALU.u_wallace._4650_ ),
    .C(\u_cpu.ALU.u_wallace._4836_ ),
    .D(\u_cpu.ALU.u_wallace._4841_ ),
    .X(\u_cpu.ALU.u_wallace._2071_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7732_  (.A1(\u_cpu.ALU.u_wallace._1691_ ),
    .A2(\u_cpu.ALU.u_wallace._0363_ ),
    .A3(\u_cpu.ALU.u_wallace._4783_ ),
    .B1(\u_cpu.ALU.u_wallace._2071_ ),
    .X(\u_cpu.ALU.u_wallace._2072_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7733_  (.A1(\u_cpu.ALU.u_wallace._2069_ ),
    .A2(\u_cpu.ALU.u_wallace._2070_ ),
    .B1(\u_cpu.ALU.u_wallace._2072_ ),
    .Y(\u_cpu.ALU.u_wallace._2073_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7734_  (.A1(\u_cpu.ALU.u_wallace._4794_ ),
    .A2(\u_cpu.ALU.u_wallace._0028_ ),
    .B1(\u_cpu.ALU.u_wallace._4838_ ),
    .B2(\u_cpu.ALU.u_wallace._4551_ ),
    .Y(\u_cpu.ALU.u_wallace._2074_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7735_  (.A(\u_cpu.ALU.u_wallace._1693_ ),
    .B(\u_cpu.ALU.u_wallace._2074_ ),
    .Y(\u_cpu.ALU.u_wallace._2075_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7736_  (.A1(\u_cpu.ALU.u_wallace._2071_ ),
    .A2(\u_cpu.ALU.u_wallace._2075_ ),
    .B1(\u_cpu.ALU.u_wallace._2070_ ),
    .C1(\u_cpu.ALU.u_wallace._2069_ ),
    .X(\u_cpu.ALU.u_wallace._2076_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7737_  (.A1(\u_cpu.ALU.u_wallace._1834_ ),
    .A2(\u_cpu.ALU.u_wallace._0735_ ),
    .A3(\u_cpu.ALU.u_wallace._4452_ ),
    .B1(\u_cpu.ALU.u_wallace._1832_ ),
    .X(\u_cpu.ALU.u_wallace._2077_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._7738_  (.A1(\u_cpu.ALU.u_wallace._2073_ ),
    .A2(\u_cpu.ALU.u_wallace._2076_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2077_ ),
    .Y(\u_cpu.ALU.u_wallace._2079_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7739_  (.A1(\u_cpu.ALU.u_wallace._2069_ ),
    .A2(\u_cpu.ALU.u_wallace._2070_ ),
    .B1(\u_cpu.ALU.u_wallace._2072_ ),
    .X(\u_cpu.ALU.u_wallace._2080_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7740_  (.A1(\u_cpu.ALU.u_wallace._2071_ ),
    .A2(\u_cpu.ALU.u_wallace._2075_ ),
    .B1(\u_cpu.ALU.u_wallace._2070_ ),
    .C1(\u_cpu.ALU.u_wallace._2069_ ),
    .Y(\u_cpu.ALU.u_wallace._2081_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7741_  (.A(\u_cpu.ALU.u_wallace._2077_ ),
    .B(\u_cpu.ALU.u_wallace._2080_ ),
    .C(\u_cpu.ALU.u_wallace._2081_ ),
    .Y(\u_cpu.ALU.u_wallace._2082_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7742_  (.A1(\u_cpu.ALU.u_wallace._1840_ ),
    .A2(\u_cpu.ALU.u_wallace._1842_ ),
    .B1(\u_cpu.ALU.u_wallace._1844_ ),
    .Y(\u_cpu.ALU.u_wallace._2083_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7743_  (.A1(\u_cpu.ALU.u_wallace._2079_ ),
    .A2(\u_cpu.ALU.u_wallace._2082_ ),
    .B1(\u_cpu.ALU.u_wallace._2083_ ),
    .Y(\u_cpu.ALU.u_wallace._2084_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7744_  (.A(\u_cpu.ALU.u_wallace._1840_ ),
    .B(\u_cpu.ALU.u_wallace._1842_ ),
    .Y(\u_cpu.ALU.u_wallace._2085_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7745_  (.A1(\u_cpu.ALU.u_wallace._1841_ ),
    .A2(\u_cpu.ALU.u_wallace._2085_ ),
    .B1(\u_cpu.ALU.u_wallace._2079_ ),
    .C1(\u_cpu.ALU.u_wallace._2082_ ),
    .X(\u_cpu.ALU.u_wallace._2086_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7746_  (.A1(\u_cpu.ALU.u_wallace._2064_ ),
    .A2(\u_cpu.ALU.u_wallace._2065_ ),
    .B1(\u_cpu.ALU.u_wallace._2084_ ),
    .B2(\u_cpu.ALU.u_wallace._2086_ ),
    .Y(\u_cpu.ALU.u_wallace._2087_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7747_  (.A1(\u_cpu.ALU.u_wallace._2079_ ),
    .A2(\u_cpu.ALU.u_wallace._2082_ ),
    .B1(\u_cpu.ALU.u_wallace._2083_ ),
    .X(\u_cpu.ALU.u_wallace._2088_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7748_  (.A1(\u_cpu.ALU.u_wallace._1841_ ),
    .A2(\u_cpu.ALU.u_wallace._2085_ ),
    .B1(\u_cpu.ALU.u_wallace._2079_ ),
    .C1(\u_cpu.ALU.u_wallace._2082_ ),
    .Y(\u_cpu.ALU.u_wallace._2090_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7749_  (.A(\u_cpu.ALU.u_wallace._2064_ ),
    .B(\u_cpu.ALU.u_wallace._2065_ ),
    .Y(\u_cpu.ALU.u_wallace._2091_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7750_  (.A(\u_cpu.ALU.u_wallace._2088_ ),
    .B(\u_cpu.ALU.u_wallace._2090_ ),
    .C(\u_cpu.ALU.u_wallace._2091_ ),
    .Y(\u_cpu.ALU.u_wallace._2092_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7751_  (.A(\u_cpu.ALU.u_wallace._2087_ ),
    .B(\u_cpu.ALU.u_wallace._2092_ ),
    .Y(\u_cpu.ALU.u_wallace._2093_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7752_  (.A(\u_cpu.ALU.u_wallace._1717_ ),
    .B(\u_cpu.ALU.u_wallace._1718_ ),
    .Y(\u_cpu.ALU.u_wallace._2094_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7753_  (.A1(\u_cpu.ALU.u_wallace._1690_ ),
    .A2(\u_cpu.ALU.u_wallace._2094_ ),
    .B1(\u_cpu.ALU.u_wallace._1807_ ),
    .Y(\u_cpu.ALU.u_wallace._2095_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7754_  (.A(\u_cpu.ALU.u_wallace._1860_ ),
    .Y(\u_cpu.ALU.u_wallace._2096_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7755_  (.A1_N(\u_cpu.ALU.u_wallace._2093_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2095_ ),
    .B1(\u_cpu.ALU.u_wallace._1851_ ),
    .B2(\u_cpu.ALU.u_wallace._2096_ ),
    .Y(\u_cpu.ALU.u_wallace._2097_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7756_  (.A(\u_cpu.ALU.u_wallace._1714_ ),
    .Y(\u_cpu.ALU.u_wallace._2098_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7757_  (.A1(\u_cpu.ALU.u_wallace._2098_ ),
    .A2(\u_cpu.ALU.u_wallace._1807_ ),
    .B1(\u_cpu.ALU.u_wallace._2087_ ),
    .C1(\u_cpu.ALU.u_wallace._2092_ ),
    .X(\u_cpu.ALU.u_wallace._2099_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7758_  (.A1(\u_cpu.ALU.u_wallace._1690_ ),
    .A2(\u_cpu.ALU.u_wallace._2094_ ),
    .B1(\u_cpu.ALU.u_wallace._1807_ ),
    .X(\u_cpu.ALU.u_wallace._2101_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7759_  (.A1(\u_cpu.ALU.u_wallace._2087_ ),
    .A2(\u_cpu.ALU.u_wallace._2092_ ),
    .B1(\u_cpu.ALU.u_wallace._2101_ ),
    .Y(\u_cpu.ALU.u_wallace._2102_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7760_  (.A1(\u_cpu.ALU.u_wallace._1853_ ),
    .A2(\u_cpu.ALU.u_wallace._1858_ ),
    .B1(\u_cpu.ALU.u_wallace._1851_ ),
    .X(\u_cpu.ALU.u_wallace._2103_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._7761_  (.A1(\u_cpu.ALU.u_wallace._2102_ ),
    .A2(\u_cpu.ALU.u_wallace._2099_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2103_ ),
    .Y(\u_cpu.ALU.u_wallace._2104_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7762_  (.A1(\u_cpu.ALU.u_wallace._1951_ ),
    .A2(\u_cpu.ALU.u_wallace._2043_ ),
    .B1(\u_cpu.ALU.u_wallace._2044_ ),
    .C1(\u_cpu.ALU.u_wallace._2025_ ),
    .Y(\u_cpu.ALU.u_wallace._2105_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._7763_  (.A1(\u_cpu.ALU.u_wallace._2029_ ),
    .A2(\u_cpu.ALU.u_wallace._2027_ ),
    .A3(\u_cpu.ALU.u_wallace._2028_ ),
    .B1(\u_cpu.ALU.u_wallace._2032_ ),
    .Y(\u_cpu.ALU.u_wallace._2106_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU.u_wallace._7764_  (.A1(\u_cpu.ALU.u_wallace._2022_ ),
    .A2(\u_cpu.ALU.u_wallace._2015_ ),
    .A3(\u_cpu.ALU.u_wallace._2106_ ),
    .B1(\u_cpu.ALU.u_wallace._2033_ ),
    .C1(\u_cpu.ALU.u_wallace._2037_ ),
    .X(\u_cpu.ALU.u_wallace._2107_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._7765_  (.A1(\u_cpu.ALU.u_wallace._1798_ ),
    .A2(\u_cpu.ALU.u_wallace._1799_ ),
    .A3(\u_cpu.ALU.u_wallace._1805_ ),
    .B1(\u_cpu.ALU.u_wallace._1789_ ),
    .B2(\u_cpu.ALU.u_wallace._1809_ ),
    .X(\u_cpu.ALU.u_wallace._2108_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.ALU.u_wallace._7766_  (.A1_N(\u_cpu.ALU.u_wallace._1956_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1958_ ),
    .B1(\u_cpu.ALU.u_wallace._2025_ ),
    .B2(\u_cpu.ALU.u_wallace._2038_ ),
    .X(\u_cpu.ALU.u_wallace._2109_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7767_  (.A1(\u_cpu.ALU.u_wallace._2105_ ),
    .A2(\u_cpu.ALU.u_wallace._2107_ ),
    .B1(\u_cpu.ALU.u_wallace._2108_ ),
    .C1(\u_cpu.ALU.u_wallace._2109_ ),
    .Y(\u_cpu.ALU.u_wallace._2110_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7768_  (.A1(\u_cpu.ALU.u_wallace._2097_ ),
    .A2(\u_cpu.ALU.u_wallace._2099_ ),
    .B1(\u_cpu.ALU.u_wallace._2104_ ),
    .C1(\u_cpu.ALU.u_wallace._2110_ ),
    .Y(\u_cpu.ALU.u_wallace._2112_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7769_  (.A1(\u_cpu.ALU.u_wallace._2087_ ),
    .A2(\u_cpu.ALU.u_wallace._2092_ ),
    .B1(\u_cpu.ALU.u_wallace._2101_ ),
    .X(\u_cpu.ALU.u_wallace._2113_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7770_  (.A1(\u_cpu.ALU.u_wallace._2098_ ),
    .A2(\u_cpu.ALU.u_wallace._1807_ ),
    .B1(\u_cpu.ALU.u_wallace._2087_ ),
    .C1(\u_cpu.ALU.u_wallace._2092_ ),
    .Y(\u_cpu.ALU.u_wallace._2114_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7771_  (.A1(\u_cpu.ALU.u_wallace._1851_ ),
    .A2(\u_cpu.ALU.u_wallace._2096_ ),
    .B1(\u_cpu.ALU.u_wallace._2113_ ),
    .C1(\u_cpu.ALU.u_wallace._2114_ ),
    .Y(\u_cpu.ALU.u_wallace._2115_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7772_  (.A1(\u_cpu.ALU.u_wallace._2039_ ),
    .A2(\u_cpu.ALU.u_wallace._2046_ ),
    .B1(\u_cpu.ALU.u_wallace._2047_ ),
    .Y(\u_cpu.ALU.u_wallace._2116_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7773_  (.A1(\u_cpu.ALU.u_wallace._2104_ ),
    .A2(\u_cpu.ALU.u_wallace._2115_ ),
    .B1(\u_cpu.ALU.u_wallace._2110_ ),
    .B2(\u_cpu.ALU.u_wallace._2116_ ),
    .X(\u_cpu.ALU.u_wallace._2117_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7774_  (.A1(\u_cpu.ALU.u_wallace._1872_ ),
    .A2(\u_cpu.ALU.u_wallace._1866_ ),
    .A3(\u_cpu.ALU.u_wallace._1876_ ),
    .B1(\u_cpu.ALU.u_wallace._1811_ ),
    .X(\u_cpu.ALU.u_wallace._2118_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7775_  (.A1(\u_cpu.ALU.u_wallace._2048_ ),
    .A2(\u_cpu.ALU.u_wallace._2112_ ),
    .B1(\u_cpu.ALU.u_wallace._2117_ ),
    .C1(\u_cpu.ALU.u_wallace._2118_ ),
    .Y(\u_cpu.ALU.u_wallace._2119_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7776_  (.A1(\u_cpu.ALU.u_wallace._2113_ ),
    .A2(\u_cpu.ALU.u_wallace._2114_ ),
    .B1(\u_cpu.ALU.u_wallace._2103_ ),
    .Y(\u_cpu.ALU.u_wallace._2120_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7777_  (.A1(\u_cpu.ALU.u_wallace._1851_ ),
    .A2(\u_cpu.ALU.u_wallace._2096_ ),
    .B1(\u_cpu.ALU.u_wallace._2113_ ),
    .C1(\u_cpu.ALU.u_wallace._2114_ ),
    .X(\u_cpu.ALU.u_wallace._2121_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._7778_  (.A1_N(\u_cpu.ALU.u_wallace._2120_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2121_ ),
    .B1(\u_cpu.ALU.u_wallace._2110_ ),
    .B2(\u_cpu.ALU.u_wallace._2116_ ),
    .Y(\u_cpu.ALU.u_wallace._2123_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._7779_  (.A1(\u_cpu.ALU.u_wallace._2097_ ),
    .A2(\u_cpu.ALU.u_wallace._2099_ ),
    .B1(\u_cpu.ALU.u_wallace._2104_ ),
    .C1(\u_cpu.ALU.u_wallace._2110_ ),
    .D1(\u_cpu.ALU.u_wallace._2116_ ),
    .X(\u_cpu.ALU.u_wallace._2124_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._7780_  (.A1(\u_cpu.ALU.u_wallace._1872_ ),
    .A2(\u_cpu.ALU.u_wallace._1866_ ),
    .A3(\u_cpu.ALU.u_wallace._1876_ ),
    .B1(\u_cpu.ALU.u_wallace._1811_ ),
    .Y(\u_cpu.ALU.u_wallace._2125_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7781_  (.A1(\u_cpu.ALU.u_wallace._2123_ ),
    .A2(\u_cpu.ALU.u_wallace._2124_ ),
    .B1(\u_cpu.ALU.u_wallace._2125_ ),
    .Y(\u_cpu.ALU.u_wallace._2126_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7782_  (.A(\u_cpu.ALU.u_wallace._1821_ ),
    .B(\u_cpu.ALU.u_wallace._1817_ ),
    .C(\u_cpu.ALU.u_wallace._1819_ ),
    .X(\u_cpu.ALU.u_wallace._2127_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7783_  (.A(\u_cpu.ALU.u_wallace._3996_ ),
    .B(\u_cpu.ALU.u_wallace._0173_ ),
    .C(\u_cpu.ALU.u_wallace._1611_ ),
    .D(\u_cpu.ALU.u_wallace._1855_ ),
    .X(\u_cpu.ALU.u_wallace._2128_ ));
 sky130_fd_sc_hd__or4_2 \u_cpu.ALU.u_wallace._7784_  (.A(\u_cpu.ALU.u_wallace._1856_ ),
    .B(\u_cpu.ALU.u_wallace._2127_ ),
    .C(\u_cpu.ALU.u_wallace._2128_ ),
    .D(\u_cpu.ALU.u_wallace._1827_ ),
    .X(\u_cpu.ALU.u_wallace._2129_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._7785_  (.A(\u_cpu.ALU.u_wallace._1823_ ),
    .B(\u_cpu.ALU.u_wallace._2128_ ),
    .X(\u_cpu.ALU.u_wallace._2130_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7786_  (.A(\u_cpu.ALU.SrcB[23] ),
    .Y(\u_cpu.ALU.u_wallace._2131_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._7787_  (.A1(\u_cpu.ALU.u_wallace._2129_ ),
    .A2(\u_cpu.ALU.u_wallace._2130_ ),
    .B1(\u_cpu.ALU.u_wallace._0043_ ),
    .C1(\u_cpu.ALU.u_wallace._2131_ ),
    .X(\u_cpu.ALU.u_wallace._2132_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7788_  (.A(\u_cpu.ALU.SrcB[23] ),
    .X(\u_cpu.ALU.u_wallace._2134_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7789_  (.A(\u_cpu.ALU.u_wallace._2129_ ),
    .B(\u_cpu.ALU.u_wallace._2130_ ),
    .Y(\u_cpu.ALU.u_wallace._2135_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7790_  (.A1(\u_cpu.ALU.u_wallace._1886_ ),
    .A2(\u_cpu.ALU.u_wallace._2134_ ),
    .B1(\u_cpu.ALU.u_wallace._2135_ ),
    .X(\u_cpu.ALU.u_wallace._2136_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7791_  (.A(\u_cpu.ALU.u_wallace._2132_ ),
    .B(\u_cpu.ALU.u_wallace._2136_ ),
    .Y(\u_cpu.ALU.u_wallace._2137_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7792_  (.A1(\u_cpu.ALU.u_wallace._1861_ ),
    .A2(\u_cpu.ALU.u_wallace._1876_ ),
    .B1(\u_cpu.ALU.u_wallace._2137_ ),
    .Y(\u_cpu.ALU.u_wallace._2138_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7793_  (.A(\u_cpu.ALU.u_wallace._1861_ ),
    .B(\u_cpu.ALU.u_wallace._1876_ ),
    .C(\u_cpu.ALU.u_wallace._2137_ ),
    .X(\u_cpu.ALU.u_wallace._2139_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7794_  (.A1_N(\u_cpu.ALU.u_wallace._2119_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2126_ ),
    .B1(\u_cpu.ALU.u_wallace._2138_ ),
    .B2(\u_cpu.ALU.u_wallace._2139_ ),
    .Y(\u_cpu.ALU.u_wallace._2140_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._7795_  (.A1(\u_cpu.ALU.u_wallace._1862_ ),
    .A2(\u_cpu.ALU.u_wallace._1877_ ),
    .B1(\u_cpu.ALU.u_wallace._2137_ ),
    .X(\u_cpu.ALU.u_wallace._2141_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7796_  (.A1(\u_cpu.ALU.u_wallace._1863_ ),
    .A2(\u_cpu.ALU.u_wallace._1864_ ),
    .B1(\u_cpu.ALU.u_wallace._1862_ ),
    .X(\u_cpu.ALU.u_wallace._2142_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7797_  (.A(\u_cpu.ALU.u_wallace._2142_ ),
    .B(\u_cpu.ALU.u_wallace._2137_ ),
    .Y(\u_cpu.ALU.u_wallace._2143_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU.u_wallace._7798_  (.A1(\u_cpu.ALU.u_wallace._2047_ ),
    .A2(\u_cpu.ALU.u_wallace._2039_ ),
    .A3(\u_cpu.ALU.u_wallace._2046_ ),
    .B1(\u_cpu.ALU.u_wallace._2104_ ),
    .C1(\u_cpu.ALU.u_wallace._2115_ ),
    .X(\u_cpu.ALU.u_wallace._2145_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7799_  (.A1(\u_cpu.ALU.u_wallace._2145_ ),
    .A2(\u_cpu.ALU.u_wallace._2116_ ),
    .B1(\u_cpu.ALU.u_wallace._2123_ ),
    .Y(\u_cpu.ALU.u_wallace._2146_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._7800_  (.A1(\u_cpu.ALU.u_wallace._2141_ ),
    .A2(\u_cpu.ALU.u_wallace._2143_ ),
    .B1(\u_cpu.ALU.u_wallace._2118_ ),
    .B2(\u_cpu.ALU.u_wallace._2146_ ),
    .C1(\u_cpu.ALU.u_wallace._2119_ ),
    .Y(\u_cpu.ALU.u_wallace._2147_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7801_  (.A1(\u_cpu.ALU.u_wallace._1901_ ),
    .A2(\u_cpu.ALU.u_wallace._1921_ ),
    .B1(\u_cpu.ALU.u_wallace._2140_ ),
    .C1(\u_cpu.ALU.u_wallace._2147_ ),
    .X(\u_cpu.ALU.u_wallace._2148_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7802_  (.A1(\u_cpu.ALU.u_wallace._1884_ ),
    .A2(\u_cpu.ALU.u_wallace._1902_ ),
    .B1(\u_cpu.ALU.u_wallace._1904_ ),
    .Y(\u_cpu.ALU.u_wallace._2149_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7803_  (.A1(\u_cpu.ALU.u_wallace._2140_ ),
    .A2(\u_cpu.ALU.u_wallace._2147_ ),
    .B1(\u_cpu.ALU.u_wallace._2149_ ),
    .Y(\u_cpu.ALU.u_wallace._2150_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7804_  (.A1(\u_cpu.ALU.u_wallace._2148_ ),
    .A2(\u_cpu.ALU.u_wallace._2150_ ),
    .B1(\u_cpu.ALU.u_wallace._1891_ ),
    .Y(\u_cpu.ALU.u_wallace._2151_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._7805_  (.A1(\u_cpu.ALU.u_wallace._1655_ ),
    .A2(\u_cpu.ALU.u_wallace._1653_ ),
    .B1(\u_cpu.ALU.u_wallace._1650_ ),
    .X(\u_cpu.ALU.u_wallace._2152_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7806_  (.A1(\u_cpu.ALU.u_wallace._1901_ ),
    .A2(\u_cpu.ALU.u_wallace._1921_ ),
    .B1(\u_cpu.ALU.u_wallace._2140_ ),
    .C1(\u_cpu.ALU.u_wallace._2147_ ),
    .Y(\u_cpu.ALU.u_wallace._2153_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7807_  (.A1(\u_cpu.ALU.u_wallace._2140_ ),
    .A2(\u_cpu.ALU.u_wallace._2147_ ),
    .B1(\u_cpu.ALU.u_wallace._2149_ ),
    .X(\u_cpu.ALU.u_wallace._2154_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7808_  (.A1(\u_cpu.ALU.u_wallace._1889_ ),
    .A2(\u_cpu.ALU.u_wallace._2152_ ),
    .B1(\u_cpu.ALU.u_wallace._2153_ ),
    .C1(\u_cpu.ALU.u_wallace._2154_ ),
    .Y(\u_cpu.ALU.u_wallace._2156_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7809_  (.A1(\u_cpu.ALU.u_wallace._1900_ ),
    .A2(\u_cpu.ALU.u_wallace._1907_ ),
    .B1(\u_cpu.ALU.u_wallace._1912_ ),
    .Y(\u_cpu.ALU.u_wallace._2157_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7810_  (.A(\u_cpu.ALU.u_wallace._2151_ ),
    .B(\u_cpu.ALU.u_wallace._2156_ ),
    .C(\u_cpu.ALU.u_wallace._2157_ ),
    .Y(\u_cpu.ALU.u_wallace._2158_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7811_  (.A1(\u_cpu.ALU.u_wallace._1906_ ),
    .A2(\u_cpu.ALU.u_wallace._1911_ ),
    .B1(\u_cpu.ALU.u_wallace._1905_ ),
    .Y(\u_cpu.ALU.u_wallace._2159_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._7812_  (.A1(\u_cpu.ALU.u_wallace._1654_ ),
    .A2(\u_cpu.ALU.u_wallace._1664_ ),
    .B1(\u_cpu.ALU.u_wallace._1888_ ),
    .C1(\u_cpu.ALU.u_wallace._2153_ ),
    .D1(\u_cpu.ALU.u_wallace._2154_ ),
    .Y(\u_cpu.ALU.u_wallace._2160_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7813_  (.A1(\u_cpu.ALU.u_wallace._1889_ ),
    .A2(\u_cpu.ALU.u_wallace._2152_ ),
    .B1(\u_cpu.ALU.u_wallace._2148_ ),
    .B2(\u_cpu.ALU.u_wallace._2150_ ),
    .Y(\u_cpu.ALU.u_wallace._2161_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7814_  (.A(\u_cpu.ALU.u_wallace._2159_ ),
    .B(\u_cpu.ALU.u_wallace._2160_ ),
    .C(\u_cpu.ALU.u_wallace._2161_ ),
    .Y(\u_cpu.ALU.u_wallace._2162_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7815_  (.A(\u_cpu.ALU.u_wallace._2158_ ),
    .B(\u_cpu.ALU.u_wallace._2162_ ),
    .Y(\u_cpu.ALU.u_wallace._2163_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._7816_  (.A1(\u_cpu.ALU.u_wallace._1674_ ),
    .A2(\u_cpu.ALU.u_wallace._1908_ ),
    .A3(\u_cpu.ALU.u_wallace._1909_ ),
    .B1(\u_cpu.ALU.u_wallace._2163_ ),
    .X(\u_cpu.ALU.u_wallace._2164_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._7817_  (.A1(\u_cpu.ALU.u_wallace._1680_ ),
    .A2(\u_cpu.ALU.u_wallace._1913_ ),
    .A3(\u_cpu.ALU.u_wallace._1915_ ),
    .A4(\u_cpu.ALU.u_wallace._2158_ ),
    .B1(\u_cpu.ALU.u_wallace._2164_ ),
    .X(\u_cpu.ALU.u_wallace._2165_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU.u_wallace._7818_  (.A1(\u_cpu.ALU.u_wallace._1906_ ),
    .A2(\u_cpu.ALU.u_wallace._1911_ ),
    .A3(\u_cpu.ALU.u_wallace._1912_ ),
    .B1(\u_cpu.ALU.u_wallace._1674_ ),
    .C1(\u_cpu.ALU.u_wallace._1689_ ),
    .X(\u_cpu.ALU.u_wallace._2167_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7819_  (.A1(\u_cpu.ALU.u_wallace._1913_ ),
    .A2(\u_cpu.ALU.u_wallace._2167_ ),
    .B1(\u_cpu.ALU.u_wallace._1920_ ),
    .B2(\u_cpu.ALU.u_wallace._1917_ ),
    .X(\u_cpu.ALU.u_wallace._2168_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu.ALU.u_wallace._7820_  (.A(\u_cpu.ALU.u_wallace._2165_ ),
    .B(\u_cpu.ALU.u_wallace._2168_ ),
    .Y(\u_cpu.ALU.Product_Wallace[23] ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7821_  (.A1(\u_cpu.ALU.u_wallace._2141_ ),
    .A2(\u_cpu.ALU.u_wallace._2143_ ),
    .B1(\u_cpu.ALU.u_wallace._2118_ ),
    .B2(\u_cpu.ALU.u_wallace._2146_ ),
    .Y(\u_cpu.ALU.u_wallace._2169_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.ALU.u_wallace._7822_  (.A1(\u_cpu.ALU.u_wallace._1945_ ),
    .A2(\u_cpu.ALU.u_wallace._1947_ ),
    .A3(\u_cpu.ALU.u_wallace._1929_ ),
    .B1(\u_cpu.ALU.u_wallace._1938_ ),
    .Y(\u_cpu.ALU.u_wallace._2170_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7823_  (.A(\u_cpu.ALU.u_wallace._2170_ ),
    .Y(\u_cpu.ALU.u_wallace._2171_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7824_  (.A(\u_cpu.ALU.u_wallace._4609_ ),
    .B(\u_cpu.ALU.u_wallace._0188_ ),
    .Y(\u_cpu.ALU.u_wallace._2172_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7825_  (.A1(\u_cpu.ALU.u_wallace._4848_ ),
    .A2(\u_cpu.ALU.u_wallace._0313_ ),
    .B1(\u_cpu.ALU.u_wallace._0330_ ),
    .B2(\u_cpu.ALU.u_wallace._4720_ ),
    .Y(\u_cpu.ALU.u_wallace._2173_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._7826_  (.A1(\u_cpu.ALU.u_wallace._2172_ ),
    .A2(\u_cpu.ALU.u_wallace._2173_ ),
    .B1(\u_cpu.ALU.u_wallace._1923_ ),
    .X(\u_cpu.ALU.u_wallace._2174_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7827_  (.A(\u_cpu.ALU.u_wallace._4720_ ),
    .B(\u_cpu.ALU.u_wallace._0045_ ),
    .C(\u_cpu.ALU.u_wallace._0330_ ),
    .D(\u_cpu.ALU.u_wallace._0448_ ),
    .Y(\u_cpu.ALU.u_wallace._2175_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7828_  (.A1(\u_cpu.ALU.u_wallace._4291_ ),
    .A2(\u_cpu.ALU.u_wallace._0324_ ),
    .B1(\u_cpu.ALU.u_wallace._0441_ ),
    .B2(\u_cpu.ALU.u_wallace._4007_ ),
    .X(\u_cpu.ALU.u_wallace._2177_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._7829_  (.A1_N(\u_cpu.ALU.u_wallace._4601_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1323_ ),
    .B1(\u_cpu.ALU.u_wallace._2175_ ),
    .B2(\u_cpu.ALU.u_wallace._2177_ ),
    .Y(\u_cpu.ALU.u_wallace._2178_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7830_  (.A1(\u_cpu.ALU.u_wallace._4848_ ),
    .A2(\u_cpu.ALU.u_wallace._0330_ ),
    .B1(\u_cpu.ALU.u_wallace._0850_ ),
    .B2(\u_cpu.ALU.u_wallace._4720_ ),
    .Y(\u_cpu.ALU.u_wallace._2179_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7831_  (.A(\u_cpu.ALU.u_wallace._4609_ ),
    .B(\u_cpu.ALU.u_wallace._0179_ ),
    .Y(\u_cpu.ALU.u_wallace._2180_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7832_  (.A(\u_cpu.ALU.u_wallace._4716_ ),
    .B(\u_cpu.ALU.u_wallace._4598_ ),
    .C(\u_cpu.ALU.u_wallace._0332_ ),
    .D(\u_cpu.ALU.u_wallace._0441_ ),
    .X(\u_cpu.ALU.u_wallace._2181_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._7833_  (.A(\u_cpu.ALU.u_wallace._2179_ ),
    .B(\u_cpu.ALU.u_wallace._2180_ ),
    .C(\u_cpu.ALU.u_wallace._2181_ ),
    .Y(\u_cpu.ALU.u_wallace._2182_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7834_  (.A(\u_cpu.ALU.u_wallace._0028_ ),
    .B(\u_cpu.ALU.u_wallace._4785_ ),
    .C(\u_cpu.ALU.u_wallace._0144_ ),
    .D(\u_cpu.ALU.u_wallace._4921_ ),
    .Y(\u_cpu.ALU.u_wallace._2183_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7835_  (.A1(\u_cpu.ALU.u_wallace._4900_ ),
    .A2(\u_cpu.ALU.u_wallace._4841_ ),
    .B1(\u_cpu.ALU.u_wallace._4907_ ),
    .B2(\u_cpu.ALU.u_wallace._0364_ ),
    .X(\u_cpu.ALU.u_wallace._2184_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7836_  (.A1(\u_cpu.ALU.u_wallace._0169_ ),
    .A2(\u_cpu.ALU.u_wallace._0037_ ),
    .B1(\u_cpu.ALU.u_wallace._2183_ ),
    .C1(\u_cpu.ALU.u_wallace._2184_ ),
    .Y(\u_cpu.ALU.u_wallace._2185_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7837_  (.A(\u_cpu.ALU.u_wallace._4653_ ),
    .B(\u_cpu.ALU.SrcB[13] ),
    .Y(\u_cpu.ALU.u_wallace._2186_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7838_  (.A1(\u_cpu.ALU.u_wallace._2183_ ),
    .A2(\u_cpu.ALU.u_wallace._2184_ ),
    .B1(\u_cpu.ALU.u_wallace._2186_ ),
    .X(\u_cpu.ALU.u_wallace._2188_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7839_  (.A(\u_cpu.ALU.u_wallace._2185_ ),
    .B(\u_cpu.ALU.u_wallace._2188_ ),
    .Y(\u_cpu.ALU.u_wallace._2189_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7840_  (.A1(\u_cpu.ALU.u_wallace._2178_ ),
    .A2(\u_cpu.ALU.u_wallace._2182_ ),
    .B1(\u_cpu.ALU.u_wallace._2174_ ),
    .Y(\u_cpu.ALU.u_wallace._2190_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU.u_wallace._7841_  (.A1(\u_cpu.ALU.u_wallace._2174_ ),
    .A2(\u_cpu.ALU.u_wallace._2178_ ),
    .A3(\u_cpu.ALU.u_wallace._2182_ ),
    .B1(\u_cpu.ALU.u_wallace._2189_ ),
    .C1(\u_cpu.ALU.u_wallace._2190_ ),
    .X(\u_cpu.ALU.u_wallace._2191_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7842_  (.A(\u_cpu.ALU.u_wallace._1973_ ),
    .B(\u_cpu.ALU.u_wallace._1975_ ),
    .Y(\u_cpu.ALU.u_wallace._2192_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7843_  (.A1(\u_cpu.ALU.u_wallace._2172_ ),
    .A2(\u_cpu.ALU.u_wallace._2173_ ),
    .B1(\u_cpu.ALU.u_wallace._1923_ ),
    .Y(\u_cpu.ALU.u_wallace._2193_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7844_  (.A1(\u_cpu.ALU.u_wallace._4604_ ),
    .A2(\u_cpu.ALU.u_wallace._0320_ ),
    .B1(\u_cpu.ALU.u_wallace._2175_ ),
    .B2(\u_cpu.ALU.u_wallace._2177_ ),
    .X(\u_cpu.ALU.u_wallace._2194_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7845_  (.A(\u_cpu.ALU.u_wallace._2177_ ),
    .B(\u_cpu.ALU.u_wallace._0652_ ),
    .C(\u_cpu.ALU.u_wallace._0052_ ),
    .D(\u_cpu.ALU.u_wallace._2175_ ),
    .Y(\u_cpu.ALU.u_wallace._2195_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7846_  (.A(\u_cpu.ALU.u_wallace._2193_ ),
    .B(\u_cpu.ALU.u_wallace._2194_ ),
    .C(\u_cpu.ALU.u_wallace._2195_ ),
    .Y(\u_cpu.ALU.u_wallace._2196_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7847_  (.A(\u_cpu.ALU.u_wallace._0028_ ),
    .B(\u_cpu.ALU.u_wallace._4787_ ),
    .C(\u_cpu.ALU.u_wallace._0144_ ),
    .D(\u_cpu.ALU.u_wallace._4921_ ),
    .X(\u_cpu.ALU.u_wallace._2197_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7848_  (.A1(\u_cpu.ALU.u_wallace._4787_ ),
    .A2(\u_cpu.ALU.u_wallace._0029_ ),
    .B1(\u_cpu.ALU.u_wallace._0188_ ),
    .B2(\u_cpu.ALU.u_wallace._4837_ ),
    .Y(\u_cpu.ALU.u_wallace._2199_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._7849_  (.A1(\u_cpu.ALU.u_wallace._0169_ ),
    .A2(\u_cpu.ALU.u_wallace._0037_ ),
    .B1(\u_cpu.ALU.u_wallace._2197_ ),
    .B2(\u_cpu.ALU.u_wallace._2199_ ),
    .X(\u_cpu.ALU.u_wallace._2200_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7850_  (.A(\u_cpu.ALU.u_wallace._2184_ ),
    .B(\u_cpu.ALU.u_wallace._0057_ ),
    .C(\u_cpu.ALU.u_wallace._1129_ ),
    .D(\u_cpu.ALU.u_wallace._2183_ ),
    .X(\u_cpu.ALU.u_wallace._2201_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7851_  (.A1_N(\u_cpu.ALU.u_wallace._2196_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2190_ ),
    .B1(\u_cpu.ALU.u_wallace._2200_ ),
    .B2(\u_cpu.ALU.u_wallace._2201_ ),
    .Y(\u_cpu.ALU.u_wallace._2202_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7852_  (.A1(\u_cpu.ALU.u_wallace._1972_ ),
    .A2(\u_cpu.ALU.u_wallace._2192_ ),
    .B1(\u_cpu.ALU.u_wallace._2202_ ),
    .Y(\u_cpu.ALU.u_wallace._2203_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7853_  (.A1(\u_cpu.ALU.u_wallace._2196_ ),
    .A2(\u_cpu.ALU.u_wallace._2190_ ),
    .B1(\u_cpu.ALU.u_wallace._2189_ ),
    .Y(\u_cpu.ALU.u_wallace._2204_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7854_  (.A1(\u_cpu.ALU.u_wallace._1966_ ),
    .A2(\u_cpu.ALU.u_wallace._1969_ ),
    .B1(\u_cpu.ALU.u_wallace._1972_ ),
    .Y(\u_cpu.ALU.u_wallace._2205_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7855_  (.A1(\u_cpu.ALU.u_wallace._2191_ ),
    .A2(\u_cpu.ALU.u_wallace._2204_ ),
    .B1(\u_cpu.ALU.u_wallace._2205_ ),
    .Y(\u_cpu.ALU.u_wallace._2206_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7856_  (.A1(\u_cpu.ALU.u_wallace._2191_ ),
    .A2(\u_cpu.ALU.u_wallace._2203_ ),
    .B1(\u_cpu.ALU.u_wallace._2206_ ),
    .Y(\u_cpu.ALU.u_wallace._2207_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._7857_  (.A1(\u_cpu.ALU.u_wallace._2172_ ),
    .A2(\u_cpu.ALU.u_wallace._2173_ ),
    .B1(\u_cpu.ALU.u_wallace._2178_ ),
    .B2(\u_cpu.ALU.u_wallace._2182_ ),
    .C1(\u_cpu.ALU.u_wallace._1923_ ),
    .X(\u_cpu.ALU.u_wallace._2208_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7858_  (.A(\u_cpu.ALU.u_wallace._2196_ ),
    .B(\u_cpu.ALU.u_wallace._2189_ ),
    .Y(\u_cpu.ALU.u_wallace._2210_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7859_  (.A1(\u_cpu.ALU.u_wallace._2208_ ),
    .A2(\u_cpu.ALU.u_wallace._2210_ ),
    .B1(\u_cpu.ALU.u_wallace._2202_ ),
    .Y(\u_cpu.ALU.u_wallace._2211_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7860_  (.A1(\u_cpu.ALU.u_wallace._2019_ ),
    .A2(\u_cpu.ALU.u_wallace._2031_ ),
    .B1(\u_cpu.ALU.u_wallace._2211_ ),
    .Y(\u_cpu.ALU.u_wallace._2212_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7861_  (.A(\u_cpu.ALU.u_wallace._2206_ ),
    .B(\u_cpu.ALU.u_wallace._2170_ ),
    .Y(\u_cpu.ALU.u_wallace._2213_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7862_  (.A1_N(\u_cpu.ALU.u_wallace._2171_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2207_ ),
    .B1(\u_cpu.ALU.u_wallace._2212_ ),
    .B2(\u_cpu.ALU.u_wallace._2213_ ),
    .Y(\u_cpu.ALU.u_wallace._2214_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7863_  (.A(\u_cpu.ALU.SrcA[24] ),
    .Y(\u_cpu.ALU.u_wallace._2215_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7864_  (.A1(\u_cpu.ALU.u_wallace._2878_ ),
    .A2(\u_cpu.ALU.u_wallace._0626_ ),
    .B1(\u_cpu.ALU.u_wallace._0808_ ),
    .B2(\u_cpu.ALU.u_wallace._2768_ ),
    .Y(\u_cpu.ALU.u_wallace._2216_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7865_  (.A(\u_cpu.ALU.u_wallace._4649_ ),
    .B(\u_cpu.ALU.u_wallace._2878_ ),
    .C(\u_cpu.ALU.u_wallace._0626_ ),
    .D(\u_cpu.ALU.u_wallace._0808_ ),
    .X(\u_cpu.ALU.u_wallace._2217_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7866_  (.A1(\u_cpu.ALU.u_wallace._4923_ ),
    .A2(\u_cpu.ALU.u_wallace._2215_ ),
    .B1(\u_cpu.ALU.u_wallace._2216_ ),
    .B2(\u_cpu.ALU.u_wallace._2217_ ),
    .Y(\u_cpu.ALU.u_wallace._2218_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7867_  (.A1(\u_cpu.ALU.u_wallace._2790_ ),
    .A2(\u_cpu.ALU.u_wallace._0813_ ),
    .B1(\u_cpu.ALU.u_wallace._1084_ ),
    .B2(\u_cpu.ALU.u_wallace._2768_ ),
    .X(\u_cpu.ALU.u_wallace._2219_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7868_  (.A(\u_cpu.ALU.u_wallace._3678_ ),
    .B(\u_cpu.ALU.u_wallace._2790_ ),
    .C(\u_cpu.ALU.u_wallace._0813_ ),
    .D(\u_cpu.ALU.u_wallace._1084_ ),
    .Y(\u_cpu.ALU.u_wallace._2221_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7869_  (.A(\u_cpu.ALU.SrcA[24] ),
    .X(\u_cpu.ALU.u_wallace._2222_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7870_  (.A(\u_cpu.ALU.u_wallace._2219_ ),
    .B(\u_cpu.ALU.u_wallace._2221_ ),
    .C(\u_cpu.ALU.u_wallace._0873_ ),
    .D(\u_cpu.ALU.u_wallace._2222_ ),
    .Y(\u_cpu.ALU.u_wallace._2223_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7871_  (.A1(\u_cpu.ALU.u_wallace._1982_ ),
    .A2(\u_cpu.ALU.u_wallace._1981_ ),
    .B1(\u_cpu.ALU.u_wallace._1999_ ),
    .Y(\u_cpu.ALU.u_wallace._2224_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7872_  (.A1(\u_cpu.ALU.u_wallace._2218_ ),
    .A2(\u_cpu.ALU.u_wallace._2223_ ),
    .B1(\u_cpu.ALU.u_wallace._2224_ ),
    .Y(\u_cpu.ALU.u_wallace._2225_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7873_  (.A(\u_cpu.ALU.SrcA[24] ),
    .X(\u_cpu.ALU.u_wallace._2226_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7874_  (.A(\u_cpu.ALU.u_wallace._2747_ ),
    .B(\u_cpu.ALU.u_wallace._2226_ ),
    .Y(\u_cpu.ALU.u_wallace._2227_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._7875_  (.A(\u_cpu.ALU.u_wallace._2227_ ),
    .B(\u_cpu.ALU.u_wallace._2216_ ),
    .C(\u_cpu.ALU.u_wallace._2217_ ),
    .Y(\u_cpu.ALU.u_wallace._2228_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7876_  (.A(\u_cpu.ALU.u_wallace._4431_ ),
    .B(\u_cpu.ALU.u_wallace._0642_ ),
    .Y(\u_cpu.ALU.u_wallace._2229_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7877_  (.A(\u_cpu.ALU.u_wallace._3777_ ),
    .B(\u_cpu.ALU.u_wallace._1102_ ),
    .Y(\u_cpu.ALU.u_wallace._2230_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7878_  (.A1(\u_cpu.ALU.u_wallace._2229_ ),
    .A2(\u_cpu.ALU.u_wallace._2230_ ),
    .B1(\u_cpu.ALU.u_wallace._1982_ ),
    .Y(\u_cpu.ALU.u_wallace._2232_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7879_  (.A1(\u_cpu.ALU.u_wallace._1988_ ),
    .A2(\u_cpu.ALU.u_wallace._2232_ ),
    .B1(\u_cpu.ALU.u_wallace._2218_ ),
    .Y(\u_cpu.ALU.u_wallace._2233_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7880_  (.A1(\u_cpu.ALU.u_wallace._0807_ ),
    .A2(\u_cpu.ALU.SrcA[22] ),
    .B1(\u_cpu.ALU.u_wallace._2000_ ),
    .B2(\u_cpu.ALU.u_wallace._1903_ ),
    .X(\u_cpu.ALU.u_wallace._2234_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7881_  (.A(\u_cpu.ALU.u_wallace._4657_ ),
    .B(\u_cpu.ALU.u_wallace._4658_ ),
    .C(\u_cpu.ALU.u_wallace._1734_ ),
    .D(\u_cpu.ALU.u_wallace._2000_ ),
    .Y(\u_cpu.ALU.u_wallace._2235_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7882_  (.A1(\u_cpu.ALU.u_wallace._0840_ ),
    .A2(\u_cpu.ALU.u_wallace._1531_ ),
    .B1(\u_cpu.ALU.u_wallace._2234_ ),
    .B2(\u_cpu.ALU.u_wallace._2235_ ),
    .Y(\u_cpu.ALU.u_wallace._2236_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7883_  (.A1(\u_cpu.ALU.u_wallace._0490_ ),
    .A2(\u_cpu.ALU.SrcA[22] ),
    .B1(\u_cpu.ALU.u_wallace._2000_ ),
    .B2(\u_cpu.ALU.u_wallace._0206_ ),
    .Y(\u_cpu.ALU.u_wallace._2237_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7884_  (.A(\u_cpu.ALU.u_wallace._0457_ ),
    .B(\u_cpu.ALU.u_wallace._1730_ ),
    .Y(\u_cpu.ALU.u_wallace._2238_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7885_  (.A(\u_cpu.ALU.u_wallace._0775_ ),
    .B(\u_cpu.ALU.u_wallace._0534_ ),
    .C(\u_cpu.ALU.SrcA[22] ),
    .D(\u_cpu.ALU.SrcA[23] ),
    .X(\u_cpu.ALU.u_wallace._2239_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._7886_  (.A(\u_cpu.ALU.u_wallace._2237_ ),
    .B(\u_cpu.ALU.u_wallace._2238_ ),
    .C(\u_cpu.ALU.u_wallace._2239_ ),
    .Y(\u_cpu.ALU.u_wallace._2240_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7887_  (.A(\u_cpu.ALU.u_wallace._2236_ ),
    .B(\u_cpu.ALU.u_wallace._2240_ ),
    .Y(\u_cpu.ALU.u_wallace._2241_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7888_  (.A1(\u_cpu.ALU.u_wallace._2228_ ),
    .A2(\u_cpu.ALU.u_wallace._2233_ ),
    .B1(\u_cpu.ALU.u_wallace._2241_ ),
    .Y(\u_cpu.ALU.u_wallace._2243_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7889_  (.A1(\u_cpu.ALU.u_wallace._1988_ ),
    .A2(\u_cpu.ALU.u_wallace._2232_ ),
    .B1(\u_cpu.ALU.u_wallace._2223_ ),
    .C1(\u_cpu.ALU.u_wallace._2218_ ),
    .X(\u_cpu.ALU.u_wallace._2244_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7890_  (.A1(\u_cpu.ALU.u_wallace._2236_ ),
    .A2(\u_cpu.ALU.u_wallace._2240_ ),
    .B1(\u_cpu.ALU.u_wallace._2244_ ),
    .B2(\u_cpu.ALU.u_wallace._2225_ ),
    .Y(\u_cpu.ALU.u_wallace._2245_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7891_  (.A1(\u_cpu.ALU.u_wallace._1989_ ),
    .A2(\u_cpu.ALU.u_wallace._1986_ ),
    .B1(\u_cpu.ALU.u_wallace._2026_ ),
    .B2(\u_cpu.ALU.u_wallace._2009_ ),
    .Y(\u_cpu.ALU.u_wallace._2246_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7892_  (.A1(\u_cpu.ALU.u_wallace._2225_ ),
    .A2(\u_cpu.ALU.u_wallace._2243_ ),
    .B1(\u_cpu.ALU.u_wallace._2245_ ),
    .C1(\u_cpu.ALU.u_wallace._2246_ ),
    .X(\u_cpu.ALU.u_wallace._2247_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7893_  (.A(\u_cpu.ALU.u_wallace._1075_ ),
    .X(\u_cpu.ALU.u_wallace._2248_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7894_  (.A(\u_cpu.ALU.u_wallace._1962_ ),
    .B(\u_cpu.ALU.u_wallace._2248_ ),
    .C(\u_cpu.ALU.u_wallace._0015_ ),
    .X(\u_cpu.ALU.u_wallace._2249_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7895_  (.A(\u_cpu.ALU.u_wallace._0840_ ),
    .B(\u_cpu.ALU.u_wallace._1275_ ),
    .Y(\u_cpu.ALU.u_wallace._2250_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7896_  (.A(\u_cpu.ALU.u_wallace._2250_ ),
    .B(\u_cpu.ALU.u_wallace._1992_ ),
    .Y(\u_cpu.ALU.u_wallace._2251_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7897_  (.A1(\u_cpu.ALU.u_wallace._2078_ ),
    .A2(\u_cpu.ALU.u_wallace._1090_ ),
    .B1(\u_cpu.ALU.u_wallace._1270_ ),
    .B2(\u_cpu.ALU.u_wallace._4467_ ),
    .X(\u_cpu.ALU.u_wallace._2252_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7898_  (.A(\u_cpu.ALU.u_wallace._1530_ ),
    .B(\u_cpu.ALU.u_wallace._2056_ ),
    .C(\u_cpu.ALU.u_wallace._1090_ ),
    .D(\u_cpu.ALU.u_wallace._1543_ ),
    .Y(\u_cpu.ALU.u_wallace._2254_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7899_  (.A(\u_cpu.ALU.u_wallace._2252_ ),
    .B(\u_cpu.ALU.u_wallace._2254_ ),
    .C(\u_cpu.ALU.u_wallace._2626_ ),
    .D(\u_cpu.ALU.u_wallace._1286_ ),
    .Y(\u_cpu.ALU.u_wallace._2255_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7900_  (.A1(\u_cpu.ALU.u_wallace._2056_ ),
    .A2(\u_cpu.ALU.u_wallace._1090_ ),
    .B1(\u_cpu.ALU.u_wallace._1543_ ),
    .B2(\u_cpu.ALU.u_wallace._2045_ ),
    .Y(\u_cpu.ALU.u_wallace._2256_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7901_  (.A(\u_cpu.ALU.u_wallace._1465_ ),
    .B(\u_cpu.ALU.u_wallace._2538_ ),
    .C(\u_cpu.ALU.u_wallace._1100_ ),
    .D(\u_cpu.ALU.u_wallace._1270_ ),
    .X(\u_cpu.ALU.u_wallace._2257_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7902_  (.A1(\u_cpu.ALU.u_wallace._4471_ ),
    .A2(\u_cpu.ALU.u_wallace._0635_ ),
    .B1(\u_cpu.ALU.u_wallace._2256_ ),
    .B2(\u_cpu.ALU.u_wallace._2257_ ),
    .Y(\u_cpu.ALU.u_wallace._2258_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7903_  (.A1(\u_cpu.ALU.u_wallace._1991_ ),
    .A2(\u_cpu.ALU.u_wallace._2251_ ),
    .B1(\u_cpu.ALU.u_wallace._2255_ ),
    .C1(\u_cpu.ALU.u_wallace._2258_ ),
    .Y(\u_cpu.ALU.u_wallace._2259_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7904_  (.A1(\u_cpu.ALU.u_wallace._2250_ ),
    .A2(\u_cpu.ALU.u_wallace._1992_ ),
    .B1(\u_cpu.ALU.u_wallace._1995_ ),
    .Y(\u_cpu.ALU.u_wallace._2260_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7905_  (.A1(\u_cpu.ALU.u_wallace._2255_ ),
    .A2(\u_cpu.ALU.u_wallace._2258_ ),
    .B1(\u_cpu.ALU.u_wallace._2260_ ),
    .X(\u_cpu.ALU.u_wallace._2261_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._7906_  (.A1_N(\u_cpu.ALU.u_wallace._1960_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2249_ ),
    .B1(\u_cpu.ALU.u_wallace._2259_ ),
    .B2(\u_cpu.ALU.u_wallace._2261_ ),
    .Y(\u_cpu.ALU.u_wallace._2262_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._7907_  (.A1(\u_cpu.ALU.u_wallace._1991_ ),
    .A2(\u_cpu.ALU.u_wallace._2251_ ),
    .B1(\u_cpu.ALU.u_wallace._2258_ ),
    .X(\u_cpu.ALU.u_wallace._2263_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7908_  (.A1(\u_cpu.ALU.u_wallace._1962_ ),
    .A2(\u_cpu.ALU.u_wallace._2248_ ),
    .A3(\u_cpu.ALU.u_wallace._0015_ ),
    .B1(\u_cpu.ALU.u_wallace._1960_ ),
    .X(\u_cpu.ALU.u_wallace._2265_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7909_  (.A1(\u_cpu.ALU.u_wallace._2255_ ),
    .A2(\u_cpu.ALU.u_wallace._2258_ ),
    .B1(\u_cpu.ALU.u_wallace._2260_ ),
    .Y(\u_cpu.ALU.u_wallace._2266_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU.u_wallace._7910_  (.A1(\u_cpu.ALU.u_wallace._2263_ ),
    .A2(\u_cpu.ALU.u_wallace._2255_ ),
    .B1(\u_cpu.ALU.u_wallace._2265_ ),
    .C1(\u_cpu.ALU.u_wallace._2266_ ),
    .Y(\u_cpu.ALU.u_wallace._2267_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7911_  (.A1(\u_cpu.ALU.u_wallace._2244_ ),
    .A2(\u_cpu.ALU.u_wallace._2225_ ),
    .B1(\u_cpu.ALU.u_wallace._2241_ ),
    .Y(\u_cpu.ALU.u_wallace._2268_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7912_  (.A1(\u_cpu.ALU.u_wallace._2757_ ),
    .A2(\u_cpu.ALU.u_wallace._2222_ ),
    .B1(\u_cpu.ALU.u_wallace._2219_ ),
    .B2(\u_cpu.ALU.u_wallace._2221_ ),
    .Y(\u_cpu.ALU.u_wallace._2269_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._7913_  (.A1(\u_cpu.ALU.u_wallace._2269_ ),
    .A2(\u_cpu.ALU.u_wallace._2228_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2224_ ),
    .Y(\u_cpu.ALU.u_wallace._2270_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._7914_  (.A1(\u_cpu.ALU.u_wallace._2236_ ),
    .A2(\u_cpu.ALU.u_wallace._2240_ ),
    .B1(\u_cpu.ALU.u_wallace._2228_ ),
    .B2(\u_cpu.ALU.u_wallace._2233_ ),
    .C1(\u_cpu.ALU.u_wallace._2270_ ),
    .Y(\u_cpu.ALU.u_wallace._2271_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._7915_  (.A1(\u_cpu.ALU.u_wallace._1989_ ),
    .A2(\u_cpu.ALU.u_wallace._1986_ ),
    .B1(\u_cpu.ALU.u_wallace._2026_ ),
    .B2(\u_cpu.ALU.u_wallace._2009_ ),
    .X(\u_cpu.ALU.u_wallace._2272_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7916_  (.A(\u_cpu.ALU.u_wallace._2268_ ),
    .B(\u_cpu.ALU.u_wallace._2271_ ),
    .C(\u_cpu.ALU.u_wallace._2272_ ),
    .Y(\u_cpu.ALU.u_wallace._2273_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7917_  (.A1(\u_cpu.ALU.u_wallace._2262_ ),
    .A2(\u_cpu.ALU.u_wallace._2267_ ),
    .B1(\u_cpu.ALU.u_wallace._2273_ ),
    .Y(\u_cpu.ALU.u_wallace._2274_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7918_  (.A1(\u_cpu.ALU.u_wallace._2225_ ),
    .A2(\u_cpu.ALU.u_wallace._2243_ ),
    .B1(\u_cpu.ALU.u_wallace._2245_ ),
    .C1(\u_cpu.ALU.u_wallace._2246_ ),
    .Y(\u_cpu.ALU.u_wallace._2276_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._7919_  (.A(\u_cpu.ALU.u_wallace._2265_ ),
    .B(\u_cpu.ALU.u_wallace._2259_ ),
    .C(\u_cpu.ALU.u_wallace._2261_ ),
    .X(\u_cpu.ALU.u_wallace._2277_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7920_  (.A1(\u_cpu.ALU.u_wallace._2259_ ),
    .A2(\u_cpu.ALU.u_wallace._2261_ ),
    .B1(\u_cpu.ALU.u_wallace._2265_ ),
    .Y(\u_cpu.ALU.u_wallace._2278_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7921_  (.A1_N(\u_cpu.ALU.u_wallace._2276_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2273_ ),
    .B1(\u_cpu.ALU.u_wallace._2277_ ),
    .B2(\u_cpu.ALU.u_wallace._2278_ ),
    .Y(\u_cpu.ALU.u_wallace._2279_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._7922_  (.A1(\u_cpu.ALU.u_wallace._2247_ ),
    .A2(\u_cpu.ALU.u_wallace._2274_ ),
    .B1(\u_cpu.ALU.u_wallace._2022_ ),
    .B2(\u_cpu.ALU.u_wallace._2106_ ),
    .C1(\u_cpu.ALU.u_wallace._2279_ ),
    .Y(\u_cpu.ALU.u_wallace._2280_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7923_  (.A1(\u_cpu.ALU.u_wallace._2262_ ),
    .A2(\u_cpu.ALU.u_wallace._2267_ ),
    .B1(\u_cpu.ALU.u_wallace._2276_ ),
    .C1(\u_cpu.ALU.u_wallace._2273_ ),
    .X(\u_cpu.ALU.u_wallace._2281_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7924_  (.A1(\u_cpu.ALU.u_wallace._1991_ ),
    .A2(\u_cpu.ALU.u_wallace._2251_ ),
    .B1(\u_cpu.ALU.u_wallace._2255_ ),
    .C1(\u_cpu.ALU.u_wallace._2258_ ),
    .X(\u_cpu.ALU.u_wallace._2282_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7925_  (.A1(\u_cpu.ALU.u_wallace._2282_ ),
    .A2(\u_cpu.ALU.u_wallace._2266_ ),
    .B1(\u_cpu.ALU.u_wallace._2265_ ),
    .Y(\u_cpu.ALU.u_wallace._2283_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7926_  (.A(\u_cpu.ALU.u_wallace._4471_ ),
    .X(\u_cpu.ALU.u_wallace._2284_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._7927_  (.A1(\u_cpu.ALU.u_wallace._2284_ ),
    .A2(\u_cpu.ALU.u_wallace._0442_ ),
    .A3(\u_cpu.ALU.u_wallace._1959_ ),
    .B1(\u_cpu.ALU.u_wallace._1963_ ),
    .X(\u_cpu.ALU.u_wallace._2285_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7928_  (.A(\u_cpu.ALU.u_wallace._2261_ ),
    .B(\u_cpu.ALU.u_wallace._2285_ ),
    .C(\u_cpu.ALU.u_wallace._2259_ ),
    .Y(\u_cpu.ALU.u_wallace._2287_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7929_  (.A(\u_cpu.ALU.u_wallace._2283_ ),
    .B(\u_cpu.ALU.u_wallace._2287_ ),
    .Y(\u_cpu.ALU.u_wallace._2288_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7930_  (.A1(\u_cpu.ALU.u_wallace._2276_ ),
    .A2(\u_cpu.ALU.u_wallace._2273_ ),
    .B1(\u_cpu.ALU.u_wallace._2288_ ),
    .Y(\u_cpu.ALU.u_wallace._2289_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._7931_  (.A1(\u_cpu.ALU.u_wallace._1976_ ),
    .A2(\u_cpu.ALU.u_wallace._2031_ ),
    .A3(\u_cpu.ALU.u_wallace._2030_ ),
    .B1(\u_cpu.ALU.u_wallace._2022_ ),
    .Y(\u_cpu.ALU.u_wallace._2290_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7932_  (.A1(\u_cpu.ALU.u_wallace._2281_ ),
    .A2(\u_cpu.ALU.u_wallace._2289_ ),
    .B1(\u_cpu.ALU.u_wallace._2290_ ),
    .Y(\u_cpu.ALU.u_wallace._2291_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._7933_  (.A_N(\u_cpu.ALU.u_wallace._2214_ ),
    .B(\u_cpu.ALU.u_wallace._2280_ ),
    .C(\u_cpu.ALU.u_wallace._2291_ ),
    .Y(\u_cpu.ALU.u_wallace._2292_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7934_  (.A1(\u_cpu.ALU.u_wallace._2191_ ),
    .A2(\u_cpu.ALU.u_wallace._2203_ ),
    .B1(\u_cpu.ALU.u_wallace._2206_ ),
    .C1(\u_cpu.ALU.u_wallace._2170_ ),
    .X(\u_cpu.ALU.u_wallace._2293_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU.u_wallace._7935_  (.A1(\u_cpu.ALU.u_wallace._1945_ ),
    .A2(\u_cpu.ALU.u_wallace._1947_ ),
    .A3(\u_cpu.ALU.u_wallace._1929_ ),
    .B1(\u_cpu.ALU.u_wallace._1938_ ),
    .C1(\u_cpu.ALU.u_wallace._2207_ ),
    .X(\u_cpu.ALU.u_wallace._2294_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._7936_  (.A1(\u_cpu.ALU.u_wallace._2247_ ),
    .A2(\u_cpu.ALU.u_wallace._2274_ ),
    .B1(\u_cpu.ALU.u_wallace._2022_ ),
    .B2(\u_cpu.ALU.u_wallace._2106_ ),
    .C1(\u_cpu.ALU.u_wallace._2279_ ),
    .X(\u_cpu.ALU.u_wallace._2295_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7937_  (.A1(\u_cpu.ALU.u_wallace._2262_ ),
    .A2(\u_cpu.ALU.u_wallace._2267_ ),
    .B1(\u_cpu.ALU.u_wallace._2276_ ),
    .C1(\u_cpu.ALU.u_wallace._2273_ ),
    .Y(\u_cpu.ALU.u_wallace._2296_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7938_  (.A1(\u_cpu.ALU.u_wallace._2032_ ),
    .A2(\u_cpu.ALU.u_wallace._2015_ ),
    .B1(\u_cpu.ALU.u_wallace._2011_ ),
    .Y(\u_cpu.ALU.u_wallace._2298_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7939_  (.A1(\u_cpu.ALU.u_wallace._2296_ ),
    .A2(\u_cpu.ALU.u_wallace._2279_ ),
    .B1(\u_cpu.ALU.u_wallace._2298_ ),
    .Y(\u_cpu.ALU.u_wallace._2299_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._7940_  (.A1(\u_cpu.ALU.u_wallace._2293_ ),
    .A2(\u_cpu.ALU.u_wallace._2294_ ),
    .B1(\u_cpu.ALU.u_wallace._2295_ ),
    .B2(\u_cpu.ALU.u_wallace._2299_ ),
    .Y(\u_cpu.ALU.u_wallace._2300_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7941_  (.A(\u_cpu.ALU.u_wallace._1953_ ),
    .Y(\u_cpu.ALU.u_wallace._2301_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7942_  (.A1(\u_cpu.ALU.u_wallace._1775_ ),
    .A2(\u_cpu.ALU.u_wallace._1942_ ),
    .B1(\u_cpu.ALU.u_wallace._1949_ ),
    .Y(\u_cpu.ALU.u_wallace._2302_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7943_  (.A1(\u_cpu.ALU.u_wallace._1953_ ),
    .A2(\u_cpu.ALU.u_wallace._1949_ ),
    .B1(\u_cpu.ALU.u_wallace._1954_ ),
    .X(\u_cpu.ALU.u_wallace._2303_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7944_  (.A1(\u_cpu.ALU.u_wallace._2301_ ),
    .A2(\u_cpu.ALU.u_wallace._2302_ ),
    .B1(\u_cpu.ALU.u_wallace._2303_ ),
    .Y(\u_cpu.ALU.u_wallace._2304_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._7945_  (.A1_N(\u_cpu.ALU.u_wallace._1951_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2043_ ),
    .B1(\u_cpu.ALU.u_wallace._1922_ ),
    .B2(\u_cpu.ALU.u_wallace._2304_ ),
    .Y(\u_cpu.ALU.u_wallace._2305_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7946_  (.A1(\u_cpu.ALU.u_wallace._2013_ ),
    .A2(\u_cpu.ALU.u_wallace._2015_ ),
    .B1(\u_cpu.ALU.u_wallace._2018_ ),
    .C1(\u_cpu.ALU.u_wallace._2024_ ),
    .X(\u_cpu.ALU.u_wallace._2306_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7947_  (.A1(\u_cpu.ALU.u_wallace._2305_ ),
    .A2(\u_cpu.ALU.u_wallace._2038_ ),
    .B1(\u_cpu.ALU.u_wallace._2306_ ),
    .Y(\u_cpu.ALU.u_wallace._2307_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._7948_  (.A1(\u_cpu.ALU.u_wallace._2292_ ),
    .A2(\u_cpu.ALU.u_wallace._2300_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2307_ ),
    .Y(\u_cpu.ALU.u_wallace._2309_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7949_  (.A1(\u_cpu.ALU.u_wallace._1793_ ),
    .A2(\u_cpu.ALU.u_wallace._0957_ ),
    .B1(\u_cpu.ALU.u_wallace._1210_ ),
    .B2(\u_cpu.ALU.u_wallace._2955_ ),
    .X(\u_cpu.ALU.u_wallace._2310_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7950_  (.A(\u_cpu.ALU.u_wallace._1848_ ),
    .B(\u_cpu.ALU.u_wallace._1125_ ),
    .C(\u_cpu.ALU.u_wallace._1387_ ),
    .D(\u_cpu.ALU.u_wallace._1210_ ),
    .Y(\u_cpu.ALU.u_wallace._2311_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7951_  (.A1(\u_cpu.ALU.u_wallace._2933_ ),
    .A2(\u_cpu.ALU.u_wallace._1386_ ),
    .B1(\u_cpu.ALU.u_wallace._2310_ ),
    .B2(\u_cpu.ALU.u_wallace._2311_ ),
    .X(\u_cpu.ALU.u_wallace._2312_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7952_  (.A(\u_cpu.ALU.u_wallace._2310_ ),
    .B(\u_cpu.ALU.u_wallace._2311_ ),
    .C(\u_cpu.ALU.u_wallace._2933_ ),
    .D(\u_cpu.ALU.u_wallace._1392_ ),
    .Y(\u_cpu.ALU.u_wallace._2313_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7953_  (.A1(\u_cpu.ALU.u_wallace._2049_ ),
    .A2(\u_cpu.ALU.u_wallace._1386_ ),
    .A3(\u_cpu.ALU.u_wallace._4527_ ),
    .B1(\u_cpu.ALU.u_wallace._2055_ ),
    .X(\u_cpu.ALU.u_wallace._2314_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7954_  (.A1(\u_cpu.ALU.u_wallace._2312_ ),
    .A2(\u_cpu.ALU.u_wallace._2313_ ),
    .B1(\u_cpu.ALU.u_wallace._2314_ ),
    .X(\u_cpu.ALU.u_wallace._2315_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7955_  (.A(\u_cpu.ALU.u_wallace._2314_ ),
    .B(\u_cpu.ALU.u_wallace._2312_ ),
    .C(\u_cpu.ALU.u_wallace._2313_ ),
    .Y(\u_cpu.ALU.u_wallace._2316_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7956_  (.A(\u_cpu.ALU.u_wallace._4545_ ),
    .B(\u_cpu.ALU.u_wallace._4527_ ),
    .C(\u_cpu.ALU.SrcB[21] ),
    .D(\u_cpu.ALU.SrcB[22] ),
    .X(\u_cpu.ALU.u_wallace._2317_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7957_  (.A1(\u_cpu.ALU.u_wallace._4541_ ),
    .A2(\u_cpu.ALU.u_wallace._1610_ ),
    .B1(\u_cpu.ALU.u_wallace._1824_ ),
    .B2(\u_cpu.ALU.u_wallace._0370_ ),
    .Y(\u_cpu.ALU.u_wallace._2318_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7958_  (.A(\u_cpu.ALU.u_wallace._2317_ ),
    .B(\u_cpu.ALU.u_wallace._2318_ ),
    .Y(\u_cpu.ALU.u_wallace._2320_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7959_  (.A1(\u_cpu.ALU.u_wallace._2315_ ),
    .A2(\u_cpu.ALU.u_wallace._2316_ ),
    .B1(\u_cpu.ALU.u_wallace._2320_ ),
    .X(\u_cpu.ALU.u_wallace._2321_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7960_  (.A(\u_cpu.ALU.u_wallace._2315_ ),
    .B(\u_cpu.ALU.u_wallace._2316_ ),
    .C(\u_cpu.ALU.u_wallace._2320_ ),
    .Y(\u_cpu.ALU.u_wallace._2322_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._7961_  (.A1(\u_cpu.ALU.u_wallace._2071_ ),
    .A2(\u_cpu.ALU.u_wallace._2075_ ),
    .B1(\u_cpu.ALU.u_wallace._2070_ ),
    .X(\u_cpu.ALU.u_wallace._2323_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7962_  (.A1(\u_cpu.ALU.u_wallace._2069_ ),
    .A2(\u_cpu.ALU.u_wallace._2323_ ),
    .B1(\u_cpu.ALU.u_wallace._2080_ ),
    .B2(\u_cpu.ALU.u_wallace._2077_ ),
    .Y(\u_cpu.ALU.u_wallace._2324_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._7963_  (.A(\u_cpu.ALU.u_wallace._1932_ ),
    .B(\u_cpu.ALU.u_wallace._1943_ ),
    .Y(\u_cpu.ALU.u_wallace._2325_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._7964_  (.A1(\u_cpu.ALU.u_wallace._4550_ ),
    .A2(\u_cpu.ALU.u_wallace._0727_ ),
    .B1(\u_cpu.ALU.u_wallace._0278_ ),
    .B2(\u_cpu.ALU.u_wallace._4401_ ),
    .X(\u_cpu.ALU.u_wallace._2326_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7965_  (.A(\u_cpu.ALU.u_wallace._4562_ ),
    .B(\u_cpu.ALU.u_wallace._4553_ ),
    .C(\u_cpu.ALU.u_wallace._0727_ ),
    .D(\u_cpu.ALU.u_wallace._0728_ ),
    .Y(\u_cpu.ALU.u_wallace._2327_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._7966_  (.A(\u_cpu.ALU.u_wallace._2326_ ),
    .B(\u_cpu.ALU.u_wallace._0550_ ),
    .C(\u_cpu.ALU.u_wallace._4660_ ),
    .D(\u_cpu.ALU.u_wallace._2327_ ),
    .Y(\u_cpu.ALU.u_wallace._2328_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._7967_  (.A1_N(\u_cpu.ALU.u_wallace._2327_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2326_ ),
    .B1(\u_cpu.ALU.u_wallace._4676_ ),
    .B2(\u_cpu.ALU.u_wallace._0941_ ),
    .Y(\u_cpu.ALU.u_wallace._2329_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._7968_  (.A1(\u_cpu.ALU.u_wallace._1944_ ),
    .A2(\u_cpu.ALU.u_wallace._2325_ ),
    .B1(\u_cpu.ALU.u_wallace._2328_ ),
    .C1(\u_cpu.ALU.u_wallace._2329_ ),
    .X(\u_cpu.ALU.u_wallace._2331_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7969_  (.A1(\u_cpu.ALU.u_wallace._1930_ ),
    .A2(\u_cpu.ALU.u_wallace._0363_ ),
    .A3(\u_cpu.ALU.u_wallace._4643_ ),
    .B1(\u_cpu.ALU.u_wallace._1944_ ),
    .X(\u_cpu.ALU.u_wallace._2332_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._7970_  (.A1(\u_cpu.ALU.u_wallace._2328_ ),
    .A2(\u_cpu.ALU.u_wallace._2329_ ),
    .B1(\u_cpu.ALU.u_wallace._2332_ ),
    .Y(\u_cpu.ALU.u_wallace._2333_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7971_  (.A(\u_cpu.ALU.u_wallace._3623_ ),
    .B(\u_cpu.ALU.u_wallace._4412_ ),
    .C(\u_cpu.ALU.u_wallace._0730_ ),
    .D(\u_cpu.ALU.u_wallace._0732_ ),
    .X(\u_cpu.ALU.u_wallace._2334_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._7972_  (.A1(\u_cpu.ALU.u_wallace._2066_ ),
    .A2(\u_cpu.ALU.u_wallace._0735_ ),
    .A3(\u_cpu.ALU.u_wallace._2801_ ),
    .B1(\u_cpu.ALU.u_wallace._2334_ ),
    .X(\u_cpu.ALU.u_wallace._2335_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7973_  (.A1(\u_cpu.ALU.u_wallace._2331_ ),
    .A2(\u_cpu.ALU.u_wallace._2333_ ),
    .B1(\u_cpu.ALU.u_wallace._2335_ ),
    .Y(\u_cpu.ALU.u_wallace._2336_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7974_  (.A1(\u_cpu.ALU.u_wallace._4642_ ),
    .A2(\u_cpu.ALU.u_wallace._0120_ ),
    .B1(\u_cpu.ALU.u_wallace._0732_ ),
    .B2(\u_cpu.ALU.u_wallace._4412_ ),
    .Y(\u_cpu.ALU.u_wallace._2337_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7975_  (.A(\u_cpu.ALU.u_wallace._4449_ ),
    .B(\u_cpu.ALU.u_wallace._0550_ ),
    .Y(\u_cpu.ALU.u_wallace._2338_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._7976_  (.A(\u_cpu.ALU.u_wallace._4444_ ),
    .B(\u_cpu.ALU.u_wallace._4550_ ),
    .C(\u_cpu.ALU.u_wallace._0727_ ),
    .D(\u_cpu.ALU.u_wallace._0278_ ),
    .X(\u_cpu.ALU.u_wallace._2339_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._7977_  (.A(\u_cpu.ALU.u_wallace._2337_ ),
    .B(\u_cpu.ALU.u_wallace._2338_ ),
    .C(\u_cpu.ALU.u_wallace._2339_ ),
    .Y(\u_cpu.ALU.u_wallace._2340_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7978_  (.A1(\u_cpu.ALU.u_wallace._1944_ ),
    .A2(\u_cpu.ALU.u_wallace._2325_ ),
    .B1(\u_cpu.ALU.u_wallace._2329_ ),
    .Y(\u_cpu.ALU.u_wallace._2342_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._7979_  (.A(\u_cpu.ALU.u_wallace._4698_ ),
    .X(\u_cpu.ALU.u_wallace._2343_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._7980_  (.A1(\u_cpu.ALU.u_wallace._2066_ ),
    .A2(\u_cpu.ALU.u_wallace._0551_ ),
    .A3(\u_cpu.ALU.u_wallace._2343_ ),
    .B1(\u_cpu.ALU.u_wallace._2334_ ),
    .Y(\u_cpu.ALU.u_wallace._2344_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7981_  (.A1(\u_cpu.ALU.u_wallace._4669_ ),
    .A2(\u_cpu.ALU.u_wallace._0735_ ),
    .B1(\u_cpu.ALU.u_wallace._2327_ ),
    .B2(\u_cpu.ALU.u_wallace._2326_ ),
    .Y(\u_cpu.ALU.u_wallace._2345_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._7982_  (.A1(\u_cpu.ALU.u_wallace._4904_ ),
    .A2(\u_cpu.ALU.u_wallace._0036_ ),
    .A3(\u_cpu.ALU.u_wallace._1943_ ),
    .B1(\u_cpu.ALU.u_wallace._1931_ ),
    .X(\u_cpu.ALU.u_wallace._2346_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7983_  (.A1(\u_cpu.ALU.u_wallace._2340_ ),
    .A2(\u_cpu.ALU.u_wallace._2345_ ),
    .B1(\u_cpu.ALU.u_wallace._2346_ ),
    .Y(\u_cpu.ALU.u_wallace._2347_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7984_  (.A1(\u_cpu.ALU.u_wallace._2340_ ),
    .A2(\u_cpu.ALU.u_wallace._2342_ ),
    .B1(\u_cpu.ALU.u_wallace._2344_ ),
    .C1(\u_cpu.ALU.u_wallace._2347_ ),
    .Y(\u_cpu.ALU.u_wallace._2348_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._7985_  (.A(\u_cpu.ALU.u_wallace._2324_ ),
    .B(\u_cpu.ALU.u_wallace._2336_ ),
    .C(\u_cpu.ALU.u_wallace._2348_ ),
    .Y(\u_cpu.ALU.u_wallace._2349_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7986_  (.A(\u_cpu.ALU.u_wallace._2069_ ),
    .B(\u_cpu.ALU.u_wallace._2070_ ),
    .Y(\u_cpu.ALU.u_wallace._2350_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._7987_  (.A1(\u_cpu.ALU.u_wallace._4573_ ),
    .A2(\u_cpu.ALU.u_wallace._0037_ ),
    .A3(\u_cpu.ALU.u_wallace._2074_ ),
    .B1(\u_cpu.ALU.u_wallace._1692_ ),
    .X(\u_cpu.ALU.u_wallace._2351_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._7988_  (.A1(\u_cpu.ALU.u_wallace._2350_ ),
    .A2(\u_cpu.ALU.u_wallace._2351_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2077_ ),
    .Y(\u_cpu.ALU.u_wallace._2353_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7989_  (.A1(\u_cpu.ALU.u_wallace._2342_ ),
    .A2(\u_cpu.ALU.u_wallace._2340_ ),
    .B1(\u_cpu.ALU.u_wallace._2335_ ),
    .C1(\u_cpu.ALU.u_wallace._2347_ ),
    .Y(\u_cpu.ALU.u_wallace._2354_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._7990_  (.A1(\u_cpu.ALU.u_wallace._2331_ ),
    .A2(\u_cpu.ALU.u_wallace._2333_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2335_ ),
    .Y(\u_cpu.ALU.u_wallace._2355_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._7991_  (.A1(\u_cpu.ALU.u_wallace._2076_ ),
    .A2(\u_cpu.ALU.u_wallace._2353_ ),
    .B1(\u_cpu.ALU.u_wallace._2354_ ),
    .C1(\u_cpu.ALU.u_wallace._2355_ ),
    .Y(\u_cpu.ALU.u_wallace._2356_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._7992_  (.A1(\u_cpu.ALU.u_wallace._2321_ ),
    .A2(\u_cpu.ALU.u_wallace._2322_ ),
    .B1(\u_cpu.ALU.u_wallace._2349_ ),
    .B2(\u_cpu.ALU.u_wallace._2356_ ),
    .Y(\u_cpu.ALU.u_wallace._2357_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7993_  (.A(\u_cpu.ALU.u_wallace._2315_ ),
    .B(\u_cpu.ALU.u_wallace._2320_ ),
    .Y(\u_cpu.ALU.u_wallace._2358_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._7994_  (.A(\u_cpu.ALU.u_wallace._2316_ ),
    .Y(\u_cpu.ALU.u_wallace._2359_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._7995_  (.A1(\u_cpu.ALU.u_wallace._2358_ ),
    .A2(\u_cpu.ALU.u_wallace._2359_ ),
    .B1(\u_cpu.ALU.u_wallace._2321_ ),
    .C1(\u_cpu.ALU.u_wallace._2349_ ),
    .D1(\u_cpu.ALU.u_wallace._2356_ ),
    .X(\u_cpu.ALU.u_wallace._2360_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._7996_  (.A1(\u_cpu.ALU.u_wallace._2302_ ),
    .A2(\u_cpu.ALU.u_wallace._2301_ ),
    .B1(\u_cpu.ALU.u_wallace._1922_ ),
    .B2(\u_cpu.ALU.u_wallace._1955_ ),
    .X(\u_cpu.ALU.u_wallace._2361_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._7997_  (.A1(\u_cpu.ALU.u_wallace._2357_ ),
    .A2(\u_cpu.ALU.u_wallace._2360_ ),
    .B1(\u_cpu.ALU.u_wallace._2361_ ),
    .Y(\u_cpu.ALU.u_wallace._2362_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._7998_  (.A1(\u_cpu.ALU.u_wallace._2088_ ),
    .A2(\u_cpu.ALU.u_wallace._2091_ ),
    .B1(\u_cpu.ALU.u_wallace._2086_ ),
    .X(\u_cpu.ALU.u_wallace._2364_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._7999_  (.A(\u_cpu.ALU.u_wallace._2362_ ),
    .B(\u_cpu.ALU.u_wallace._2364_ ),
    .Y(\u_cpu.ALU.u_wallace._2365_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8000_  (.A1(\u_cpu.ALU.u_wallace._2041_ ),
    .A2(\u_cpu.ALU.u_wallace._2040_ ),
    .B1(\u_cpu.ALU.u_wallace._1922_ ),
    .Y(\u_cpu.ALU.u_wallace._2366_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8001_  (.A1(\u_cpu.ALU.u_wallace._2321_ ),
    .A2(\u_cpu.ALU.u_wallace._2322_ ),
    .B1(\u_cpu.ALU.u_wallace._2349_ ),
    .B2(\u_cpu.ALU.u_wallace._2356_ ),
    .X(\u_cpu.ALU.u_wallace._2367_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._8002_  (.A1(\u_cpu.ALU.u_wallace._2358_ ),
    .A2(\u_cpu.ALU.u_wallace._2359_ ),
    .B1(\u_cpu.ALU.u_wallace._2321_ ),
    .C1(\u_cpu.ALU.u_wallace._2349_ ),
    .D1(\u_cpu.ALU.u_wallace._2356_ ),
    .Y(\u_cpu.ALU.u_wallace._2368_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8003_  (.A1(\u_cpu.ALU.u_wallace._1951_ ),
    .A2(\u_cpu.ALU.u_wallace._2366_ ),
    .B1(\u_cpu.ALU.u_wallace._2367_ ),
    .C1(\u_cpu.ALU.u_wallace._2368_ ),
    .X(\u_cpu.ALU.u_wallace._2369_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8004_  (.A1(\u_cpu.ALU.u_wallace._1951_ ),
    .A2(\u_cpu.ALU.u_wallace._2366_ ),
    .B1(\u_cpu.ALU.u_wallace._2367_ ),
    .C1(\u_cpu.ALU.u_wallace._2368_ ),
    .Y(\u_cpu.ALU.u_wallace._2370_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8005_  (.A1(\u_cpu.ALU.u_wallace._2362_ ),
    .A2(\u_cpu.ALU.u_wallace._2370_ ),
    .B1(\u_cpu.ALU.u_wallace._2364_ ),
    .X(\u_cpu.ALU.u_wallace._2371_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8006_  (.A(\u_cpu.ALU.u_wallace._2011_ ),
    .B(\u_cpu.ALU.u_wallace._2030_ ),
    .Y(\u_cpu.ALU.u_wallace._2372_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8007_  (.A1_N(\u_cpu.ALU.u_wallace._2032_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2372_ ),
    .B1(\u_cpu.ALU.u_wallace._2013_ ),
    .B2(\u_cpu.ALU.u_wallace._2015_ ),
    .Y(\u_cpu.ALU.u_wallace._2373_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8008_  (.A1(\u_cpu.ALU.u_wallace._1951_ ),
    .A2(\u_cpu.ALU.u_wallace._2043_ ),
    .B1(\u_cpu.ALU.u_wallace._2044_ ),
    .Y(\u_cpu.ALU.u_wallace._2375_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8009_  (.A1(\u_cpu.ALU.u_wallace._2037_ ),
    .A2(\u_cpu.ALU.u_wallace._2373_ ),
    .B1(\u_cpu.ALU.u_wallace._2375_ ),
    .Y(\u_cpu.ALU.u_wallace._2376_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8010_  (.A1(\u_cpu.ALU.u_wallace._2306_ ),
    .A2(\u_cpu.ALU.u_wallace._2376_ ),
    .B1(\u_cpu.ALU.u_wallace._2292_ ),
    .C1(\u_cpu.ALU.u_wallace._2300_ ),
    .Y(\u_cpu.ALU.u_wallace._2377_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8011_  (.A1(\u_cpu.ALU.u_wallace._2365_ ),
    .A2(\u_cpu.ALU.u_wallace._2369_ ),
    .B1(\u_cpu.ALU.u_wallace._2371_ ),
    .C1(\u_cpu.ALU.u_wallace._2377_ ),
    .Y(\u_cpu.ALU.u_wallace._2378_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8012_  (.A1(\u_cpu.ALU.u_wallace._1951_ ),
    .A2(\u_cpu.ALU.u_wallace._2366_ ),
    .B1(\u_cpu.ALU.u_wallace._2367_ ),
    .Y(\u_cpu.ALU.u_wallace._2379_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._8013_  (.A(\u_cpu.ALU.u_wallace._2092_ ),
    .Y(\u_cpu.ALU.u_wallace._2380_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._8014_  (.A1(\u_cpu.ALU.u_wallace._2360_ ),
    .A2(\u_cpu.ALU.u_wallace._2379_ ),
    .B1(\u_cpu.ALU.u_wallace._2086_ ),
    .B2(\u_cpu.ALU.u_wallace._2380_ ),
    .C1(\u_cpu.ALU.u_wallace._2362_ ),
    .Y(\u_cpu.ALU.u_wallace._2381_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._8015_  (.A1(\u_cpu.ALU.u_wallace._2295_ ),
    .A2(\u_cpu.ALU.u_wallace._2299_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2214_ ),
    .Y(\u_cpu.ALU.u_wallace._2382_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8016_  (.A1(\u_cpu.ALU.u_wallace._2293_ ),
    .A2(\u_cpu.ALU.u_wallace._2294_ ),
    .B1(\u_cpu.ALU.u_wallace._2280_ ),
    .C1(\u_cpu.ALU.u_wallace._2291_ ),
    .Y(\u_cpu.ALU.u_wallace._2383_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8017_  (.A(\u_cpu.ALU.u_wallace._2382_ ),
    .B(\u_cpu.ALU.u_wallace._2383_ ),
    .C(\u_cpu.ALU.u_wallace._2307_ ),
    .Y(\u_cpu.ALU.u_wallace._2384_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8018_  (.A1(\u_cpu.ALU.u_wallace._2371_ ),
    .A2(\u_cpu.ALU.u_wallace._2381_ ),
    .B1(\u_cpu.ALU.u_wallace._2384_ ),
    .B2(\u_cpu.ALU.u_wallace._2377_ ),
    .X(\u_cpu.ALU.u_wallace._2386_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8019_  (.A1(\u_cpu.ALU.u_wallace._2309_ ),
    .A2(\u_cpu.ALU.u_wallace._2378_ ),
    .B1(\u_cpu.ALU.u_wallace._2386_ ),
    .Y(\u_cpu.ALU.u_wallace._2387_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8020_  (.A1(\u_cpu.ALU.u_wallace._2099_ ),
    .A2(\u_cpu.ALU.u_wallace._2097_ ),
    .B1(\u_cpu.ALU.u_wallace._2104_ ),
    .Y(\u_cpu.ALU.u_wallace._2388_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.ALU.u_wallace._8021_  (.A1(\u_cpu.ALU.u_wallace._2047_ ),
    .A2(\u_cpu.ALU.u_wallace._2039_ ),
    .A3(\u_cpu.ALU.u_wallace._2046_ ),
    .B1(\u_cpu.ALU.u_wallace._2388_ ),
    .B2(\u_cpu.ALU.u_wallace._2048_ ),
    .X(\u_cpu.ALU.u_wallace._2389_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8022_  (.A(\u_cpu.ALU.u_wallace._4545_ ),
    .B(\u_cpu.ALU.u_wallace._0162_ ),
    .C(\u_cpu.ALU.u_wallace._1610_ ),
    .D(\u_cpu.ALU.u_wallace._1824_ ),
    .X(\u_cpu.ALU.u_wallace._2390_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8023_  (.A1(\u_cpu.ALU.u_wallace._2058_ ),
    .A2(\u_cpu.ALU.u_wallace._2052_ ),
    .A3(\u_cpu.ALU.u_wallace._2057_ ),
    .B1(\u_cpu.ALU.u_wallace._2390_ ),
    .X(\u_cpu.ALU.u_wallace._2391_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8024_  (.A(\u_cpu.ALU.u_wallace._2058_ ),
    .B(\u_cpu.ALU.u_wallace._2052_ ),
    .C(\u_cpu.ALU.u_wallace._2057_ ),
    .D(\u_cpu.ALU.u_wallace._2390_ ),
    .Y(\u_cpu.ALU.u_wallace._2392_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._8025_  (.A1(\u_cpu.ALU.u_wallace._2059_ ),
    .A2(\u_cpu.ALU.u_wallace._2063_ ),
    .A3(\u_cpu.ALU.u_wallace._2060_ ),
    .B1(\u_cpu.ALU.u_wallace._2391_ ),
    .B2(\u_cpu.ALU.u_wallace._2392_ ),
    .X(\u_cpu.ALU.u_wallace._2393_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8026_  (.A1(\u_cpu.ALU.u_wallace._1855_ ),
    .A2(\u_cpu.ALU.u_wallace._2127_ ),
    .A3(\u_cpu.ALU.u_wallace._1825_ ),
    .B1(\u_cpu.ALU.u_wallace._2393_ ),
    .X(\u_cpu.ALU.u_wallace._2394_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8027_  (.A(\u_cpu.ALU.u_wallace._2393_ ),
    .B(\u_cpu.ALU.u_wallace._1825_ ),
    .C(\u_cpu.ALU.u_wallace._2127_ ),
    .D(\u_cpu.ALU.u_wallace._1855_ ),
    .Y(\u_cpu.ALU.u_wallace._2395_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8028_  (.A(\u_cpu.ALU.SrcB[24] ),
    .X(\u_cpu.ALU.u_wallace._2397_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8029_  (.A(\u_cpu.ALU.u_wallace._3996_ ),
    .B(\u_cpu.ALU.u_wallace._2397_ ),
    .Y(\u_cpu.ALU.u_wallace._2398_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8030_  (.A(\u_cpu.ALU.u_wallace._0173_ ),
    .B(\u_cpu.ALU.SrcB[23] ),
    .Y(\u_cpu.ALU.u_wallace._2399_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU.u_wallace._8031_  (.A(\u_cpu.ALU.u_wallace._2398_ ),
    .B(\u_cpu.ALU.u_wallace._2399_ ),
    .X(\u_cpu.ALU.u_wallace._2400_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8032_  (.A(\u_cpu.ALU.u_wallace._2400_ ),
    .X(\u_cpu.ALU.u_wallace._2401_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8033_  (.A(\u_cpu.ALU.u_wallace._2397_ ),
    .X(\u_cpu.ALU.u_wallace._2402_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8034_  (.A1(\u_cpu.ALU.u_wallace._0184_ ),
    .A2(\u_cpu.ALU.u_wallace._2134_ ),
    .B1(\u_cpu.ALU.u_wallace._2402_ ),
    .B2(\u_cpu.ALU.u_wallace._0129_ ),
    .X(\u_cpu.ALU.u_wallace._2403_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8035_  (.A1(\u_cpu.ALU.u_wallace._2394_ ),
    .A2(\u_cpu.ALU.u_wallace._2395_ ),
    .B1(\u_cpu.ALU.u_wallace._2401_ ),
    .B2(\u_cpu.ALU.u_wallace._2403_ ),
    .X(\u_cpu.ALU.u_wallace._2404_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8036_  (.A(\u_cpu.ALU.u_wallace._2394_ ),
    .B(\u_cpu.ALU.u_wallace._2395_ ),
    .C(\u_cpu.ALU.u_wallace._2401_ ),
    .D(\u_cpu.ALU.u_wallace._2403_ ),
    .Y(\u_cpu.ALU.u_wallace._2405_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8037_  (.A(\u_cpu.ALU.u_wallace._2404_ ),
    .B(\u_cpu.ALU.u_wallace._2405_ ),
    .Y(\u_cpu.ALU.u_wallace._2406_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8038_  (.A1(\u_cpu.ALU.u_wallace._2114_ ),
    .A2(\u_cpu.ALU.u_wallace._2097_ ),
    .B1(\u_cpu.ALU.u_wallace._2406_ ),
    .X(\u_cpu.ALU.u_wallace._2408_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8039_  (.A1(\u_cpu.ALU.u_wallace._2093_ ),
    .A2(\u_cpu.ALU.u_wallace._2095_ ),
    .B1(\u_cpu.ALU.u_wallace._2406_ ),
    .C1(\u_cpu.ALU.u_wallace._2097_ ),
    .Y(\u_cpu.ALU.u_wallace._2409_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8040_  (.A(\u_cpu.ALU.u_wallace._2408_ ),
    .B(\u_cpu.ALU.u_wallace._2409_ ),
    .Y(\u_cpu.ALU.u_wallace._2410_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8041_  (.A1(\u_cpu.ALU.u_wallace._2114_ ),
    .A2(\u_cpu.ALU.u_wallace._2097_ ),
    .A3(\u_cpu.ALU.u_wallace._2406_ ),
    .B1(\u_cpu.ALU.u_wallace._2132_ ),
    .X(\u_cpu.ALU.u_wallace._2411_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8042_  (.A1(\u_cpu.ALU.u_wallace._2114_ ),
    .A2(\u_cpu.ALU.u_wallace._2097_ ),
    .B1(\u_cpu.ALU.u_wallace._2406_ ),
    .Y(\u_cpu.ALU.u_wallace._2412_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8043_  (.A1_N(\u_cpu.ALU.u_wallace._2132_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2410_ ),
    .B1(\u_cpu.ALU.u_wallace._2411_ ),
    .B2(\u_cpu.ALU.u_wallace._2412_ ),
    .Y(\u_cpu.ALU.u_wallace._2413_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8044_  (.A1(\u_cpu.ALU.u_wallace._2387_ ),
    .A2(\u_cpu.ALU.u_wallace._2389_ ),
    .B1(\u_cpu.ALU.u_wallace._2413_ ),
    .Y(\u_cpu.ALU.u_wallace._2414_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8045_  (.A1(\u_cpu.ALU.u_wallace._2388_ ),
    .A2(\u_cpu.ALU.u_wallace._2048_ ),
    .B1(\u_cpu.ALU.u_wallace._2110_ ),
    .Y(\u_cpu.ALU.u_wallace._2415_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8046_  (.A1(\u_cpu.ALU.u_wallace._2309_ ),
    .A2(\u_cpu.ALU.u_wallace._2378_ ),
    .B1(\u_cpu.ALU.u_wallace._2386_ ),
    .C1(\u_cpu.ALU.u_wallace._2415_ ),
    .Y(\u_cpu.ALU.u_wallace._2416_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8047_  (.A(\u_cpu.ALU.u_wallace._2134_ ),
    .X(\u_cpu.ALU.u_wallace._2417_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._8048_  (.A1(\u_cpu.ALU.u_wallace._1886_ ),
    .A2(\u_cpu.ALU.u_wallace._2417_ ),
    .A3(\u_cpu.ALU.u_wallace._2135_ ),
    .B1(\u_cpu.ALU.u_wallace._2408_ ),
    .B2(\u_cpu.ALU.u_wallace._2409_ ),
    .X(\u_cpu.ALU.u_wallace._2419_ ));
 sky130_fd_sc_hd__a311o_2 \u_cpu.ALU.u_wallace._8049_  (.A1(\u_cpu.ALU.u_wallace._2114_ ),
    .A2(\u_cpu.ALU.u_wallace._2097_ ),
    .A3(\u_cpu.ALU.u_wallace._2406_ ),
    .B1(\u_cpu.ALU.u_wallace._2132_ ),
    .C1(\u_cpu.ALU.u_wallace._2412_ ),
    .X(\u_cpu.ALU.u_wallace._2420_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8050_  (.A1(\u_cpu.ALU.u_wallace._2362_ ),
    .A2(\u_cpu.ALU.u_wallace._2370_ ),
    .B1(\u_cpu.ALU.u_wallace._2364_ ),
    .Y(\u_cpu.ALU.u_wallace._2421_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._8051_  (.A1(\u_cpu.ALU.u_wallace._2360_ ),
    .A2(\u_cpu.ALU.u_wallace._2379_ ),
    .B1(\u_cpu.ALU.u_wallace._2086_ ),
    .B2(\u_cpu.ALU.u_wallace._2380_ ),
    .C1(\u_cpu.ALU.u_wallace._2362_ ),
    .X(\u_cpu.ALU.u_wallace._2422_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._8052_  (.A1_N(\u_cpu.ALU.u_wallace._2421_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2422_ ),
    .B1(\u_cpu.ALU.u_wallace._2384_ ),
    .B2(\u_cpu.ALU.u_wallace._2377_ ),
    .Y(\u_cpu.ALU.u_wallace._2423_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._8053_  (.A1(\u_cpu.ALU.u_wallace._2365_ ),
    .A2(\u_cpu.ALU.u_wallace._2369_ ),
    .B1(\u_cpu.ALU.u_wallace._2371_ ),
    .C1(\u_cpu.ALU.u_wallace._2384_ ),
    .D1(\u_cpu.ALU.u_wallace._2377_ ),
    .X(\u_cpu.ALU.u_wallace._2424_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._8054_  (.A1(\u_cpu.ALU.u_wallace._2048_ ),
    .A2(\u_cpu.ALU.u_wallace._2388_ ),
    .B1(\u_cpu.ALU.u_wallace._2423_ ),
    .B2(\u_cpu.ALU.u_wallace._2424_ ),
    .C1(\u_cpu.ALU.u_wallace._2110_ ),
    .Y(\u_cpu.ALU.u_wallace._2425_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8055_  (.A1(\u_cpu.ALU.u_wallace._2419_ ),
    .A2(\u_cpu.ALU.u_wallace._2420_ ),
    .B1(\u_cpu.ALU.u_wallace._2425_ ),
    .B2(\u_cpu.ALU.u_wallace._2416_ ),
    .Y(\u_cpu.ALU.u_wallace._2426_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.ALU.u_wallace._8056_  (.A1(\u_cpu.ALU.u_wallace._2119_ ),
    .A2(\u_cpu.ALU.u_wallace._2169_ ),
    .B1(\u_cpu.ALU.u_wallace._2414_ ),
    .B2(\u_cpu.ALU.u_wallace._2416_ ),
    .C1(\u_cpu.ALU.u_wallace._2426_ ),
    .Y(\u_cpu.ALU.u_wallace._2427_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8057_  (.A(\u_cpu.ALU.u_wallace._2119_ ),
    .B(\u_cpu.ALU.u_wallace._2169_ ),
    .Y(\u_cpu.ALU.u_wallace._2428_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8058_  (.A(\u_cpu.ALU.u_wallace._2415_ ),
    .B(\u_cpu.ALU.u_wallace._2386_ ),
    .Y(\u_cpu.ALU.u_wallace._2430_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8059_  (.A1(\u_cpu.ALU.u_wallace._2424_ ),
    .A2(\u_cpu.ALU.u_wallace._2430_ ),
    .B1(\u_cpu.ALU.u_wallace._2425_ ),
    .Y(\u_cpu.ALU.u_wallace._2431_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8060_  (.A1(\u_cpu.ALU.u_wallace._2414_ ),
    .A2(\u_cpu.ALU.u_wallace._2416_ ),
    .B1(\u_cpu.ALU.u_wallace._2413_ ),
    .B2(\u_cpu.ALU.u_wallace._2431_ ),
    .Y(\u_cpu.ALU.u_wallace._2432_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8061_  (.A1(\u_cpu.ALU.u_wallace._2428_ ),
    .A2(\u_cpu.ALU.u_wallace._2432_ ),
    .B1(\u_cpu.ALU.u_wallace._2138_ ),
    .Y(\u_cpu.ALU.u_wallace._2433_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._8062_  (.A(\u_cpu.ALU.u_wallace._2142_ ),
    .Y(\u_cpu.ALU.u_wallace._2434_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8063_  (.A1(\u_cpu.ALU.u_wallace._2389_ ),
    .A2(\u_cpu.ALU.u_wallace._2387_ ),
    .B1(\u_cpu.ALU.u_wallace._2414_ ),
    .Y(\u_cpu.ALU.u_wallace._2435_ ));
 sky130_fd_sc_hd__a32oi_2 \u_cpu.ALU.u_wallace._8064_  (.A1(\u_cpu.ALU.u_wallace._1886_ ),
    .A2(\u_cpu.ALU.u_wallace._2417_ ),
    .A3(\u_cpu.ALU.u_wallace._2135_ ),
    .B1(\u_cpu.ALU.u_wallace._2408_ ),
    .B2(\u_cpu.ALU.u_wallace._2409_ ),
    .Y(\u_cpu.ALU.u_wallace._2436_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8065_  (.A(\u_cpu.ALU.u_wallace._1886_ ),
    .B(\u_cpu.ALU.u_wallace._2417_ ),
    .Y(\u_cpu.ALU.u_wallace._2437_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.ALU.u_wallace._8066_  (.A_N(\u_cpu.ALU.u_wallace._2437_ ),
    .B(\u_cpu.ALU.u_wallace._2135_ ),
    .C(\u_cpu.ALU.u_wallace._2408_ ),
    .D(\u_cpu.ALU.u_wallace._2409_ ),
    .X(\u_cpu.ALU.u_wallace._2438_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._8067_  (.A1(\u_cpu.ALU.u_wallace._2365_ ),
    .A2(\u_cpu.ALU.u_wallace._2369_ ),
    .B1(\u_cpu.ALU.u_wallace._2371_ ),
    .C1(\u_cpu.ALU.u_wallace._2384_ ),
    .D1(\u_cpu.ALU.u_wallace._2377_ ),
    .Y(\u_cpu.ALU.u_wallace._2439_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8068_  (.A1(\u_cpu.ALU.u_wallace._2439_ ),
    .A2(\u_cpu.ALU.u_wallace._2386_ ),
    .B1(\u_cpu.ALU.u_wallace._2415_ ),
    .Y(\u_cpu.ALU.u_wallace._2441_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8069_  (.A1(\u_cpu.ALU.u_wallace._2309_ ),
    .A2(\u_cpu.ALU.u_wallace._2378_ ),
    .B1(\u_cpu.ALU.u_wallace._2386_ ),
    .C1(\u_cpu.ALU.u_wallace._2415_ ),
    .X(\u_cpu.ALU.u_wallace._2442_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8070_  (.A1(\u_cpu.ALU.u_wallace._2436_ ),
    .A2(\u_cpu.ALU.u_wallace._2438_ ),
    .B1(\u_cpu.ALU.u_wallace._2441_ ),
    .B2(\u_cpu.ALU.u_wallace._2442_ ),
    .Y(\u_cpu.ALU.u_wallace._2443_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8071_  (.A1(\u_cpu.ALU.u_wallace._2435_ ),
    .A2(\u_cpu.ALU.u_wallace._2443_ ),
    .B1(\u_cpu.ALU.u_wallace._2428_ ),
    .Y(\u_cpu.ALU.u_wallace._2444_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8072_  (.A1(\u_cpu.ALU.u_wallace._2434_ ),
    .A2(\u_cpu.ALU.u_wallace._2137_ ),
    .B1(\u_cpu.ALU.u_wallace._2427_ ),
    .B2(\u_cpu.ALU.u_wallace._2444_ ),
    .Y(\u_cpu.ALU.u_wallace._2445_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8073_  (.A1(\u_cpu.ALU.u_wallace._2427_ ),
    .A2(\u_cpu.ALU.u_wallace._2433_ ),
    .B1(\u_cpu.ALU.u_wallace._2445_ ),
    .Y(\u_cpu.ALU.u_wallace._2446_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._8074_  (.A1(\u_cpu.ALU.u_wallace._1889_ ),
    .A2(\u_cpu.ALU.u_wallace._2152_ ),
    .A3(\u_cpu.ALU.u_wallace._2150_ ),
    .B1(\u_cpu.ALU.u_wallace._2153_ ),
    .X(\u_cpu.ALU.u_wallace._2447_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8075_  (.A1(\u_cpu.ALU.u_wallace._2446_ ),
    .A2(\u_cpu.ALU.u_wallace._2447_ ),
    .B1(\u_cpu.ALU.u_wallace._2162_ ),
    .Y(\u_cpu.ALU.u_wallace._2448_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU.u_wallace._8076_  (.A(\u_cpu.ALU.u_wallace._2447_ ),
    .B(\u_cpu.ALU.u_wallace._2446_ ),
    .X(\u_cpu.ALU.u_wallace._2449_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8077_  (.A(\u_cpu.ALU.u_wallace._2159_ ),
    .B(\u_cpu.ALU.u_wallace._2160_ ),
    .C(\u_cpu.ALU.u_wallace._2161_ ),
    .X(\u_cpu.ALU.u_wallace._2450_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8078_  (.A(\u_cpu.ALU.u_wallace._2447_ ),
    .B(\u_cpu.ALU.u_wallace._2446_ ),
    .Y(\u_cpu.ALU.u_wallace._2452_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU.u_wallace._8079_  (.A1(\u_cpu.ALU.u_wallace._1889_ ),
    .A2(\u_cpu.ALU.u_wallace._2152_ ),
    .A3(\u_cpu.ALU.u_wallace._2150_ ),
    .B1(\u_cpu.ALU.u_wallace._2446_ ),
    .C1(\u_cpu.ALU.u_wallace._2153_ ),
    .X(\u_cpu.ALU.u_wallace._2453_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8080_  (.A(\u_cpu.ALU.u_wallace._2452_ ),
    .B(\u_cpu.ALU.u_wallace._2453_ ),
    .Y(\u_cpu.ALU.u_wallace._2454_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8081_  (.A1_N(\u_cpu.ALU.u_wallace._2448_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2449_ ),
    .B1(\u_cpu.ALU.u_wallace._2450_ ),
    .B2(\u_cpu.ALU.u_wallace._2454_ ),
    .Y(\u_cpu.ALU.u_wallace._2455_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8082_  (.A1_N(\u_cpu.ALU.u_wallace._1685_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1683_ ),
    .B1(\u_cpu.ALU.u_wallace._1919_ ),
    .B2(\u_cpu.ALU.u_wallace._1918_ ),
    .Y(\u_cpu.ALU.u_wallace._2456_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8083_  (.A1(\u_cpu.ALU.u_wallace._1910_ ),
    .A2(\u_cpu.ALU.u_wallace._1916_ ),
    .B1(\u_cpu.ALU.u_wallace._2163_ ),
    .Y(\u_cpu.ALU.u_wallace._2457_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8084_  (.A1(\u_cpu.ALU.u_wallace._1446_ ),
    .A2(\u_cpu.ALU.u_wallace._1453_ ),
    .A3(\u_cpu.ALU.u_wallace._1687_ ),
    .B1(\u_cpu.ALU.u_wallace._1457_ ),
    .X(\u_cpu.ALU.u_wallace._2458_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8085_  (.A(\u_cpu.ALU.u_wallace._1913_ ),
    .B(\u_cpu.ALU.u_wallace._1915_ ),
    .Y(\u_cpu.ALU.u_wallace._2459_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU.u_wallace._8086_  (.A1(\u_cpu.ALU.u_wallace._1674_ ),
    .A2(\u_cpu.ALU.u_wallace._2458_ ),
    .B1(\u_cpu.ALU.u_wallace._2459_ ),
    .C1(\u_cpu.ALU.u_wallace._2163_ ),
    .Y(\u_cpu.ALU.u_wallace._2460_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8087_  (.A1(\u_cpu.ALU.u_wallace._2456_ ),
    .A2(\u_cpu.ALU.u_wallace._2457_ ),
    .B1(\u_cpu.ALU.u_wallace._2460_ ),
    .Y(\u_cpu.ALU.u_wallace._2461_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8088_  (.A(\u_cpu.ALU.u_wallace._1461_ ),
    .B(\u_cpu.ALU.u_wallace._1466_ ),
    .Y(\u_cpu.ALU.u_wallace._2463_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._8089_  (.A(\u_cpu.ALU.u_wallace._2463_ ),
    .B(\u_cpu.ALU.u_wallace._1683_ ),
    .X(\u_cpu.ALU.u_wallace._2464_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8090_  (.A(\u_cpu.ALU.u_wallace._1474_ ),
    .B(\u_cpu.ALU.u_wallace._2457_ ),
    .C(\u_cpu.ALU.u_wallace._2464_ ),
    .Y(\u_cpu.ALU.u_wallace._2465_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._8091_  (.A_N(\u_cpu.ALU.u_wallace._2163_ ),
    .B(\u_cpu.ALU.u_wallace._1917_ ),
    .C(\u_cpu.ALU.u_wallace._1683_ ),
    .D(\u_cpu.ALU.u_wallace._2463_ ),
    .Y(\u_cpu.ALU.u_wallace._2466_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._8092_  (.A_N(\u_cpu.ALU.u_wallace._2466_ ),
    .B(\u_cpu.ALU.u_wallace._0601_ ),
    .C(\u_cpu.ALU.u_wallace._0595_ ),
    .D(\u_cpu.ALU.u_wallace._1468_ ),
    .Y(\u_cpu.ALU.u_wallace._2467_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8093_  (.A(\u_cpu.ALU.u_wallace._2467_ ),
    .B(\u_cpu.ALU.u_wallace._2461_ ),
    .C(\u_cpu.ALU.u_wallace._2465_ ),
    .Y(\u_cpu.ALU.u_wallace._2468_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._8094_  (.A1(\u_cpu.ALU.u_wallace._2450_ ),
    .A2(\u_cpu.ALU.u_wallace._2454_ ),
    .B1(\u_cpu.ALU.u_wallace._2468_ ),
    .X(\u_cpu.ALU.u_wallace._2469_ ));
 sky130_fd_sc_hd__a41oi_2 \u_cpu.ALU.u_wallace._8095_  (.A1(\u_cpu.ALU.u_wallace._2455_ ),
    .A2(\u_cpu.ALU.u_wallace._2461_ ),
    .A3(\u_cpu.ALU.u_wallace._2465_ ),
    .A4(\u_cpu.ALU.u_wallace._2467_ ),
    .B1(\u_cpu.ALU.u_wallace._2469_ ),
    .Y(\u_cpu.ALU.Product_Wallace[24] ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8096_  (.A1(\u_cpu.ALU.u_wallace._2449_ ),
    .A2(\u_cpu.ALU.u_wallace._2448_ ),
    .B1(\u_cpu.ALU.u_wallace._2469_ ),
    .X(\u_cpu.ALU.u_wallace._2470_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._8097_  (.A(\u_cpu.ALU.u_wallace._2138_ ),
    .Y(\u_cpu.ALU.u_wallace._2471_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._8098_  (.A1(\u_cpu.ALU.u_wallace._2471_ ),
    .A2(\u_cpu.ALU.u_wallace._2444_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2427_ ),
    .Y(\u_cpu.ALU.u_wallace._2473_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8099_  (.A(\u_cpu.ALU.u_wallace._2409_ ),
    .B(\u_cpu.ALU.u_wallace._2417_ ),
    .C(\u_cpu.ALU.u_wallace._1886_ ),
    .D(\u_cpu.ALU.u_wallace._2135_ ),
    .X(\u_cpu.ALU.u_wallace._2474_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8100_  (.A1(\u_cpu.ALU.u_wallace._2314_ ),
    .A2(\u_cpu.ALU.u_wallace._2312_ ),
    .A3(\u_cpu.ALU.u_wallace._2313_ ),
    .B1(\u_cpu.ALU.u_wallace._2317_ ),
    .X(\u_cpu.ALU.u_wallace._2475_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8101_  (.A(\u_cpu.ALU.u_wallace._2314_ ),
    .B(\u_cpu.ALU.u_wallace._2312_ ),
    .C(\u_cpu.ALU.u_wallace._2313_ ),
    .D(\u_cpu.ALU.u_wallace._2317_ ),
    .Y(\u_cpu.ALU.u_wallace._2476_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8102_  (.A(\u_cpu.ALU.u_wallace._2475_ ),
    .B(\u_cpu.ALU.u_wallace._2476_ ),
    .Y(\u_cpu.ALU.u_wallace._2477_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._8103_  (.A1(\u_cpu.ALU.u_wallace._2322_ ),
    .A2(\u_cpu.ALU.u_wallace._2477_ ),
    .B1(\u_cpu.ALU.u_wallace._2060_ ),
    .C1(\u_cpu.ALU.u_wallace._2061_ ),
    .X(\u_cpu.ALU.u_wallace._2478_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8104_  (.A1(\u_cpu.ALU.u_wallace._2060_ ),
    .A2(\u_cpu.ALU.u_wallace._2061_ ),
    .B1(\u_cpu.ALU.u_wallace._2322_ ),
    .C1(\u_cpu.ALU.u_wallace._2477_ ),
    .Y(\u_cpu.ALU.u_wallace._2479_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8105_  (.A(\u_cpu.ALU.SrcB[25] ),
    .X(\u_cpu.ALU.u_wallace._2480_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._8106_  (.A(\u_cpu.ALU.u_wallace._2480_ ),
    .Y(\u_cpu.ALU.u_wallace._2481_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8107_  (.A(\u_cpu.ALU.u_wallace._2481_ ),
    .X(\u_cpu.ALU.u_wallace._2482_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8108_  (.A(\u_cpu.ALU.u_wallace._0118_ ),
    .B(\u_cpu.ALU.u_wallace._0272_ ),
    .C(\u_cpu.ALU.u_wallace._2397_ ),
    .Y(\u_cpu.ALU.u_wallace._2484_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8109_  (.A1(\u_cpu.ALU.u_wallace._0173_ ),
    .A2(\u_cpu.ALU.u_wallace._2397_ ),
    .B1(\u_cpu.ALU.u_wallace._2480_ ),
    .B2(\u_cpu.ALU.u_wallace._0118_ ),
    .X(\u_cpu.ALU.u_wallace._2485_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._8110_  (.A1(\u_cpu.ALU.u_wallace._2482_ ),
    .A2(\u_cpu.ALU.u_wallace._2484_ ),
    .B1(\u_cpu.ALU.u_wallace._0370_ ),
    .C1(\u_cpu.ALU.u_wallace._2134_ ),
    .D1(\u_cpu.ALU.u_wallace._2485_ ),
    .X(\u_cpu.ALU.u_wallace._2486_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU.u_wallace._8111_  (.A1_N(\u_cpu.ALU.u_wallace._0173_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2397_ ),
    .B1(\u_cpu.ALU.u_wallace._2482_ ),
    .B2(\u_cpu.ALU.u_wallace._0043_ ),
    .X(\u_cpu.ALU.u_wallace._2487_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8112_  (.A(\u_cpu.ALU.u_wallace._0108_ ),
    .B(\u_cpu.ALU.u_wallace._4463_ ),
    .C(\u_cpu.ALU.SrcB[24] ),
    .D(\u_cpu.ALU.u_wallace._2480_ ),
    .X(\u_cpu.ALU.u_wallace._2488_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._8113_  (.A1(\u_cpu.ALU.u_wallace._0414_ ),
    .A2(\u_cpu.ALU.u_wallace._2131_ ),
    .B1(\u_cpu.ALU.u_wallace._2487_ ),
    .B2(\u_cpu.ALU.u_wallace._2488_ ),
    .X(\u_cpu.ALU.u_wallace._2489_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8114_  (.A(\u_cpu.ALU.u_wallace._2486_ ),
    .B(\u_cpu.ALU.u_wallace._2489_ ),
    .Y(\u_cpu.ALU.u_wallace._2490_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8115_  (.A1(\u_cpu.ALU.u_wallace._2478_ ),
    .A2(\u_cpu.ALU.u_wallace._2479_ ),
    .B1(\u_cpu.ALU.u_wallace._2490_ ),
    .X(\u_cpu.ALU.u_wallace._2491_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8116_  (.A(\u_cpu.ALU.u_wallace._2478_ ),
    .B(\u_cpu.ALU.u_wallace._2479_ ),
    .C(\u_cpu.ALU.u_wallace._2490_ ),
    .Y(\u_cpu.ALU.u_wallace._2492_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8117_  (.A(\u_cpu.ALU.u_wallace._2491_ ),
    .B(\u_cpu.ALU.u_wallace._2492_ ),
    .Y(\u_cpu.ALU.u_wallace._2493_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8118_  (.A(\u_cpu.ALU.u_wallace._2370_ ),
    .B(\u_cpu.ALU.u_wallace._2365_ ),
    .C(\u_cpu.ALU.u_wallace._2493_ ),
    .X(\u_cpu.ALU.u_wallace._2495_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8119_  (.A1(\u_cpu.ALU.u_wallace._2362_ ),
    .A2(\u_cpu.ALU.u_wallace._2364_ ),
    .B1(\u_cpu.ALU.u_wallace._2369_ ),
    .Y(\u_cpu.ALU.u_wallace._2496_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.ALU.u_wallace._8120_  (.A1_N(\u_cpu.ALU.u_wallace._2493_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2496_ ),
    .B1(\u_cpu.ALU.u_wallace._2405_ ),
    .B2(\u_cpu.ALU.u_wallace._2395_ ),
    .X(\u_cpu.ALU.u_wallace._2497_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8121_  (.A1(\u_cpu.ALU.u_wallace._2370_ ),
    .A2(\u_cpu.ALU.u_wallace._2365_ ),
    .B1(\u_cpu.ALU.u_wallace._2493_ ),
    .Y(\u_cpu.ALU.u_wallace._2498_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._8122_  (.A(\u_cpu.ALU.u_wallace._2395_ ),
    .B(\u_cpu.ALU.u_wallace._2405_ ),
    .X(\u_cpu.ALU.u_wallace._2499_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8123_  (.A1(\u_cpu.ALU.u_wallace._2498_ ),
    .A2(\u_cpu.ALU.u_wallace._2495_ ),
    .B1(\u_cpu.ALU.u_wallace._2499_ ),
    .Y(\u_cpu.ALU.u_wallace._2500_ ));
 sky130_fd_sc_hd__a311oi_2 \u_cpu.ALU.u_wallace._8124_  (.A1(\u_cpu.ALU.u_wallace._2298_ ),
    .A2(\u_cpu.ALU.u_wallace._2296_ ),
    .A3(\u_cpu.ALU.u_wallace._2279_ ),
    .B1(\u_cpu.ALU.u_wallace._2214_ ),
    .C1(\u_cpu.ALU.u_wallace._2299_ ),
    .Y(\u_cpu.ALU.u_wallace._2501_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._8125_  (.A1(\u_cpu.ALU.u_wallace._2293_ ),
    .A2(\u_cpu.ALU.u_wallace._2294_ ),
    .B1(\u_cpu.ALU.u_wallace._2295_ ),
    .B2(\u_cpu.ALU.u_wallace._2299_ ),
    .X(\u_cpu.ALU.u_wallace._2502_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8126_  (.A1(\u_cpu.ALU.u_wallace._2369_ ),
    .A2(\u_cpu.ALU.u_wallace._2365_ ),
    .B1(\u_cpu.ALU.u_wallace._2371_ ),
    .Y(\u_cpu.ALU.u_wallace._2503_ ));
 sky130_fd_sc_hd__o32ai_2 \u_cpu.ALU.u_wallace._8127_  (.A1(\u_cpu.ALU.u_wallace._2307_ ),
    .A2(\u_cpu.ALU.u_wallace._2501_ ),
    .A3(\u_cpu.ALU.u_wallace._2502_ ),
    .B1(\u_cpu.ALU.u_wallace._2503_ ),
    .B2(\u_cpu.ALU.u_wallace._2309_ ),
    .Y(\u_cpu.ALU.u_wallace._2504_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8128_  (.A1(\u_cpu.ALU.u_wallace._4450_ ),
    .A2(\u_cpu.ALU.u_wallace._0957_ ),
    .B1(\u_cpu.ALU.u_wallace._1210_ ),
    .B2(\u_cpu.ALU.u_wallace._3777_ ),
    .X(\u_cpu.ALU.u_wallace._2506_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8129_  (.A(\u_cpu.ALU.u_wallace._2725_ ),
    .B(\u_cpu.ALU.u_wallace._3832_ ),
    .C(\u_cpu.ALU.u_wallace._1387_ ),
    .D(\u_cpu.ALU.u_wallace._1210_ ),
    .Y(\u_cpu.ALU.u_wallace._2507_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8130_  (.A(\u_cpu.ALU.u_wallace._2506_ ),
    .B(\u_cpu.ALU.u_wallace._1392_ ),
    .C(\u_cpu.ALU.u_wallace._1136_ ),
    .D(\u_cpu.ALU.u_wallace._2507_ ),
    .Y(\u_cpu.ALU.u_wallace._2508_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8131_  (.A1(\u_cpu.ALU.u_wallace._1136_ ),
    .A2(\u_cpu.ALU.u_wallace._1386_ ),
    .B1(\u_cpu.ALU.u_wallace._2507_ ),
    .B2(\u_cpu.ALU.u_wallace._2506_ ),
    .X(\u_cpu.ALU.u_wallace._2509_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8132_  (.A(\u_cpu.ALU.u_wallace._3832_ ),
    .B(\u_cpu.ALU.u_wallace._1979_ ),
    .C(\u_cpu.ALU.u_wallace._1387_ ),
    .D(\u_cpu.ALU.u_wallace._1210_ ),
    .X(\u_cpu.ALU.u_wallace._2510_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8133_  (.A1(\u_cpu.ALU.u_wallace._2310_ ),
    .A2(\u_cpu.ALU.u_wallace._1392_ ),
    .A3(\u_cpu.ALU.u_wallace._2933_ ),
    .B1(\u_cpu.ALU.u_wallace._2510_ ),
    .X(\u_cpu.ALU.u_wallace._2511_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8134_  (.A1(\u_cpu.ALU.u_wallace._2508_ ),
    .A2(\u_cpu.ALU.u_wallace._2509_ ),
    .B1(\u_cpu.ALU.u_wallace._2511_ ),
    .X(\u_cpu.ALU.u_wallace._2512_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8135_  (.A(\u_cpu.ALU.u_wallace._2511_ ),
    .B(\u_cpu.ALU.u_wallace._2508_ ),
    .C(\u_cpu.ALU.u_wallace._2509_ ),
    .Y(\u_cpu.ALU.u_wallace._2513_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8136_  (.A(\u_cpu.ALU.u_wallace._0917_ ),
    .B(\u_cpu.ALU.u_wallace._4527_ ),
    .C(\u_cpu.ALU.u_wallace._1610_ ),
    .D(\u_cpu.ALU.SrcB[22] ),
    .X(\u_cpu.ALU.u_wallace._2514_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8137_  (.A1(\u_cpu.ALU.u_wallace._0917_ ),
    .A2(\u_cpu.ALU.u_wallace._1610_ ),
    .B1(\u_cpu.ALU.u_wallace._1824_ ),
    .B2(\u_cpu.ALU.u_wallace._4541_ ),
    .Y(\u_cpu.ALU.u_wallace._2515_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8138_  (.A(\u_cpu.ALU.u_wallace._2514_ ),
    .B(\u_cpu.ALU.u_wallace._2515_ ),
    .Y(\u_cpu.ALU.u_wallace._2517_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8139_  (.A1(\u_cpu.ALU.u_wallace._2512_ ),
    .A2(\u_cpu.ALU.u_wallace._2513_ ),
    .B1(\u_cpu.ALU.u_wallace._2517_ ),
    .X(\u_cpu.ALU.u_wallace._2518_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8140_  (.A(\u_cpu.ALU.u_wallace._2512_ ),
    .B(\u_cpu.ALU.u_wallace._2513_ ),
    .C(\u_cpu.ALU.u_wallace._2517_ ),
    .Y(\u_cpu.ALU.u_wallace._2519_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._8141_  (.A1_N(\u_cpu.ALU.u_wallace._2342_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2340_ ),
    .B1(\u_cpu.ALU.u_wallace._2335_ ),
    .B2(\u_cpu.ALU.u_wallace._2347_ ),
    .Y(\u_cpu.ALU.u_wallace._2520_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8142_  (.A(\u_cpu.ALU.u_wallace._2326_ ),
    .B(\u_cpu.ALU.u_wallace._0551_ ),
    .C(\u_cpu.ALU.u_wallace._4661_ ),
    .X(\u_cpu.ALU.u_wallace._2521_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8143_  (.A(\u_cpu.ALU.u_wallace._4787_ ),
    .B(\u_cpu.ALU.u_wallace._0029_ ),
    .Y(\u_cpu.ALU.u_wallace._2522_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8144_  (.A(\u_cpu.ALU.u_wallace._0028_ ),
    .B(\u_cpu.ALU.u_wallace._4921_ ),
    .Y(\u_cpu.ALU.u_wallace._2523_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8145_  (.A1(\u_cpu.ALU.u_wallace._2522_ ),
    .A2(\u_cpu.ALU.u_wallace._2523_ ),
    .B1(\u_cpu.ALU.u_wallace._2186_ ),
    .Y(\u_cpu.ALU.u_wallace._2524_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8146_  (.A1(\u_cpu.ALU.u_wallace._4650_ ),
    .A2(\u_cpu.ALU.u_wallace._0727_ ),
    .B1(\u_cpu.ALU.u_wallace._0728_ ),
    .B2(\u_cpu.ALU.u_wallace._4553_ ),
    .X(\u_cpu.ALU.u_wallace._2525_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8147_  (.A(\u_cpu.ALU.u_wallace._4642_ ),
    .B(\u_cpu.ALU.u_wallace._4797_ ),
    .C(\u_cpu.ALU.u_wallace._0120_ ),
    .D(\u_cpu.ALU.u_wallace._0728_ ),
    .Y(\u_cpu.ALU.u_wallace._2526_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8148_  (.A(\u_cpu.ALU.u_wallace._2525_ ),
    .B(\u_cpu.ALU.u_wallace._2526_ ),
    .C(\u_cpu.ALU.u_wallace._4567_ ),
    .D(\u_cpu.ALU.u_wallace._0550_ ),
    .Y(\u_cpu.ALU.u_wallace._2528_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8149_  (.A1(\u_cpu.ALU.u_wallace._4647_ ),
    .A2(\u_cpu.ALU.u_wallace._0120_ ),
    .B1(\u_cpu.ALU.u_wallace._0732_ ),
    .B2(\u_cpu.ALU.u_wallace._4642_ ),
    .Y(\u_cpu.ALU.u_wallace._2529_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8150_  (.A(\u_cpu.ALU.u_wallace._4553_ ),
    .B(\u_cpu.ALU.u_wallace._4650_ ),
    .C(\u_cpu.ALU.u_wallace._0727_ ),
    .D(\u_cpu.ALU.u_wallace._0278_ ),
    .X(\u_cpu.ALU.u_wallace._2530_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8151_  (.A1(\u_cpu.ALU.u_wallace._4573_ ),
    .A2(\u_cpu.ALU.u_wallace._0941_ ),
    .B1(\u_cpu.ALU.u_wallace._2529_ ),
    .B2(\u_cpu.ALU.u_wallace._2530_ ),
    .Y(\u_cpu.ALU.u_wallace._2531_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8152_  (.A1(\u_cpu.ALU.u_wallace._2197_ ),
    .A2(\u_cpu.ALU.u_wallace._2524_ ),
    .B1(\u_cpu.ALU.u_wallace._2528_ ),
    .C1(\u_cpu.ALU.u_wallace._2531_ ),
    .X(\u_cpu.ALU.u_wallace._2532_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8153_  (.A1(\u_cpu.ALU.u_wallace._2186_ ),
    .A2(\u_cpu.ALU.u_wallace._2199_ ),
    .B1(\u_cpu.ALU.u_wallace._2183_ ),
    .Y(\u_cpu.ALU.u_wallace._2533_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8154_  (.A1(\u_cpu.ALU.u_wallace._2528_ ),
    .A2(\u_cpu.ALU.u_wallace._2531_ ),
    .B1(\u_cpu.ALU.u_wallace._2533_ ),
    .Y(\u_cpu.ALU.u_wallace._2534_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8155_  (.A1(\u_cpu.ALU.u_wallace._2339_ ),
    .A2(\u_cpu.ALU.u_wallace._2521_ ),
    .B1(\u_cpu.ALU.u_wallace._2532_ ),
    .B2(\u_cpu.ALU.u_wallace._2534_ ),
    .Y(\u_cpu.ALU.u_wallace._2535_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8156_  (.A1(\u_cpu.ALU.u_wallace._2528_ ),
    .A2(\u_cpu.ALU.u_wallace._2531_ ),
    .B1(\u_cpu.ALU.u_wallace._2533_ ),
    .X(\u_cpu.ALU.u_wallace._2536_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._8157_  (.A1(\u_cpu.ALU.u_wallace._4677_ ),
    .A2(\u_cpu.ALU.u_wallace._0554_ ),
    .A3(\u_cpu.ALU.u_wallace._2337_ ),
    .B1(\u_cpu.ALU.u_wallace._2327_ ),
    .X(\u_cpu.ALU.u_wallace._2537_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8158_  (.A1(\u_cpu.ALU.u_wallace._2197_ ),
    .A2(\u_cpu.ALU.u_wallace._2524_ ),
    .B1(\u_cpu.ALU.u_wallace._2528_ ),
    .C1(\u_cpu.ALU.u_wallace._2531_ ),
    .Y(\u_cpu.ALU.u_wallace._2539_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8159_  (.A(\u_cpu.ALU.u_wallace._2536_ ),
    .B(\u_cpu.ALU.u_wallace._2537_ ),
    .C(\u_cpu.ALU.u_wallace._2539_ ),
    .Y(\u_cpu.ALU.u_wallace._2540_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8160_  (.A(\u_cpu.ALU.u_wallace._2520_ ),
    .B(\u_cpu.ALU.u_wallace._2535_ ),
    .C(\u_cpu.ALU.u_wallace._2540_ ),
    .Y(\u_cpu.ALU.u_wallace._2541_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8161_  (.A(\u_cpu.ALU.u_wallace._2066_ ),
    .B(\u_cpu.ALU.u_wallace._0551_ ),
    .C(\u_cpu.ALU.u_wallace._4698_ ),
    .Y(\u_cpu.ALU.u_wallace._2542_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8162_  (.A(\u_cpu.ALU.u_wallace._2328_ ),
    .B(\u_cpu.ALU.u_wallace._2329_ ),
    .Y(\u_cpu.ALU.u_wallace._2543_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8163_  (.A1(\u_cpu.ALU.u_wallace._2068_ ),
    .A2(\u_cpu.ALU.u_wallace._2542_ ),
    .B1(\u_cpu.ALU.u_wallace._2543_ ),
    .B2(\u_cpu.ALU.u_wallace._2346_ ),
    .Y(\u_cpu.ALU.u_wallace._2544_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8164_  (.A1(\u_cpu.ALU.u_wallace._2339_ ),
    .A2(\u_cpu.ALU.u_wallace._2521_ ),
    .B1(\u_cpu.ALU.u_wallace._2539_ ),
    .C1(\u_cpu.ALU.u_wallace._2536_ ),
    .Y(\u_cpu.ALU.u_wallace._2545_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8165_  (.A1(\u_cpu.ALU.u_wallace._2532_ ),
    .A2(\u_cpu.ALU.u_wallace._2534_ ),
    .B1(\u_cpu.ALU.u_wallace._2537_ ),
    .Y(\u_cpu.ALU.u_wallace._2546_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8166_  (.A1(\u_cpu.ALU.u_wallace._2331_ ),
    .A2(\u_cpu.ALU.u_wallace._2544_ ),
    .B1(\u_cpu.ALU.u_wallace._2545_ ),
    .C1(\u_cpu.ALU.u_wallace._2546_ ),
    .Y(\u_cpu.ALU.u_wallace._2547_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8167_  (.A1(\u_cpu.ALU.u_wallace._2518_ ),
    .A2(\u_cpu.ALU.u_wallace._2519_ ),
    .B1(\u_cpu.ALU.u_wallace._2541_ ),
    .B2(\u_cpu.ALU.u_wallace._2547_ ),
    .Y(\u_cpu.ALU.u_wallace._2548_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8168_  (.A(\u_cpu.ALU.u_wallace._2506_ ),
    .B(\u_cpu.ALU.u_wallace._1392_ ),
    .C(\u_cpu.ALU.u_wallace._1136_ ),
    .D(\u_cpu.ALU.u_wallace._2507_ ),
    .X(\u_cpu.ALU.u_wallace._2550_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8169_  (.A(\u_cpu.ALU.u_wallace._2801_ ),
    .B(\u_cpu.ALU.u_wallace._4452_ ),
    .C(\u_cpu.ALU.u_wallace._2050_ ),
    .D(\u_cpu.ALU.u_wallace._1175_ ),
    .X(\u_cpu.ALU.u_wallace._2551_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8170_  (.A1(\u_cpu.ALU.u_wallace._3821_ ),
    .A2(\u_cpu.ALU.u_wallace._2050_ ),
    .B1(\u_cpu.ALU.u_wallace._1175_ ),
    .B2(\u_cpu.ALU.u_wallace._1848_ ),
    .Y(\u_cpu.ALU.u_wallace._2552_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._8171_  (.A1(\u_cpu.ALU.u_wallace._4813_ ),
    .A2(\u_cpu.ALU.u_wallace._2053_ ),
    .B1(\u_cpu.ALU.u_wallace._2551_ ),
    .B2(\u_cpu.ALU.u_wallace._2552_ ),
    .X(\u_cpu.ALU.u_wallace._2553_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8172_  (.A(\u_cpu.ALU.u_wallace._2550_ ),
    .B(\u_cpu.ALU.u_wallace._2553_ ),
    .Y(\u_cpu.ALU.u_wallace._2554_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8173_  (.A1(\u_cpu.ALU.u_wallace._2511_ ),
    .A2(\u_cpu.ALU.u_wallace._2554_ ),
    .B1(\u_cpu.ALU.u_wallace._2517_ ),
    .Y(\u_cpu.ALU.u_wallace._2555_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._8174_  (.A(\u_cpu.ALU.u_wallace._2513_ ),
    .Y(\u_cpu.ALU.u_wallace._2556_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._8175_  (.A1(\u_cpu.ALU.u_wallace._2555_ ),
    .A2(\u_cpu.ALU.u_wallace._2556_ ),
    .B1(\u_cpu.ALU.u_wallace._2518_ ),
    .C1(\u_cpu.ALU.u_wallace._2541_ ),
    .D1(\u_cpu.ALU.u_wallace._2547_ ),
    .X(\u_cpu.ALU.u_wallace._2557_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8176_  (.A1(\u_cpu.ALU.u_wallace._2206_ ),
    .A2(\u_cpu.ALU.u_wallace._2170_ ),
    .B1(\u_cpu.ALU.u_wallace._2212_ ),
    .Y(\u_cpu.ALU.u_wallace._2558_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8177_  (.A1(\u_cpu.ALU.u_wallace._2548_ ),
    .A2(\u_cpu.ALU.u_wallace._2557_ ),
    .B1(\u_cpu.ALU.u_wallace._2558_ ),
    .Y(\u_cpu.ALU.u_wallace._2559_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8178_  (.A(\u_cpu.ALU.u_wallace._2356_ ),
    .B(\u_cpu.ALU.u_wallace._2368_ ),
    .Y(\u_cpu.ALU.u_wallace._2561_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8179_  (.A(\u_cpu.ALU.u_wallace._2559_ ),
    .B(\u_cpu.ALU.u_wallace._2561_ ),
    .Y(\u_cpu.ALU.u_wallace._2562_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._8180_  (.A1(\u_cpu.ALU.u_wallace._2211_ ),
    .A2(\u_cpu.ALU.u_wallace._2205_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2170_ ),
    .Y(\u_cpu.ALU.u_wallace._2563_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8181_  (.A1(\u_cpu.ALU.u_wallace._2518_ ),
    .A2(\u_cpu.ALU.u_wallace._2519_ ),
    .B1(\u_cpu.ALU.u_wallace._2541_ ),
    .B2(\u_cpu.ALU.u_wallace._2547_ ),
    .X(\u_cpu.ALU.u_wallace._2564_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._8182_  (.A1(\u_cpu.ALU.u_wallace._2555_ ),
    .A2(\u_cpu.ALU.u_wallace._2556_ ),
    .B1(\u_cpu.ALU.u_wallace._2518_ ),
    .C1(\u_cpu.ALU.u_wallace._2541_ ),
    .D1(\u_cpu.ALU.u_wallace._2547_ ),
    .Y(\u_cpu.ALU.u_wallace._2565_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8183_  (.A1(\u_cpu.ALU.u_wallace._2212_ ),
    .A2(\u_cpu.ALU.u_wallace._2563_ ),
    .B1(\u_cpu.ALU.u_wallace._2564_ ),
    .C1(\u_cpu.ALU.u_wallace._2565_ ),
    .X(\u_cpu.ALU.u_wallace._2566_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8184_  (.A1(\u_cpu.ALU.u_wallace._2225_ ),
    .A2(\u_cpu.ALU.u_wallace._2243_ ),
    .B1(\u_cpu.ALU.u_wallace._2245_ ),
    .Y(\u_cpu.ALU.u_wallace._2567_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._8185_  (.A1_N(\u_cpu.ALU.u_wallace._2262_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2267_ ),
    .B1(\u_cpu.ALU.u_wallace._2272_ ),
    .B2(\u_cpu.ALU.u_wallace._2567_ ),
    .Y(\u_cpu.ALU.u_wallace._2568_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8186_  (.A(\u_cpu.ALU.u_wallace._2226_ ),
    .X(\u_cpu.ALU.u_wallace._2569_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._8187_  (.A1(\u_cpu.ALU.u_wallace._0097_ ),
    .A2(\u_cpu.ALU.u_wallace._2569_ ),
    .A3(\u_cpu.ALU.u_wallace._2219_ ),
    .A4(\u_cpu.ALU.u_wallace._2221_ ),
    .B1(\u_cpu.ALU.u_wallace._2233_ ),
    .X(\u_cpu.ALU.u_wallace._2570_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8188_  (.A(\u_cpu.ALU.u_wallace._2270_ ),
    .B(\u_cpu.ALU.u_wallace._2241_ ),
    .Y(\u_cpu.ALU.u_wallace._2572_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8189_  (.A(\u_cpu.ALU.u_wallace._4431_ ),
    .B(\u_cpu.ALU.u_wallace._0802_ ),
    .Y(\u_cpu.ALU.u_wallace._2573_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8190_  (.A(\u_cpu.ALU.u_wallace._4450_ ),
    .B(\u_cpu.ALU.u_wallace._1102_ ),
    .Y(\u_cpu.ALU.u_wallace._2574_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8191_  (.A1(\u_cpu.ALU.u_wallace._2573_ ),
    .A2(\u_cpu.ALU.u_wallace._2574_ ),
    .B1(\u_cpu.ALU.u_wallace._2227_ ),
    .Y(\u_cpu.ALU.u_wallace._2575_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8192_  (.A1(\u_cpu.ALU.SrcA[8] ),
    .A2(\u_cpu.ALU.u_wallace._0628_ ),
    .B1(\u_cpu.ALU.SrcA[19] ),
    .B2(\u_cpu.ALU.u_wallace._1815_ ),
    .X(\u_cpu.ALU.u_wallace._2576_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8193_  (.A(\u_cpu.ALU.u_wallace._2768_ ),
    .B(\u_cpu.ALU.u_wallace._3645_ ),
    .C(\u_cpu.ALU.u_wallace._0626_ ),
    .D(\u_cpu.ALU.u_wallace._1100_ ),
    .Y(\u_cpu.ALU.u_wallace._2577_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8194_  (.A(\u_cpu.ALU.SrcA[25] ),
    .X(\u_cpu.ALU.u_wallace._2578_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8195_  (.A(\u_cpu.ALU.u_wallace._2576_ ),
    .B(\u_cpu.ALU.u_wallace._2577_ ),
    .C(\u_cpu.ALU.u_wallace._1859_ ),
    .D(\u_cpu.ALU.u_wallace._2578_ ),
    .Y(\u_cpu.ALU.u_wallace._2579_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._8196_  (.A(\u_cpu.ALU.SrcA[25] ),
    .Y(\u_cpu.ALU.u_wallace._2580_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8197_  (.A1(\u_cpu.ALU.u_wallace._3645_ ),
    .A2(\u_cpu.ALU.u_wallace._0626_ ),
    .B1(\u_cpu.ALU.u_wallace._1100_ ),
    .B2(\u_cpu.ALU.u_wallace._4649_ ),
    .Y(\u_cpu.ALU.u_wallace._2581_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8198_  (.A(\u_cpu.ALU.u_wallace._1815_ ),
    .B(\u_cpu.ALU.SrcA[8] ),
    .C(\u_cpu.ALU.u_wallace._0628_ ),
    .D(\u_cpu.ALU.SrcA[19] ),
    .X(\u_cpu.ALU.u_wallace._2583_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8199_  (.A1(\u_cpu.ALU.u_wallace._0634_ ),
    .A2(\u_cpu.ALU.u_wallace._2580_ ),
    .B1(\u_cpu.ALU.u_wallace._2581_ ),
    .B2(\u_cpu.ALU.u_wallace._2583_ ),
    .Y(\u_cpu.ALU.u_wallace._2584_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8200_  (.A1(\u_cpu.ALU.u_wallace._2217_ ),
    .A2(\u_cpu.ALU.u_wallace._2575_ ),
    .B1(\u_cpu.ALU.u_wallace._2579_ ),
    .C1(\u_cpu.ALU.u_wallace._2584_ ),
    .X(\u_cpu.ALU.u_wallace._2585_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8201_  (.A1(\u_cpu.ALU.u_wallace._2227_ ),
    .A2(\u_cpu.ALU.u_wallace._2216_ ),
    .B1(\u_cpu.ALU.u_wallace._2221_ ),
    .Y(\u_cpu.ALU.u_wallace._2586_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8202_  (.A1(\u_cpu.ALU.u_wallace._2584_ ),
    .A2(\u_cpu.ALU.u_wallace._2579_ ),
    .B1(\u_cpu.ALU.u_wallace._2586_ ),
    .Y(\u_cpu.ALU.u_wallace._2587_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8203_  (.A1(\u_cpu.ALU.u_wallace._1914_ ),
    .A2(\u_cpu.ALU.u_wallace._2000_ ),
    .B1(\u_cpu.ALU.u_wallace._2226_ ),
    .B2(\u_cpu.ALU.u_wallace._1903_ ),
    .Y(\u_cpu.ALU.u_wallace._2588_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8204_  (.A(\u_cpu.ALU.u_wallace._0742_ ),
    .B(\u_cpu.ALU.SrcA[22] ),
    .Y(\u_cpu.ALU.u_wallace._2589_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._8205_  (.A1(\u_cpu.ALU.u_wallace._0187_ ),
    .A2(\u_cpu.ALU.u_wallace._0304_ ),
    .A3(\u_cpu.ALU.u_wallace._2000_ ),
    .A4(\u_cpu.ALU.u_wallace._2222_ ),
    .B1(\u_cpu.ALU.u_wallace._2589_ ),
    .X(\u_cpu.ALU.u_wallace._2590_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8206_  (.A(\u_cpu.ALU.u_wallace._1903_ ),
    .B(\u_cpu.ALU.u_wallace._0807_ ),
    .C(\u_cpu.ALU.SrcA[23] ),
    .D(\u_cpu.ALU.u_wallace._2226_ ),
    .X(\u_cpu.ALU.u_wallace._2591_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8207_  (.A1(\u_cpu.ALU.u_wallace._2588_ ),
    .A2(\u_cpu.ALU.u_wallace._2591_ ),
    .B1(\u_cpu.ALU.u_wallace._2589_ ),
    .Y(\u_cpu.ALU.u_wallace._2592_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._8208_  (.A1(\u_cpu.ALU.u_wallace._2588_ ),
    .A2(\u_cpu.ALU.u_wallace._2590_ ),
    .B1(\u_cpu.ALU.u_wallace._2592_ ),
    .X(\u_cpu.ALU.u_wallace._2594_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8209_  (.A1(\u_cpu.ALU.u_wallace._2585_ ),
    .A2(\u_cpu.ALU.u_wallace._2587_ ),
    .B1(\u_cpu.ALU.u_wallace._2594_ ),
    .Y(\u_cpu.ALU.u_wallace._2595_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._8210_  (.A1(\u_cpu.ALU.u_wallace._1892_ ),
    .A2(\u_cpu.ALU.u_wallace._1737_ ),
    .B1(\u_cpu.ALU.u_wallace._2588_ ),
    .B2(\u_cpu.ALU.u_wallace._2591_ ),
    .X(\u_cpu.ALU.u_wallace._2596_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8211_  (.A(\u_cpu.ALU.u_wallace._0187_ ),
    .B(\u_cpu.ALU.u_wallace._1169_ ),
    .C(\u_cpu.ALU.u_wallace._2000_ ),
    .D(\u_cpu.ALU.u_wallace._2226_ ),
    .Y(\u_cpu.ALU.u_wallace._2597_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8212_  (.A(\u_cpu.ALU.u_wallace._1734_ ),
    .X(\u_cpu.ALU.u_wallace._2598_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.ALU.u_wallace._8213_  (.A_N(\u_cpu.ALU.u_wallace._2588_ ),
    .B(\u_cpu.ALU.u_wallace._2597_ ),
    .C(\u_cpu.ALU.u_wallace._0578_ ),
    .D(\u_cpu.ALU.u_wallace._2598_ ),
    .X(\u_cpu.ALU.u_wallace._2599_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8214_  (.A1(\u_cpu.ALU.u_wallace._2217_ ),
    .A2(\u_cpu.ALU.u_wallace._2575_ ),
    .B1(\u_cpu.ALU.u_wallace._2579_ ),
    .C1(\u_cpu.ALU.u_wallace._2584_ ),
    .Y(\u_cpu.ALU.u_wallace._2600_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8215_  (.A1(\u_cpu.ALU.u_wallace._0086_ ),
    .A2(\u_cpu.ALU.u_wallace._2578_ ),
    .B1(\u_cpu.ALU.u_wallace._2576_ ),
    .B2(\u_cpu.ALU.u_wallace._2577_ ),
    .Y(\u_cpu.ALU.u_wallace._2601_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8216_  (.A(\u_cpu.ALU.u_wallace._1749_ ),
    .B(\u_cpu.ALU.u_wallace._2578_ ),
    .Y(\u_cpu.ALU.u_wallace._2602_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._8217_  (.A(\u_cpu.ALU.u_wallace._2602_ ),
    .B(\u_cpu.ALU.u_wallace._2581_ ),
    .C(\u_cpu.ALU.u_wallace._2583_ ),
    .Y(\u_cpu.ALU.u_wallace._2603_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._8218_  (.A1(\u_cpu.ALU.u_wallace._4923_ ),
    .A2(\u_cpu.ALU.u_wallace._2215_ ),
    .A3(\u_cpu.ALU.u_wallace._2216_ ),
    .B1(\u_cpu.ALU.u_wallace._2221_ ),
    .X(\u_cpu.ALU.u_wallace._2605_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8219_  (.A1(\u_cpu.ALU.u_wallace._2601_ ),
    .A2(\u_cpu.ALU.u_wallace._2603_ ),
    .B1(\u_cpu.ALU.u_wallace._2605_ ),
    .Y(\u_cpu.ALU.u_wallace._2606_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8220_  (.A1(\u_cpu.ALU.u_wallace._2596_ ),
    .A2(\u_cpu.ALU.u_wallace._2599_ ),
    .B1(\u_cpu.ALU.u_wallace._2600_ ),
    .C1(\u_cpu.ALU.u_wallace._2606_ ),
    .Y(\u_cpu.ALU.u_wallace._2607_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8221_  (.A1(\u_cpu.ALU.u_wallace._2570_ ),
    .A2(\u_cpu.ALU.u_wallace._2572_ ),
    .B1(\u_cpu.ALU.u_wallace._2595_ ),
    .B2(\u_cpu.ALU.u_wallace._2607_ ),
    .Y(\u_cpu.ALU.u_wallace._2608_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8222_  (.A(\u_cpu.ALU.u_wallace._2238_ ),
    .B(\u_cpu.ALU.u_wallace._2237_ ),
    .Y(\u_cpu.ALU.u_wallace._2609_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8223_  (.A1(\u_cpu.ALU.u_wallace._1552_ ),
    .A2(\u_cpu.ALU.u_wallace._1543_ ),
    .B1(\u_cpu.ALU.u_wallace._1535_ ),
    .B2(\u_cpu.ALU.u_wallace._1530_ ),
    .X(\u_cpu.ALU.u_wallace._2610_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8224_  (.A(\u_cpu.ALU.u_wallace._2155_ ),
    .B(\u_cpu.ALU.u_wallace._2187_ ),
    .C(\u_cpu.ALU.u_wallace._1543_ ),
    .D(\u_cpu.ALU.u_wallace._1531_ ),
    .Y(\u_cpu.ALU.u_wallace._2611_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8225_  (.A(\u_cpu.ALU.u_wallace._2610_ ),
    .B(\u_cpu.ALU.u_wallace._2611_ ),
    .C(\u_cpu.ALU.u_wallace._2604_ ),
    .D(\u_cpu.ALU.u_wallace._0815_ ),
    .Y(\u_cpu.ALU.u_wallace._2612_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8226_  (.A1(\u_cpu.ALU.u_wallace._2187_ ),
    .A2(\u_cpu.ALU.u_wallace._1543_ ),
    .B1(\u_cpu.ALU.u_wallace._1531_ ),
    .B2(\u_cpu.ALU.u_wallace._2155_ ),
    .Y(\u_cpu.ALU.u_wallace._2613_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8227_  (.A(\u_cpu.ALU.u_wallace._2045_ ),
    .B(\u_cpu.ALU.u_wallace._2582_ ),
    .C(\u_cpu.ALU.u_wallace._1543_ ),
    .D(\u_cpu.ALU.u_wallace._1730_ ),
    .X(\u_cpu.ALU.u_wallace._2614_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8228_  (.A1(\u_cpu.ALU.u_wallace._4539_ ),
    .A2(\u_cpu.ALU.u_wallace._0809_ ),
    .B1(\u_cpu.ALU.u_wallace._2613_ ),
    .B2(\u_cpu.ALU.u_wallace._2614_ ),
    .Y(\u_cpu.ALU.u_wallace._2616_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8229_  (.A1(\u_cpu.ALU.u_wallace._2239_ ),
    .A2(\u_cpu.ALU.u_wallace._2609_ ),
    .B1(\u_cpu.ALU.u_wallace._2612_ ),
    .C1(\u_cpu.ALU.u_wallace._2616_ ),
    .X(\u_cpu.ALU.u_wallace._2617_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8230_  (.A(\u_cpu.ALU.u_wallace._1535_ ),
    .X(\u_cpu.ALU.u_wallace._2618_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8231_  (.A1(\u_cpu.ALU.u_wallace._2234_ ),
    .A2(\u_cpu.ALU.u_wallace._2618_ ),
    .A3(\u_cpu.ALU.u_wallace._0983_ ),
    .B1(\u_cpu.ALU.u_wallace._2239_ ),
    .X(\u_cpu.ALU.u_wallace._2619_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8232_  (.A1(\u_cpu.ALU.u_wallace._2612_ ),
    .A2(\u_cpu.ALU.u_wallace._2616_ ),
    .B1(\u_cpu.ALU.u_wallace._2619_ ),
    .Y(\u_cpu.ALU.u_wallace._2620_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8233_  (.A(\u_cpu.ALU.u_wallace._1286_ ),
    .X(\u_cpu.ALU.u_wallace._2621_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8234_  (.A1(\u_cpu.ALU.u_wallace._2252_ ),
    .A2(\u_cpu.ALU.u_wallace._2621_ ),
    .A3(\u_cpu.ALU.u_wallace._0015_ ),
    .B1(\u_cpu.ALU.u_wallace._2257_ ),
    .X(\u_cpu.ALU.u_wallace._2622_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._8235_  (.A1(\u_cpu.ALU.u_wallace._2617_ ),
    .A2(\u_cpu.ALU.u_wallace._2620_ ),
    .B1(\u_cpu.ALU.u_wallace._2622_ ),
    .X(\u_cpu.ALU.u_wallace._2623_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8236_  (.A1(\u_cpu.ALU.u_wallace._2612_ ),
    .A2(\u_cpu.ALU.u_wallace._2616_ ),
    .B1(\u_cpu.ALU.u_wallace._2619_ ),
    .X(\u_cpu.ALU.u_wallace._2624_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._8237_  (.A1(\u_cpu.ALU.u_wallace._2284_ ),
    .A2(\u_cpu.ALU.u_wallace._0635_ ),
    .A3(\u_cpu.ALU.u_wallace._2256_ ),
    .B1(\u_cpu.ALU.u_wallace._2254_ ),
    .X(\u_cpu.ALU.u_wallace._2625_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8238_  (.A1(\u_cpu.ALU.u_wallace._2239_ ),
    .A2(\u_cpu.ALU.u_wallace._2609_ ),
    .B1(\u_cpu.ALU.u_wallace._2612_ ),
    .C1(\u_cpu.ALU.u_wallace._2616_ ),
    .Y(\u_cpu.ALU.u_wallace._2627_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8239_  (.A(\u_cpu.ALU.u_wallace._2624_ ),
    .B(\u_cpu.ALU.u_wallace._2625_ ),
    .C(\u_cpu.ALU.u_wallace._2627_ ),
    .X(\u_cpu.ALU.u_wallace._2628_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._8240_  (.A1_N(\u_cpu.ALU.u_wallace._2228_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2233_ ),
    .B1(\u_cpu.ALU.u_wallace._2241_ ),
    .B2(\u_cpu.ALU.u_wallace._2270_ ),
    .Y(\u_cpu.ALU.u_wallace._2629_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8241_  (.A(\u_cpu.ALU.u_wallace._2595_ ),
    .B(\u_cpu.ALU.u_wallace._2607_ ),
    .C(\u_cpu.ALU.u_wallace._2629_ ),
    .Y(\u_cpu.ALU.u_wallace._2630_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8242_  (.A1(\u_cpu.ALU.u_wallace._2623_ ),
    .A2(\u_cpu.ALU.u_wallace._2628_ ),
    .B1(\u_cpu.ALU.u_wallace._2630_ ),
    .Y(\u_cpu.ALU.u_wallace._2631_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8243_  (.A(\u_cpu.ALU.u_wallace._2622_ ),
    .B(\u_cpu.ALU.u_wallace._2627_ ),
    .C(\u_cpu.ALU.u_wallace._2624_ ),
    .X(\u_cpu.ALU.u_wallace._2632_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._8244_  (.A1(\u_cpu.ALU.u_wallace._2617_ ),
    .A2(\u_cpu.ALU.u_wallace._2620_ ),
    .B1(\u_cpu.ALU.u_wallace._2625_ ),
    .X(\u_cpu.ALU.u_wallace._2633_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._8245_  (.A1(\u_cpu.ALU.u_wallace._2590_ ),
    .A2(\u_cpu.ALU.u_wallace._2588_ ),
    .B1(\u_cpu.ALU.u_wallace._2592_ ),
    .C1(\u_cpu.ALU.u_wallace._2600_ ),
    .D1(\u_cpu.ALU.u_wallace._2606_ ),
    .Y(\u_cpu.ALU.u_wallace._2634_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8246_  (.A1(\u_cpu.ALU.u_wallace._2596_ ),
    .A2(\u_cpu.ALU.u_wallace._2599_ ),
    .B1(\u_cpu.ALU.u_wallace._2585_ ),
    .B2(\u_cpu.ALU.u_wallace._2587_ ),
    .Y(\u_cpu.ALU.u_wallace._2635_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8247_  (.A1_N(\u_cpu.ALU.u_wallace._2241_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2270_ ),
    .B1(\u_cpu.ALU.u_wallace._2233_ ),
    .B2(\u_cpu.ALU.u_wallace._2228_ ),
    .Y(\u_cpu.ALU.u_wallace._2636_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8248_  (.A1(\u_cpu.ALU.u_wallace._2634_ ),
    .A2(\u_cpu.ALU.u_wallace._2635_ ),
    .B1(\u_cpu.ALU.u_wallace._2636_ ),
    .Y(\u_cpu.ALU.u_wallace._2638_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8249_  (.A1(\u_cpu.ALU.u_wallace._2632_ ),
    .A2(\u_cpu.ALU.u_wallace._2633_ ),
    .B1(\u_cpu.ALU.u_wallace._2608_ ),
    .B2(\u_cpu.ALU.u_wallace._2638_ ),
    .Y(\u_cpu.ALU.u_wallace._2639_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._8250_  (.A1(\u_cpu.ALU.u_wallace._2247_ ),
    .A2(\u_cpu.ALU.u_wallace._2568_ ),
    .B1(\u_cpu.ALU.u_wallace._2608_ ),
    .B2(\u_cpu.ALU.u_wallace._2631_ ),
    .C1(\u_cpu.ALU.u_wallace._2639_ ),
    .X(\u_cpu.ALU.u_wallace._2640_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._8251_  (.A(\u_cpu.ALU.u_wallace._2196_ ),
    .Y(\u_cpu.ALU.u_wallace._2641_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8252_  (.A1(\u_cpu.ALU.u_wallace._1129_ ),
    .A2(\u_cpu.ALU.u_wallace._0117_ ),
    .B1(\u_cpu.ALU.u_wallace._2183_ ),
    .B2(\u_cpu.ALU.u_wallace._2184_ ),
    .X(\u_cpu.ALU.u_wallace._2642_ ));
 sky130_fd_sc_hd__or4_2 \u_cpu.ALU.u_wallace._8253_  (.A(\u_cpu.ALU.u_wallace._0169_ ),
    .B(\u_cpu.ALU.u_wallace._2199_ ),
    .C(\u_cpu.ALU.u_wallace._0124_ ),
    .D(\u_cpu.ALU.u_wallace._2197_ ),
    .X(\u_cpu.ALU.u_wallace._2643_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8254_  (.A(\u_cpu.ALU.u_wallace._2190_ ),
    .B(\u_cpu.ALU.u_wallace._2642_ ),
    .C(\u_cpu.ALU.u_wallace._2643_ ),
    .X(\u_cpu.ALU.u_wallace._2644_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8255_  (.A(\u_cpu.ALU.u_wallace._2180_ ),
    .B(\u_cpu.ALU.u_wallace._2179_ ),
    .Y(\u_cpu.ALU.u_wallace._2645_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8256_  (.A(\u_cpu.ALU.u_wallace._4847_ ),
    .B(\u_cpu.ALU.u_wallace._4598_ ),
    .C(\u_cpu.ALU.u_wallace._0441_ ),
    .D(\u_cpu.ALU.u_wallace._0630_ ),
    .X(\u_cpu.ALU.u_wallace._2646_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8257_  (.A1(\u_cpu.ALU.u_wallace._4848_ ),
    .A2(\u_cpu.ALU.u_wallace._0448_ ),
    .B1(\u_cpu.ALU.u_wallace._0642_ ),
    .B2(\u_cpu.ALU.u_wallace._4720_ ),
    .Y(\u_cpu.ALU.u_wallace._2647_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8258_  (.A1(\u_cpu.ALU.u_wallace._4602_ ),
    .A2(\u_cpu.ALU.u_wallace._1324_ ),
    .B1(\u_cpu.ALU.u_wallace._2646_ ),
    .B2(\u_cpu.ALU.u_wallace._2647_ ),
    .Y(\u_cpu.ALU.u_wallace._2649_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8259_  (.A1(\u_cpu.ALU.u_wallace._4848_ ),
    .A2(\u_cpu.ALU.u_wallace._0448_ ),
    .B1(\u_cpu.ALU.u_wallace._0642_ ),
    .B2(\u_cpu.ALU.u_wallace._4720_ ),
    .X(\u_cpu.ALU.u_wallace._2650_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8260_  (.A(\u_cpu.ALU.u_wallace._4018_ ),
    .B(\u_cpu.ALU.u_wallace._4595_ ),
    .C(\u_cpu.ALU.u_wallace._0850_ ),
    .D(\u_cpu.ALU.u_wallace._0642_ ),
    .Y(\u_cpu.ALU.u_wallace._2651_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8261_  (.A(\u_cpu.ALU.u_wallace._2650_ ),
    .B(\u_cpu.ALU.u_wallace._0826_ ),
    .C(\u_cpu.ALU.u_wallace._0052_ ),
    .D(\u_cpu.ALU.u_wallace._2651_ ),
    .Y(\u_cpu.ALU.u_wallace._2652_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8262_  (.A1(\u_cpu.ALU.u_wallace._2181_ ),
    .A2(\u_cpu.ALU.u_wallace._2645_ ),
    .B1(\u_cpu.ALU.u_wallace._2649_ ),
    .C1(\u_cpu.ALU.u_wallace._2652_ ),
    .X(\u_cpu.ALU.u_wallace._2653_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._8263_  (.A1(\u_cpu.ALU.u_wallace._4602_ ),
    .A2(\u_cpu.ALU.u_wallace._1323_ ),
    .A3(\u_cpu.ALU.u_wallace._2179_ ),
    .B1(\u_cpu.ALU.u_wallace._2175_ ),
    .X(\u_cpu.ALU.u_wallace._2654_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8264_  (.A(\u_cpu.ALU.u_wallace._2649_ ),
    .B(\u_cpu.ALU.u_wallace._2652_ ),
    .Y(\u_cpu.ALU.u_wallace._2655_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8265_  (.A1(\u_cpu.ALU.u_wallace._0144_ ),
    .A2(\u_cpu.ALU.u_wallace._4921_ ),
    .B1(\u_cpu.ALU.u_wallace._0179_ ),
    .B2(\u_cpu.ALU.u_wallace._0028_ ),
    .Y(\u_cpu.ALU.u_wallace._2656_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8266_  (.A(\u_cpu.ALU.u_wallace._4837_ ),
    .B(\u_cpu.ALU.u_wallace._0029_ ),
    .C(\u_cpu.ALU.u_wallace._0188_ ),
    .D(\u_cpu.ALU.u_wallace._0179_ ),
    .X(\u_cpu.ALU.u_wallace._2657_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8267_  (.A(\u_cpu.ALU.u_wallace._0475_ ),
    .X(\u_cpu.ALU.u_wallace._2658_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8268_  (.A1(\u_cpu.ALU.u_wallace._2656_ ),
    .A2(\u_cpu.ALU.u_wallace._2657_ ),
    .B1(\u_cpu.ALU.u_wallace._2658_ ),
    .C1(\u_cpu.ALU.u_wallace._0034_ ),
    .X(\u_cpu.ALU.u_wallace._2660_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU.u_wallace._8269_  (.A1(\u_cpu.ALU.u_wallace._2658_ ),
    .A2(\u_cpu.ALU.u_wallace._0034_ ),
    .B1(\u_cpu.ALU.u_wallace._2656_ ),
    .C1(\u_cpu.ALU.u_wallace._2657_ ),
    .Y(\u_cpu.ALU.u_wallace._2661_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8270_  (.A1_N(\u_cpu.ALU.u_wallace._2654_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2655_ ),
    .B1(\u_cpu.ALU.u_wallace._2660_ ),
    .B2(\u_cpu.ALU.u_wallace._2661_ ),
    .Y(\u_cpu.ALU.u_wallace._2662_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8271_  (.A(\u_cpu.ALU.u_wallace._2285_ ),
    .B(\u_cpu.ALU.u_wallace._2266_ ),
    .Y(\u_cpu.ALU.u_wallace._2663_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._8272_  (.A1(\u_cpu.ALU.u_wallace._4913_ ),
    .A2(\u_cpu.ALU.u_wallace._0124_ ),
    .B1(\u_cpu.ALU.u_wallace._2656_ ),
    .B2(\u_cpu.ALU.u_wallace._2657_ ),
    .X(\u_cpu.ALU.u_wallace._2664_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8273_  (.A(\u_cpu.ALU.u_wallace._4840_ ),
    .B(\u_cpu.ALU.u_wallace._4842_ ),
    .C(\u_cpu.ALU.u_wallace._0319_ ),
    .D(\u_cpu.ALU.u_wallace._0320_ ),
    .Y(\u_cpu.ALU.u_wallace._2665_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.ALU.u_wallace._8274_  (.A_N(\u_cpu.ALU.u_wallace._2656_ ),
    .B(\u_cpu.ALU.u_wallace._2665_ ),
    .C(\u_cpu.ALU.u_wallace._2658_ ),
    .D(\u_cpu.ALU.u_wallace._0034_ ),
    .X(\u_cpu.ALU.u_wallace._2666_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8275_  (.A1(\u_cpu.ALU.u_wallace._2177_ ),
    .A2(\u_cpu.ALU.u_wallace._0652_ ),
    .A3(\u_cpu.ALU.u_wallace._0052_ ),
    .B1(\u_cpu.ALU.u_wallace._2181_ ),
    .X(\u_cpu.ALU.u_wallace._2667_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8276_  (.A1(\u_cpu.ALU.u_wallace._2649_ ),
    .A2(\u_cpu.ALU.u_wallace._2652_ ),
    .B1(\u_cpu.ALU.u_wallace._2667_ ),
    .Y(\u_cpu.ALU.u_wallace._2668_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8277_  (.A1(\u_cpu.ALU.u_wallace._2664_ ),
    .A2(\u_cpu.ALU.u_wallace._2666_ ),
    .B1(\u_cpu.ALU.u_wallace._2653_ ),
    .B2(\u_cpu.ALU.u_wallace._2668_ ),
    .Y(\u_cpu.ALU.u_wallace._2669_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._8278_  (.A1(\u_cpu.ALU.u_wallace._2653_ ),
    .A2(\u_cpu.ALU.u_wallace._2662_ ),
    .B1(\u_cpu.ALU.u_wallace._2282_ ),
    .B2(\u_cpu.ALU.u_wallace._2663_ ),
    .C1(\u_cpu.ALU.u_wallace._2669_ ),
    .Y(\u_cpu.ALU.u_wallace._2671_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8279_  (.A1(\u_cpu.ALU.u_wallace._2660_ ),
    .A2(\u_cpu.ALU.u_wallace._2661_ ),
    .B1(\u_cpu.ALU.u_wallace._2653_ ),
    .B2(\u_cpu.ALU.u_wallace._2668_ ),
    .Y(\u_cpu.ALU.u_wallace._2672_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8280_  (.A1(\u_cpu.ALU.u_wallace._2181_ ),
    .A2(\u_cpu.ALU.u_wallace._2645_ ),
    .B1(\u_cpu.ALU.u_wallace._2649_ ),
    .C1(\u_cpu.ALU.u_wallace._2652_ ),
    .Y(\u_cpu.ALU.u_wallace._2673_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8281_  (.A1(\u_cpu.ALU.u_wallace._2649_ ),
    .A2(\u_cpu.ALU.u_wallace._2652_ ),
    .B1(\u_cpu.ALU.u_wallace._2667_ ),
    .X(\u_cpu.ALU.u_wallace._2674_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8282_  (.A1(\u_cpu.ALU.u_wallace._2664_ ),
    .A2(\u_cpu.ALU.u_wallace._2666_ ),
    .B1(\u_cpu.ALU.u_wallace._2673_ ),
    .C1(\u_cpu.ALU.u_wallace._2674_ ),
    .Y(\u_cpu.ALU.u_wallace._2675_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8283_  (.A1(\u_cpu.ALU.u_wallace._2255_ ),
    .A2(\u_cpu.ALU.u_wallace._2263_ ),
    .B1(\u_cpu.ALU.u_wallace._2261_ ),
    .B2(\u_cpu.ALU.u_wallace._2265_ ),
    .Y(\u_cpu.ALU.u_wallace._2676_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8284_  (.A(\u_cpu.ALU.u_wallace._2672_ ),
    .B(\u_cpu.ALU.u_wallace._2675_ ),
    .C(\u_cpu.ALU.u_wallace._2676_ ),
    .Y(\u_cpu.ALU.u_wallace._2677_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._8285_  (.A1_N(\u_cpu.ALU.u_wallace._2641_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2644_ ),
    .B1(\u_cpu.ALU.u_wallace._2671_ ),
    .B2(\u_cpu.ALU.u_wallace._2677_ ),
    .Y(\u_cpu.ALU.u_wallace._2678_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU.u_wallace._8286_  (.A(\u_cpu.ALU.u_wallace._2200_ ),
    .B(\u_cpu.ALU.u_wallace._2201_ ),
    .X(\u_cpu.ALU.u_wallace._2679_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._8287_  (.A1(\u_cpu.ALU.u_wallace._2679_ ),
    .A2(\u_cpu.ALU.u_wallace._2208_ ),
    .B1(\u_cpu.ALU.u_wallace._2196_ ),
    .C1(\u_cpu.ALU.u_wallace._2677_ ),
    .D1(\u_cpu.ALU.u_wallace._2671_ ),
    .X(\u_cpu.ALU.u_wallace._2680_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8288_  (.A1(\u_cpu.ALU.u_wallace._2617_ ),
    .A2(\u_cpu.ALU.u_wallace._2620_ ),
    .B1(\u_cpu.ALU.u_wallace._2622_ ),
    .Y(\u_cpu.ALU.u_wallace._2682_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8289_  (.A(\u_cpu.ALU.u_wallace._2624_ ),
    .B(\u_cpu.ALU.u_wallace._2625_ ),
    .C(\u_cpu.ALU.u_wallace._2627_ ),
    .Y(\u_cpu.ALU.u_wallace._2683_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8290_  (.A(\u_cpu.ALU.u_wallace._2636_ ),
    .B(\u_cpu.ALU.u_wallace._2634_ ),
    .C(\u_cpu.ALU.u_wallace._2635_ ),
    .Y(\u_cpu.ALU.u_wallace._2684_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8291_  (.A1(\u_cpu.ALU.u_wallace._2682_ ),
    .A2(\u_cpu.ALU.u_wallace._2683_ ),
    .B1(\u_cpu.ALU.u_wallace._2684_ ),
    .B2(\u_cpu.ALU.u_wallace._2630_ ),
    .X(\u_cpu.ALU.u_wallace._2685_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8292_  (.A(\u_cpu.ALU.u_wallace._2682_ ),
    .B(\u_cpu.ALU.u_wallace._2683_ ),
    .C(\u_cpu.ALU.u_wallace._2684_ ),
    .D(\u_cpu.ALU.u_wallace._2630_ ),
    .Y(\u_cpu.ALU.u_wallace._2686_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8293_  (.A1(\u_cpu.ALU.u_wallace._2273_ ),
    .A2(\u_cpu.ALU.u_wallace._2288_ ),
    .B1(\u_cpu.ALU.u_wallace._2247_ ),
    .Y(\u_cpu.ALU.u_wallace._2687_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8294_  (.A(\u_cpu.ALU.u_wallace._2685_ ),
    .B(\u_cpu.ALU.u_wallace._2686_ ),
    .C(\u_cpu.ALU.u_wallace._2687_ ),
    .Y(\u_cpu.ALU.u_wallace._2688_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8295_  (.A1(\u_cpu.ALU.u_wallace._2678_ ),
    .A2(\u_cpu.ALU.u_wallace._2680_ ),
    .B1(\u_cpu.ALU.u_wallace._2688_ ),
    .Y(\u_cpu.ALU.u_wallace._2689_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8296_  (.A1(\u_cpu.ALU.u_wallace._2623_ ),
    .A2(\u_cpu.ALU.u_wallace._2628_ ),
    .B1(\u_cpu.ALU.u_wallace._2684_ ),
    .C1(\u_cpu.ALU.u_wallace._2630_ ),
    .Y(\u_cpu.ALU.u_wallace._2690_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8297_  (.A1(\u_cpu.ALU.u_wallace._2247_ ),
    .A2(\u_cpu.ALU.u_wallace._2568_ ),
    .B1(\u_cpu.ALU.u_wallace._2690_ ),
    .C1(\u_cpu.ALU.u_wallace._2639_ ),
    .Y(\u_cpu.ALU.u_wallace._2691_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8298_  (.A1(\u_cpu.ALU.u_wallace._2190_ ),
    .A2(\u_cpu.ALU.u_wallace._2642_ ),
    .A3(\u_cpu.ALU.u_wallace._2643_ ),
    .B1(\u_cpu.ALU.u_wallace._2641_ ),
    .X(\u_cpu.ALU.u_wallace._2693_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8299_  (.A(\u_cpu.ALU.u_wallace._2693_ ),
    .B(\u_cpu.ALU.u_wallace._2671_ ),
    .C(\u_cpu.ALU.u_wallace._2677_ ),
    .X(\u_cpu.ALU.u_wallace._2694_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8300_  (.A1(\u_cpu.ALU.u_wallace._2671_ ),
    .A2(\u_cpu.ALU.u_wallace._2677_ ),
    .B1(\u_cpu.ALU.u_wallace._2693_ ),
    .Y(\u_cpu.ALU.u_wallace._2695_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8301_  (.A1_N(\u_cpu.ALU.u_wallace._2691_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2688_ ),
    .B1(\u_cpu.ALU.u_wallace._2694_ ),
    .B2(\u_cpu.ALU.u_wallace._2695_ ),
    .Y(\u_cpu.ALU.u_wallace._2696_ ));
 sky130_fd_sc_hd__o32ai_2 \u_cpu.ALU.u_wallace._8302_  (.A1(\u_cpu.ALU.u_wallace._2290_ ),
    .A2(\u_cpu.ALU.u_wallace._2281_ ),
    .A3(\u_cpu.ALU.u_wallace._2289_ ),
    .B1(\u_cpu.ALU.u_wallace._2214_ ),
    .B2(\u_cpu.ALU.u_wallace._2299_ ),
    .Y(\u_cpu.ALU.u_wallace._2697_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8303_  (.A1(\u_cpu.ALU.u_wallace._2640_ ),
    .A2(\u_cpu.ALU.u_wallace._2689_ ),
    .B1(\u_cpu.ALU.u_wallace._2696_ ),
    .C1(\u_cpu.ALU.u_wallace._2697_ ),
    .Y(\u_cpu.ALU.u_wallace._2698_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8304_  (.A1(\u_cpu.ALU.u_wallace._2212_ ),
    .A2(\u_cpu.ALU.u_wallace._2563_ ),
    .B1(\u_cpu.ALU.u_wallace._2564_ ),
    .C1(\u_cpu.ALU.u_wallace._2565_ ),
    .Y(\u_cpu.ALU.u_wallace._2699_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8305_  (.A1(\u_cpu.ALU.u_wallace._2559_ ),
    .A2(\u_cpu.ALU.u_wallace._2699_ ),
    .B1(\u_cpu.ALU.u_wallace._2561_ ),
    .X(\u_cpu.ALU.u_wallace._2700_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8306_  (.A1(\u_cpu.ALU.u_wallace._2678_ ),
    .A2(\u_cpu.ALU.u_wallace._2680_ ),
    .B1(\u_cpu.ALU.u_wallace._2691_ ),
    .C1(\u_cpu.ALU.u_wallace._2688_ ),
    .X(\u_cpu.ALU.u_wallace._2701_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8307_  (.A1(\u_cpu.ALU.u_wallace._2641_ ),
    .A2(\u_cpu.ALU.u_wallace._2644_ ),
    .B1(\u_cpu.ALU.u_wallace._2677_ ),
    .Y(\u_cpu.ALU.u_wallace._2702_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8308_  (.A1(\u_cpu.ALU.u_wallace._2671_ ),
    .A2(\u_cpu.ALU.u_wallace._2677_ ),
    .A3(\u_cpu.ALU.u_wallace._2702_ ),
    .B1(\u_cpu.ALU.u_wallace._2678_ ),
    .X(\u_cpu.ALU.u_wallace._2704_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8309_  (.A1(\u_cpu.ALU.u_wallace._2691_ ),
    .A2(\u_cpu.ALU.u_wallace._2688_ ),
    .B1(\u_cpu.ALU.u_wallace._2704_ ),
    .Y(\u_cpu.ALU.u_wallace._2705_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._8310_  (.A1(\u_cpu.ALU.u_wallace._2701_ ),
    .A2(\u_cpu.ALU.u_wallace._2705_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2697_ ),
    .Y(\u_cpu.ALU.u_wallace._2706_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._8311_  (.A1(\u_cpu.ALU.u_wallace._2562_ ),
    .A2(\u_cpu.ALU.u_wallace._2566_ ),
    .B1(\u_cpu.ALU.u_wallace._2698_ ),
    .C1(\u_cpu.ALU.u_wallace._2700_ ),
    .D1(\u_cpu.ALU.u_wallace._2706_ ),
    .Y(\u_cpu.ALU.u_wallace._2707_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8312_  (.A1(\u_cpu.ALU.u_wallace._2559_ ),
    .A2(\u_cpu.ALU.u_wallace._2699_ ),
    .B1(\u_cpu.ALU.u_wallace._2561_ ),
    .Y(\u_cpu.ALU.u_wallace._2708_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8313_  (.A(\u_cpu.ALU.u_wallace._2559_ ),
    .B(\u_cpu.ALU.u_wallace._2699_ ),
    .C(\u_cpu.ALU.u_wallace._2561_ ),
    .X(\u_cpu.ALU.u_wallace._2709_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8314_  (.A1(\u_cpu.ALU.u_wallace._2678_ ),
    .A2(\u_cpu.ALU.u_wallace._2680_ ),
    .B1(\u_cpu.ALU.u_wallace._2691_ ),
    .C1(\u_cpu.ALU.u_wallace._2688_ ),
    .Y(\u_cpu.ALU.u_wallace._2710_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8315_  (.A1(\u_cpu.ALU.u_wallace._2710_ ),
    .A2(\u_cpu.ALU.u_wallace._2696_ ),
    .B1(\u_cpu.ALU.u_wallace._2697_ ),
    .Y(\u_cpu.ALU.u_wallace._2711_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8316_  (.A1(\u_cpu.ALU.u_wallace._2640_ ),
    .A2(\u_cpu.ALU.u_wallace._2689_ ),
    .B1(\u_cpu.ALU.u_wallace._2696_ ),
    .C1(\u_cpu.ALU.u_wallace._2697_ ),
    .X(\u_cpu.ALU.u_wallace._2712_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8317_  (.A1(\u_cpu.ALU.u_wallace._2708_ ),
    .A2(\u_cpu.ALU.u_wallace._2709_ ),
    .B1(\u_cpu.ALU.u_wallace._2711_ ),
    .B2(\u_cpu.ALU.u_wallace._2712_ ),
    .Y(\u_cpu.ALU.u_wallace._2713_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8318_  (.A(\u_cpu.ALU.u_wallace._2504_ ),
    .B(\u_cpu.ALU.u_wallace._2707_ ),
    .C(\u_cpu.ALU.u_wallace._2713_ ),
    .Y(\u_cpu.ALU.u_wallace._2715_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8319_  (.A(\u_cpu.ALU.u_wallace._2697_ ),
    .B(\u_cpu.ALU.u_wallace._2696_ ),
    .Y(\u_cpu.ALU.u_wallace._2716_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8320_  (.A(\u_cpu.ALU.u_wallace._2564_ ),
    .B(\u_cpu.ALU.u_wallace._2565_ ),
    .Y(\u_cpu.ALU.u_wallace._2717_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8321_  (.A1(\u_cpu.ALU.u_wallace._2356_ ),
    .A2(\u_cpu.ALU.u_wallace._2368_ ),
    .B1(\u_cpu.ALU.u_wallace._2717_ ),
    .B2(\u_cpu.ALU.u_wallace._2558_ ),
    .Y(\u_cpu.ALU.u_wallace._2718_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8322_  (.A1(\u_cpu.ALU.u_wallace._2699_ ),
    .A2(\u_cpu.ALU.u_wallace._2718_ ),
    .B1(\u_cpu.ALU.u_wallace._2708_ ),
    .Y(\u_cpu.ALU.u_wallace._2719_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8323_  (.A1(\u_cpu.ALU.u_wallace._2701_ ),
    .A2(\u_cpu.ALU.u_wallace._2716_ ),
    .B1(\u_cpu.ALU.u_wallace._2719_ ),
    .C1(\u_cpu.ALU.u_wallace._2706_ ),
    .X(\u_cpu.ALU.u_wallace._2720_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8324_  (.A1(\u_cpu.ALU.u_wallace._2558_ ),
    .A2(\u_cpu.ALU.u_wallace._2717_ ),
    .B1(\u_cpu.ALU.u_wallace._2718_ ),
    .Y(\u_cpu.ALU.u_wallace._2721_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8325_  (.A1(\u_cpu.ALU.u_wallace._2700_ ),
    .A2(\u_cpu.ALU.u_wallace._2721_ ),
    .B1(\u_cpu.ALU.u_wallace._2706_ ),
    .B2(\u_cpu.ALU.u_wallace._2698_ ),
    .Y(\u_cpu.ALU.u_wallace._2722_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._8326_  (.A1(\u_cpu.ALU.u_wallace._2720_ ),
    .A2(\u_cpu.ALU.u_wallace._2722_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2504_ ),
    .Y(\u_cpu.ALU.u_wallace._2723_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._8327_  (.A1(\u_cpu.ALU.u_wallace._2495_ ),
    .A2(\u_cpu.ALU.u_wallace._2497_ ),
    .B1(\u_cpu.ALU.u_wallace._2500_ ),
    .C1(\u_cpu.ALU.u_wallace._2715_ ),
    .D1(\u_cpu.ALU.u_wallace._2723_ ),
    .Y(\u_cpu.ALU.u_wallace._2724_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8328_  (.A1(\u_cpu.ALU.u_wallace._2498_ ),
    .A2(\u_cpu.ALU.u_wallace._2495_ ),
    .B1(\u_cpu.ALU.u_wallace._2395_ ),
    .C1(\u_cpu.ALU.u_wallace._2405_ ),
    .X(\u_cpu.ALU.u_wallace._2726_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8329_  (.A1(\u_cpu.ALU.u_wallace._2496_ ),
    .A2(\u_cpu.ALU.u_wallace._2493_ ),
    .B1(\u_cpu.ALU.u_wallace._2497_ ),
    .Y(\u_cpu.ALU.u_wallace._2727_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8330_  (.A1_N(\u_cpu.ALU.u_wallace._2715_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2723_ ),
    .B1(\u_cpu.ALU.u_wallace._2726_ ),
    .B2(\u_cpu.ALU.u_wallace._2727_ ),
    .Y(\u_cpu.ALU.u_wallace._2728_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8331_  (.A1(\u_cpu.ALU.u_wallace._2442_ ),
    .A2(\u_cpu.ALU.u_wallace._2414_ ),
    .B1(\u_cpu.ALU.u_wallace._2724_ ),
    .C1(\u_cpu.ALU.u_wallace._2728_ ),
    .Y(\u_cpu.ALU.u_wallace._2729_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8332_  (.A1(\u_cpu.ALU.u_wallace._2365_ ),
    .A2(\u_cpu.ALU.u_wallace._2369_ ),
    .B1(\u_cpu.ALU.u_wallace._2371_ ),
    .C1(\u_cpu.ALU.u_wallace._2384_ ),
    .Y(\u_cpu.ALU.u_wallace._2730_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8333_  (.A1(\u_cpu.ALU.u_wallace._2377_ ),
    .A2(\u_cpu.ALU.u_wallace._2730_ ),
    .B1(\u_cpu.ALU.u_wallace._2722_ ),
    .Y(\u_cpu.ALU.u_wallace._2731_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8334_  (.A1(\u_cpu.ALU.u_wallace._2495_ ),
    .A2(\u_cpu.ALU.u_wallace._2497_ ),
    .B1(\u_cpu.ALU.u_wallace._2500_ ),
    .Y(\u_cpu.ALU.u_wallace._2732_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8335_  (.A1(\u_cpu.ALU.u_wallace._2707_ ),
    .A2(\u_cpu.ALU.u_wallace._2713_ ),
    .B1(\u_cpu.ALU.u_wallace._2504_ ),
    .Y(\u_cpu.ALU.u_wallace._2733_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU.u_wallace._8336_  (.A1(\u_cpu.ALU.u_wallace._2731_ ),
    .A2(\u_cpu.ALU.u_wallace._2707_ ),
    .B1(\u_cpu.ALU.u_wallace._2732_ ),
    .C1(\u_cpu.ALU.u_wallace._2733_ ),
    .Y(\u_cpu.ALU.u_wallace._2734_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._8337_  (.A1(\u_cpu.ALU.u_wallace._2715_ ),
    .A2(\u_cpu.ALU.u_wallace._2723_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2732_ ),
    .Y(\u_cpu.ALU.u_wallace._2735_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8338_  (.A1(\u_cpu.ALU.u_wallace._2424_ ),
    .A2(\u_cpu.ALU.u_wallace._2430_ ),
    .B1(\u_cpu.ALU.u_wallace._2413_ ),
    .B2(\u_cpu.ALU.u_wallace._2441_ ),
    .Y(\u_cpu.ALU.u_wallace._2737_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._8339_  (.A1(\u_cpu.ALU.u_wallace._2734_ ),
    .A2(\u_cpu.ALU.u_wallace._2735_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2737_ ),
    .Y(\u_cpu.ALU.u_wallace._2738_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8340_  (.A1(\u_cpu.ALU.u_wallace._2412_ ),
    .A2(\u_cpu.ALU.u_wallace._2474_ ),
    .B1(\u_cpu.ALU.u_wallace._2729_ ),
    .C1(\u_cpu.ALU.u_wallace._2738_ ),
    .Y(\u_cpu.ALU.u_wallace._2739_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8341_  (.A1(\u_cpu.ALU.u_wallace._2442_ ),
    .A2(\u_cpu.ALU.u_wallace._2414_ ),
    .B1(\u_cpu.ALU.u_wallace._2724_ ),
    .C1(\u_cpu.ALU.u_wallace._2728_ ),
    .X(\u_cpu.ALU.u_wallace._2740_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8342_  (.A1(\u_cpu.ALU.u_wallace._2724_ ),
    .A2(\u_cpu.ALU.u_wallace._2728_ ),
    .B1(\u_cpu.ALU.u_wallace._2737_ ),
    .Y(\u_cpu.ALU.u_wallace._2741_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._8343_  (.A1(\u_cpu.ALU.u_wallace._1886_ ),
    .A2(\u_cpu.ALU.u_wallace._2409_ ),
    .A3(\u_cpu.ALU.u_wallace._2417_ ),
    .A4(\u_cpu.ALU.u_wallace._2135_ ),
    .B1(\u_cpu.ALU.u_wallace._2412_ ),
    .X(\u_cpu.ALU.u_wallace._2742_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._8344_  (.A(\u_cpu.ALU.u_wallace._2742_ ),
    .Y(\u_cpu.ALU.u_wallace._2743_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8345_  (.A1(\u_cpu.ALU.u_wallace._2740_ ),
    .A2(\u_cpu.ALU.u_wallace._2741_ ),
    .B1(\u_cpu.ALU.u_wallace._2743_ ),
    .Y(\u_cpu.ALU.u_wallace._2744_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8346_  (.A(\u_cpu.ALU.u_wallace._2473_ ),
    .B(\u_cpu.ALU.u_wallace._2739_ ),
    .C(\u_cpu.ALU.u_wallace._2744_ ),
    .Y(\u_cpu.ALU.u_wallace._2745_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8347_  (.A1(\u_cpu.ALU.u_wallace._2412_ ),
    .A2(\u_cpu.ALU.u_wallace._2474_ ),
    .B1(\u_cpu.ALU.u_wallace._2729_ ),
    .C1(\u_cpu.ALU.u_wallace._2738_ ),
    .X(\u_cpu.ALU.u_wallace._2746_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8348_  (.A1(\u_cpu.ALU.u_wallace._2729_ ),
    .A2(\u_cpu.ALU.u_wallace._2738_ ),
    .B1(\u_cpu.ALU.u_wallace._2742_ ),
    .Y(\u_cpu.ALU.u_wallace._2748_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._8349_  (.A1(\u_cpu.ALU.u_wallace._2746_ ),
    .A2(\u_cpu.ALU.u_wallace._2748_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2473_ ),
    .Y(\u_cpu.ALU.u_wallace._2749_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8350_  (.A1_N(\u_cpu.ALU.u_wallace._2745_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2749_ ),
    .B1(\u_cpu.ALU.u_wallace._2398_ ),
    .B2(\u_cpu.ALU.u_wallace._2399_ ),
    .Y(\u_cpu.ALU.u_wallace._2750_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._8351_  (.A_N(\u_cpu.ALU.u_wallace._2401_ ),
    .B(\u_cpu.ALU.u_wallace._2745_ ),
    .C(\u_cpu.ALU.u_wallace._2749_ ),
    .Y(\u_cpu.ALU.u_wallace._2751_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8352_  (.A1(\u_cpu.ALU.u_wallace._2750_ ),
    .A2(\u_cpu.ALU.u_wallace._2751_ ),
    .B1(\u_cpu.ALU.u_wallace._2449_ ),
    .X(\u_cpu.ALU.u_wallace._2752_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8353_  (.A1(\u_cpu.ALU.u_wallace._2446_ ),
    .A2(\u_cpu.ALU.u_wallace._2447_ ),
    .B1(\u_cpu.ALU.u_wallace._2751_ ),
    .C1(\u_cpu.ALU.u_wallace._2750_ ),
    .Y(\u_cpu.ALU.u_wallace._2753_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8354_  (.A(\u_cpu.ALU.u_wallace._2752_ ),
    .B(\u_cpu.ALU.u_wallace._2753_ ),
    .Y(\u_cpu.ALU.u_wallace._2754_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._8355_  (.A(\u_cpu.ALU.u_wallace._2470_ ),
    .B(\u_cpu.ALU.u_wallace._2754_ ),
    .X(\u_cpu.ALU.Product_Wallace[25] ));
 sky130_fd_sc_hd__or3_2 \u_cpu.ALU.u_wallace._8356_  (.A(\u_cpu.ALU.u_wallace._0414_ ),
    .B(\u_cpu.ALU.u_wallace._2131_ ),
    .C(\u_cpu.ALU.u_wallace._2487_ ),
    .X(\u_cpu.ALU.u_wallace._2755_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8357_  (.A1(\u_cpu.ALU.u_wallace._2743_ ),
    .A2(\u_cpu.ALU.u_wallace._2741_ ),
    .B1(\u_cpu.ALU.u_wallace._2729_ ),
    .Y(\u_cpu.ALU.u_wallace._2756_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._8358_  (.A1(\u_cpu.ALU.u_wallace._2653_ ),
    .A2(\u_cpu.ALU.u_wallace._2662_ ),
    .B1(\u_cpu.ALU.u_wallace._2282_ ),
    .B2(\u_cpu.ALU.u_wallace._2663_ ),
    .C1(\u_cpu.ALU.u_wallace._2669_ ),
    .X(\u_cpu.ALU.u_wallace._2758_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8359_  (.A1(\u_cpu.ALU.u_wallace._2693_ ),
    .A2(\u_cpu.ALU.u_wallace._2677_ ),
    .B1(\u_cpu.ALU.u_wallace._2758_ ),
    .Y(\u_cpu.ALU.u_wallace._2759_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8360_  (.A1(\u_cpu.ALU.u_wallace._4785_ ),
    .A2(\u_cpu.ALU.u_wallace._0730_ ),
    .B1(\u_cpu.ALU.u_wallace._0732_ ),
    .B2(\u_cpu.ALU.u_wallace._4647_ ),
    .X(\u_cpu.ALU.u_wallace._2760_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8361_  (.A(\u_cpu.ALU.u_wallace._4794_ ),
    .B(\u_cpu.ALU.u_wallace._4787_ ),
    .C(\u_cpu.ALU.u_wallace._0546_ ),
    .D(\u_cpu.ALU.u_wallace._0547_ ),
    .Y(\u_cpu.ALU.u_wallace._2761_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8362_  (.A(\u_cpu.ALU.u_wallace._2760_ ),
    .B(\u_cpu.ALU.u_wallace._0735_ ),
    .C(\u_cpu.ALU.u_wallace._4643_ ),
    .D(\u_cpu.ALU.u_wallace._2761_ ),
    .Y(\u_cpu.ALU.u_wallace._2762_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8363_  (.A1_N(\u_cpu.ALU.u_wallace._2761_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2760_ ),
    .B1(\u_cpu.ALU.u_wallace._4904_ ),
    .B2(\u_cpu.ALU.u_wallace._0941_ ),
    .Y(\u_cpu.ALU.u_wallace._2763_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8364_  (.A(\u_cpu.ALU.u_wallace._0475_ ),
    .B(\u_cpu.ALU.u_wallace._0033_ ),
    .Y(\u_cpu.ALU.u_wallace._2764_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8365_  (.A1(\u_cpu.ALU.u_wallace._2764_ ),
    .A2(\u_cpu.ALU.u_wallace._2656_ ),
    .B1(\u_cpu.ALU.u_wallace._2665_ ),
    .Y(\u_cpu.ALU.u_wallace._2765_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8366_  (.A1(\u_cpu.ALU.u_wallace._2762_ ),
    .A2(\u_cpu.ALU.u_wallace._2763_ ),
    .B1(\u_cpu.ALU.u_wallace._2765_ ),
    .Y(\u_cpu.ALU.u_wallace._2766_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8367_  (.A(\u_cpu.ALU.u_wallace._2762_ ),
    .B(\u_cpu.ALU.u_wallace._2763_ ),
    .C(\u_cpu.ALU.u_wallace._2765_ ),
    .X(\u_cpu.ALU.u_wallace._2767_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._8368_  (.A1(\u_cpu.ALU.u_wallace._4573_ ),
    .A2(\u_cpu.ALU.u_wallace._0554_ ),
    .A3(\u_cpu.ALU.u_wallace._2529_ ),
    .B1(\u_cpu.ALU.u_wallace._2526_ ),
    .X(\u_cpu.ALU.u_wallace._2769_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8369_  (.A1(\u_cpu.ALU.u_wallace._2766_ ),
    .A2(\u_cpu.ALU.u_wallace._2767_ ),
    .B1(\u_cpu.ALU.u_wallace._2769_ ),
    .Y(\u_cpu.ALU.u_wallace._2770_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8370_  (.A1(\u_cpu.ALU.u_wallace._2762_ ),
    .A2(\u_cpu.ALU.u_wallace._2763_ ),
    .B1(\u_cpu.ALU.u_wallace._2765_ ),
    .X(\u_cpu.ALU.u_wallace._2771_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8371_  (.A(\u_cpu.ALU.u_wallace._2762_ ),
    .B(\u_cpu.ALU.u_wallace._2763_ ),
    .C(\u_cpu.ALU.u_wallace._2765_ ),
    .Y(\u_cpu.ALU.u_wallace._2772_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._8372_  (.A_N(\u_cpu.ALU.u_wallace._2769_ ),
    .B(\u_cpu.ALU.u_wallace._2771_ ),
    .C(\u_cpu.ALU.u_wallace._2772_ ),
    .Y(\u_cpu.ALU.u_wallace._2773_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8373_  (.A1(\u_cpu.ALU.u_wallace._2537_ ),
    .A2(\u_cpu.ALU.u_wallace._2534_ ),
    .B1(\u_cpu.ALU.u_wallace._2539_ ),
    .Y(\u_cpu.ALU.u_wallace._2774_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8374_  (.A1(\u_cpu.ALU.u_wallace._2770_ ),
    .A2(\u_cpu.ALU.u_wallace._2773_ ),
    .B1(\u_cpu.ALU.u_wallace._2774_ ),
    .Y(\u_cpu.ALU.u_wallace._2775_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._8375_  (.A1(\u_cpu.ALU.u_wallace._2766_ ),
    .A2(\u_cpu.ALU.u_wallace._2767_ ),
    .B1(\u_cpu.ALU.u_wallace._2769_ ),
    .X(\u_cpu.ALU.u_wallace._2776_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8376_  (.A(\u_cpu.ALU.u_wallace._2537_ ),
    .B(\u_cpu.ALU.u_wallace._2534_ ),
    .Y(\u_cpu.ALU.u_wallace._2777_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8377_  (.A1(\u_cpu.ALU.u_wallace._2532_ ),
    .A2(\u_cpu.ALU.u_wallace._2777_ ),
    .B1(\u_cpu.ALU.u_wallace._2773_ ),
    .Y(\u_cpu.ALU.u_wallace._2778_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8378_  (.A(\u_cpu.ALU.u_wallace._4669_ ),
    .B(\u_cpu.ALU.u_wallace._2801_ ),
    .C(\u_cpu.ALU.u_wallace._2050_ ),
    .Y(\u_cpu.ALU.u_wallace._2780_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._8379_  (.A(\u_cpu.ALU.u_wallace._1848_ ),
    .B(\u_cpu.ALU.u_wallace._1386_ ),
    .X(\u_cpu.ALU.u_wallace._2781_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8380_  (.A1(\u_cpu.ALU.u_wallace._4449_ ),
    .A2(\u_cpu.ALU.u_wallace._1387_ ),
    .B1(\u_cpu.ALU.u_wallace._1210_ ),
    .B2(\u_cpu.ALU.u_wallace._2725_ ),
    .X(\u_cpu.ALU.u_wallace._2782_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8381_  (.A1(\u_cpu.ALU.u_wallace._1211_ ),
    .A2(\u_cpu.ALU.u_wallace._2780_ ),
    .B1(\u_cpu.ALU.u_wallace._2781_ ),
    .C1(\u_cpu.ALU.u_wallace._2782_ ),
    .X(\u_cpu.ALU.u_wallace._2783_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8382_  (.A(\u_cpu.ALU.u_wallace._4660_ ),
    .B(\u_cpu.ALU.u_wallace._3821_ ),
    .C(\u_cpu.ALU.u_wallace._2050_ ),
    .D(\u_cpu.ALU.u_wallace._1175_ ),
    .Y(\u_cpu.ALU.u_wallace._2784_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8383_  (.A1(\u_cpu.ALU.u_wallace._2784_ ),
    .A2(\u_cpu.ALU.u_wallace._2782_ ),
    .B1(\u_cpu.ALU.u_wallace._2781_ ),
    .Y(\u_cpu.ALU.u_wallace._2785_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8384_  (.A(\u_cpu.ALU.u_wallace._1322_ ),
    .B(\u_cpu.ALU.u_wallace._1386_ ),
    .Y(\u_cpu.ALU.u_wallace._2786_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8385_  (.A1(\u_cpu.ALU.u_wallace._2786_ ),
    .A2(\u_cpu.ALU.u_wallace._2552_ ),
    .B1(\u_cpu.ALU.u_wallace._2507_ ),
    .Y(\u_cpu.ALU.u_wallace._2787_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._8386_  (.A1(\u_cpu.ALU.u_wallace._2783_ ),
    .A2(\u_cpu.ALU.u_wallace._2785_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2787_ ),
    .Y(\u_cpu.ALU.u_wallace._2788_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._8387_  (.A1(\u_cpu.ALU.u_wallace._1211_ ),
    .A2(\u_cpu.ALU.u_wallace._2780_ ),
    .B1(\u_cpu.ALU.u_wallace._1392_ ),
    .C1(\u_cpu.ALU.u_wallace._0198_ ),
    .D1(\u_cpu.ALU.u_wallace._2782_ ),
    .Y(\u_cpu.ALU.u_wallace._2789_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8388_  (.A1(\u_cpu.ALU.u_wallace._0198_ ),
    .A2(\u_cpu.ALU.u_wallace._1392_ ),
    .B1(\u_cpu.ALU.u_wallace._2784_ ),
    .B2(\u_cpu.ALU.u_wallace._2782_ ),
    .X(\u_cpu.ALU.u_wallace._2791_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8389_  (.A(\u_cpu.ALU.u_wallace._2787_ ),
    .B(\u_cpu.ALU.u_wallace._2789_ ),
    .C(\u_cpu.ALU.u_wallace._2791_ ),
    .Y(\u_cpu.ALU.u_wallace._2792_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8390_  (.A(\u_cpu.ALU.u_wallace._1322_ ),
    .B(\u_cpu.ALU.u_wallace._0906_ ),
    .C(\u_cpu.ALU.SrcB[21] ),
    .D(\u_cpu.ALU.SrcB[22] ),
    .X(\u_cpu.ALU.u_wallace._2793_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8391_  (.A(\u_cpu.ALU.u_wallace._2793_ ),
    .X(\u_cpu.ALU.u_wallace._2794_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8392_  (.A1(\u_cpu.ALU.u_wallace._1333_ ),
    .A2(\u_cpu.ALU.u_wallace._1610_ ),
    .B1(\u_cpu.ALU.u_wallace._1824_ ),
    .B2(\u_cpu.ALU.u_wallace._0917_ ),
    .Y(\u_cpu.ALU.u_wallace._2795_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8393_  (.A1_N(\u_cpu.ALU.u_wallace._2788_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2792_ ),
    .B1(\u_cpu.ALU.u_wallace._2794_ ),
    .B2(\u_cpu.ALU.u_wallace._2795_ ),
    .Y(\u_cpu.ALU.u_wallace._2796_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8394_  (.A(\u_cpu.ALU.u_wallace._2794_ ),
    .B(\u_cpu.ALU.u_wallace._2795_ ),
    .Y(\u_cpu.ALU.u_wallace._2797_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8395_  (.A(\u_cpu.ALU.u_wallace._2788_ ),
    .B(\u_cpu.ALU.u_wallace._2792_ ),
    .C(\u_cpu.ALU.u_wallace._2797_ ),
    .Y(\u_cpu.ALU.u_wallace._2798_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._8396_  (.A(\u_cpu.ALU.u_wallace._2796_ ),
    .B(\u_cpu.ALU.u_wallace._2798_ ),
    .X(\u_cpu.ALU.u_wallace._2799_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8397_  (.A1(\u_cpu.ALU.u_wallace._2776_ ),
    .A2(\u_cpu.ALU.u_wallace._2778_ ),
    .B1(\u_cpu.ALU.u_wallace._2799_ ),
    .Y(\u_cpu.ALU.u_wallace._2800_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU.u_wallace._8398_  (.A1_N(\u_cpu.ALU.u_wallace._2788_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2792_ ),
    .B1(\u_cpu.ALU.u_wallace._2794_ ),
    .B2(\u_cpu.ALU.u_wallace._2795_ ),
    .X(\u_cpu.ALU.u_wallace._2802_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8399_  (.A(\u_cpu.ALU.u_wallace._2788_ ),
    .B(\u_cpu.ALU.u_wallace._2792_ ),
    .C(\u_cpu.ALU.u_wallace._2797_ ),
    .X(\u_cpu.ALU.u_wallace._2803_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8400_  (.A1(\u_cpu.ALU.u_wallace._2532_ ),
    .A2(\u_cpu.ALU.u_wallace._2777_ ),
    .B1(\u_cpu.ALU.u_wallace._2770_ ),
    .C1(\u_cpu.ALU.u_wallace._2773_ ),
    .X(\u_cpu.ALU.u_wallace._2804_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8401_  (.A1(\u_cpu.ALU.u_wallace._2802_ ),
    .A2(\u_cpu.ALU.u_wallace._2803_ ),
    .B1(\u_cpu.ALU.u_wallace._2775_ ),
    .B2(\u_cpu.ALU.u_wallace._2804_ ),
    .Y(\u_cpu.ALU.u_wallace._2805_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8402_  (.A1(\u_cpu.ALU.u_wallace._2775_ ),
    .A2(\u_cpu.ALU.u_wallace._2800_ ),
    .B1(\u_cpu.ALU.u_wallace._2805_ ),
    .Y(\u_cpu.ALU.u_wallace._2806_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._8403_  (.A(\u_cpu.ALU.u_wallace._2547_ ),
    .Y(\u_cpu.ALU.u_wallace._2807_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8404_  (.A1_N(\u_cpu.ALU.u_wallace._2759_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2806_ ),
    .B1(\u_cpu.ALU.u_wallace._2557_ ),
    .B2(\u_cpu.ALU.u_wallace._2807_ ),
    .Y(\u_cpu.ALU.u_wallace._2808_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8405_  (.A1(\u_cpu.ALU.u_wallace._2693_ ),
    .A2(\u_cpu.ALU.u_wallace._2677_ ),
    .B1(\u_cpu.ALU.u_wallace._2758_ ),
    .X(\u_cpu.ALU.u_wallace._2809_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8406_  (.A1(\u_cpu.ALU.u_wallace._2775_ ),
    .A2(\u_cpu.ALU.u_wallace._2800_ ),
    .B1(\u_cpu.ALU.u_wallace._2805_ ),
    .C1(\u_cpu.ALU.u_wallace._2809_ ),
    .X(\u_cpu.ALU.u_wallace._2810_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8407_  (.A1(\u_cpu.ALU.u_wallace._2770_ ),
    .A2(\u_cpu.ALU.u_wallace._2773_ ),
    .B1(\u_cpu.ALU.u_wallace._2774_ ),
    .X(\u_cpu.ALU.u_wallace._2811_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8408_  (.A1(\u_cpu.ALU.u_wallace._2776_ ),
    .A2(\u_cpu.ALU.u_wallace._2778_ ),
    .B1(\u_cpu.ALU.u_wallace._2799_ ),
    .C1(\u_cpu.ALU.u_wallace._2811_ ),
    .Y(\u_cpu.ALU.u_wallace._2813_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8409_  (.A1(\u_cpu.ALU.u_wallace._2805_ ),
    .A2(\u_cpu.ALU.u_wallace._2813_ ),
    .B1(\u_cpu.ALU.u_wallace._2809_ ),
    .Y(\u_cpu.ALU.u_wallace._2814_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8410_  (.A1(\u_cpu.ALU.u_wallace._2518_ ),
    .A2(\u_cpu.ALU.u_wallace._2519_ ),
    .A3(\u_cpu.ALU.u_wallace._2541_ ),
    .B1(\u_cpu.ALU.u_wallace._2807_ ),
    .X(\u_cpu.ALU.u_wallace._2815_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._8411_  (.A1(\u_cpu.ALU.u_wallace._2814_ ),
    .A2(\u_cpu.ALU.u_wallace._2810_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2815_ ),
    .Y(\u_cpu.ALU.u_wallace._2816_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8412_  (.A1(\u_cpu.ALU.u_wallace._2625_ ),
    .A2(\u_cpu.ALU.u_wallace._2620_ ),
    .B1(\u_cpu.ALU.u_wallace._2627_ ),
    .Y(\u_cpu.ALU.u_wallace._2817_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._8413_  (.A1(\u_cpu.ALU.u_wallace._2620_ ),
    .A2(\u_cpu.ALU.u_wallace._2817_ ),
    .B1(\u_cpu.ALU.u_wallace._2682_ ),
    .X(\u_cpu.ALU.u_wallace._2818_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8414_  (.A(\u_cpu.ALU.u_wallace._2684_ ),
    .B(\u_cpu.ALU.u_wallace._2630_ ),
    .Y(\u_cpu.ALU.u_wallace._2819_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8415_  (.A1_N(\u_cpu.ALU.u_wallace._2818_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2819_ ),
    .B1(\u_cpu.ALU.u_wallace._2608_ ),
    .B2(\u_cpu.ALU.u_wallace._2631_ ),
    .Y(\u_cpu.ALU.u_wallace._2820_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._8416_  (.A1_N(\u_cpu.ALU.u_wallace._2678_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2680_ ),
    .B1(\u_cpu.ALU.u_wallace._2687_ ),
    .B2(\u_cpu.ALU.u_wallace._2820_ ),
    .Y(\u_cpu.ALU.u_wallace._2821_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8417_  (.A(\u_cpu.ALU.u_wallace._4609_ ),
    .B(\u_cpu.ALU.u_wallace._0325_ ),
    .Y(\u_cpu.ALU.u_wallace._2822_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8418_  (.A(\u_cpu.ALU.u_wallace._2822_ ),
    .B(\u_cpu.ALU.u_wallace._2647_ ),
    .Y(\u_cpu.ALU.u_wallace._2824_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8419_  (.A1(\u_cpu.ALU.u_wallace._4848_ ),
    .A2(\u_cpu.ALU.u_wallace._1073_ ),
    .B1(\u_cpu.ALU.u_wallace._0802_ ),
    .B2(\u_cpu.ALU.u_wallace._4720_ ),
    .X(\u_cpu.ALU.u_wallace._2825_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8420_  (.A(\u_cpu.ALU.u_wallace._4594_ ),
    .B(\u_cpu.ALU.u_wallace._4848_ ),
    .C(\u_cpu.ALU.u_wallace._0642_ ),
    .D(\u_cpu.ALU.u_wallace._0802_ ),
    .Y(\u_cpu.ALU.u_wallace._2826_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8421_  (.A(\u_cpu.ALU.u_wallace._2825_ ),
    .B(\u_cpu.ALU.u_wallace._1075_ ),
    .C(\u_cpu.ALU.u_wallace._4604_ ),
    .D(\u_cpu.ALU.u_wallace._2826_ ),
    .Y(\u_cpu.ALU.u_wallace._2827_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8422_  (.A(\u_cpu.ALU.u_wallace._4847_ ),
    .B(\u_cpu.ALU.u_wallace._0045_ ),
    .C(\u_cpu.ALU.u_wallace._1073_ ),
    .D(\u_cpu.ALU.u_wallace._1084_ ),
    .X(\u_cpu.ALU.u_wallace._2828_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8423_  (.A1(\u_cpu.ALU.u_wallace._4848_ ),
    .A2(\u_cpu.ALU.u_wallace._1073_ ),
    .B1(\u_cpu.ALU.u_wallace._0802_ ),
    .B2(\u_cpu.ALU.u_wallace._4720_ ),
    .Y(\u_cpu.ALU.u_wallace._2829_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8424_  (.A1(\u_cpu.ALU.u_wallace._4602_ ),
    .A2(\u_cpu.ALU.u_wallace._0442_ ),
    .B1(\u_cpu.ALU.u_wallace._2828_ ),
    .B2(\u_cpu.ALU.u_wallace._2829_ ),
    .Y(\u_cpu.ALU.u_wallace._2830_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8425_  (.A1(\u_cpu.ALU.u_wallace._2646_ ),
    .A2(\u_cpu.ALU.u_wallace._2824_ ),
    .B1(\u_cpu.ALU.u_wallace._2827_ ),
    .C1(\u_cpu.ALU.u_wallace._2830_ ),
    .X(\u_cpu.ALU.u_wallace._2831_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._8426_  (.A1_N(\u_cpu.ALU.u_wallace._4602_ ),
    .A2_N(\u_cpu.ALU.u_wallace._0442_ ),
    .B1(\u_cpu.ALU.u_wallace._2826_ ),
    .B2(\u_cpu.ALU.u_wallace._2825_ ),
    .Y(\u_cpu.ALU.u_wallace._2832_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8427_  (.A(\u_cpu.ALU.u_wallace._4604_ ),
    .B(\u_cpu.ALU.u_wallace._0850_ ),
    .Y(\u_cpu.ALU.u_wallace._2833_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._8428_  (.A(\u_cpu.ALU.u_wallace._2829_ ),
    .B(\u_cpu.ALU.u_wallace._2833_ ),
    .C(\u_cpu.ALU.u_wallace._2828_ ),
    .Y(\u_cpu.ALU.u_wallace._2835_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._8429_  (.A1(\u_cpu.ALU.u_wallace._2647_ ),
    .A2(\u_cpu.ALU.u_wallace._2822_ ),
    .B1(\u_cpu.ALU.u_wallace._2832_ ),
    .B2(\u_cpu.ALU.u_wallace._2835_ ),
    .C1(\u_cpu.ALU.u_wallace._2651_ ),
    .Y(\u_cpu.ALU.u_wallace._2836_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8430_  (.A1(\u_cpu.ALU.u_wallace._0144_ ),
    .A2(\u_cpu.ALU.u_wallace._0313_ ),
    .B1(\u_cpu.ALU.u_wallace._0330_ ),
    .B2(\u_cpu.ALU.u_wallace._4731_ ),
    .X(\u_cpu.ALU.u_wallace._2837_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8431_  (.A(\u_cpu.ALU.u_wallace._4837_ ),
    .B(\u_cpu.ALU.u_wallace._0029_ ),
    .C(\u_cpu.ALU.u_wallace._0179_ ),
    .D(\u_cpu.ALU.u_wallace._0325_ ),
    .Y(\u_cpu.ALU.u_wallace._2838_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8432_  (.A(\u_cpu.ALU.u_wallace._0319_ ),
    .B(\u_cpu.ALU.u_wallace._0033_ ),
    .Y(\u_cpu.ALU.u_wallace._2839_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8433_  (.A1(\u_cpu.ALU.u_wallace._2837_ ),
    .A2(\u_cpu.ALU.u_wallace._2838_ ),
    .B1(\u_cpu.ALU.u_wallace._2839_ ),
    .X(\u_cpu.ALU.u_wallace._2840_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8434_  (.A1(\u_cpu.ALU.u_wallace._0365_ ),
    .A2(\u_cpu.ALU.u_wallace._0313_ ),
    .B1(\u_cpu.ALU.u_wallace._0330_ ),
    .B2(\u_cpu.ALU.u_wallace._4731_ ),
    .Y(\u_cpu.ALU.u_wallace._2841_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8435_  (.A(\u_cpu.ALU.u_wallace._4836_ ),
    .B(\u_cpu.ALU.u_wallace._4841_ ),
    .C(\u_cpu.ALU.u_wallace._0177_ ),
    .D(\u_cpu.ALU.u_wallace._0332_ ),
    .X(\u_cpu.ALU.u_wallace._2842_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._8436_  (.A1(\u_cpu.ALU.u_wallace._0319_ ),
    .A2(\u_cpu.ALU.u_wallace._0363_ ),
    .B1(\u_cpu.ALU.u_wallace._2841_ ),
    .C1(\u_cpu.ALU.u_wallace._2842_ ),
    .X(\u_cpu.ALU.u_wallace._2843_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8437_  (.A(\u_cpu.ALU.u_wallace._2840_ ),
    .B(\u_cpu.ALU.u_wallace._2843_ ),
    .Y(\u_cpu.ALU.u_wallace._2844_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8438_  (.A(\u_cpu.ALU.u_wallace._2836_ ),
    .B(\u_cpu.ALU.u_wallace._2844_ ),
    .Y(\u_cpu.ALU.u_wallace._2846_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8439_  (.A1(\u_cpu.ALU.u_wallace._2650_ ),
    .A2(\u_cpu.ALU.u_wallace._1974_ ),
    .A3(\u_cpu.ALU.u_wallace._4610_ ),
    .B1(\u_cpu.ALU.u_wallace._2646_ ),
    .X(\u_cpu.ALU.u_wallace._2847_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8440_  (.A1(\u_cpu.ALU.u_wallace._2827_ ),
    .A2(\u_cpu.ALU.u_wallace._2830_ ),
    .B1(\u_cpu.ALU.u_wallace._2847_ ),
    .Y(\u_cpu.ALU.u_wallace._2848_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._8441_  (.A1(\u_cpu.ALU.u_wallace._2831_ ),
    .A2(\u_cpu.ALU.u_wallace._2848_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2844_ ),
    .Y(\u_cpu.ALU.u_wallace._2849_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8442_  (.A1(\u_cpu.ALU.u_wallace._2831_ ),
    .A2(\u_cpu.ALU.u_wallace._2846_ ),
    .B1(\u_cpu.ALU.u_wallace._2849_ ),
    .C1(\u_cpu.ALU.u_wallace._2817_ ),
    .X(\u_cpu.ALU.u_wallace._2850_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8443_  (.A1(\u_cpu.ALU.u_wallace._2831_ ),
    .A2(\u_cpu.ALU.u_wallace._2846_ ),
    .B1(\u_cpu.ALU.u_wallace._2849_ ),
    .Y(\u_cpu.ALU.u_wallace._2851_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._8444_  (.A1(\u_cpu.ALU.u_wallace._2625_ ),
    .A2(\u_cpu.ALU.u_wallace._2620_ ),
    .B1(\u_cpu.ALU.u_wallace._2627_ ),
    .X(\u_cpu.ALU.u_wallace._2852_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8445_  (.A1(\u_cpu.ALU.u_wallace._2673_ ),
    .A2(\u_cpu.ALU.u_wallace._2662_ ),
    .B1(\u_cpu.ALU.u_wallace._2851_ ),
    .B2(\u_cpu.ALU.u_wallace._2852_ ),
    .X(\u_cpu.ALU.u_wallace._2853_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8446_  (.A1(\u_cpu.ALU.u_wallace._2646_ ),
    .A2(\u_cpu.ALU.u_wallace._2824_ ),
    .B1(\u_cpu.ALU.u_wallace._2830_ ),
    .Y(\u_cpu.ALU.u_wallace._2854_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8447_  (.A1(\u_cpu.ALU.u_wallace._2835_ ),
    .A2(\u_cpu.ALU.u_wallace._2854_ ),
    .B1(\u_cpu.ALU.u_wallace._2844_ ),
    .C1(\u_cpu.ALU.u_wallace._2836_ ),
    .Y(\u_cpu.ALU.u_wallace._2855_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8448_  (.A1(\u_cpu.ALU.u_wallace._2855_ ),
    .A2(\u_cpu.ALU.u_wallace._2849_ ),
    .B1(\u_cpu.ALU.u_wallace._2817_ ),
    .Y(\u_cpu.ALU.u_wallace._2857_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._8449_  (.A1(\u_cpu.ALU.u_wallace._2664_ ),
    .A2(\u_cpu.ALU.u_wallace._2666_ ),
    .A3(\u_cpu.ALU.u_wallace._2668_ ),
    .B1(\u_cpu.ALU.u_wallace._2673_ ),
    .X(\u_cpu.ALU.u_wallace._2858_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8450_  (.A1(\u_cpu.ALU.u_wallace._2850_ ),
    .A2(\u_cpu.ALU.u_wallace._2857_ ),
    .B1(\u_cpu.ALU.u_wallace._2858_ ),
    .Y(\u_cpu.ALU.u_wallace._2859_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8451_  (.A(\u_cpu.ALU.u_wallace._2584_ ),
    .B(\u_cpu.ALU.u_wallace._2579_ ),
    .Y(\u_cpu.ALU.u_wallace._2860_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8452_  (.A1(\u_cpu.ALU.u_wallace._2588_ ),
    .A2(\u_cpu.ALU.u_wallace._2590_ ),
    .B1(\u_cpu.ALU.u_wallace._2592_ ),
    .Y(\u_cpu.ALU.u_wallace._2861_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8453_  (.A1(\u_cpu.ALU.u_wallace._2860_ ),
    .A2(\u_cpu.ALU.u_wallace._2605_ ),
    .B1(\u_cpu.ALU.u_wallace._2861_ ),
    .Y(\u_cpu.ALU.u_wallace._2862_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8454_  (.A(\u_cpu.ALU.u_wallace._1826_ ),
    .B(\u_cpu.ALU.u_wallace._1090_ ),
    .Y(\u_cpu.ALU.u_wallace._2863_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8455_  (.A(\u_cpu.ALU.u_wallace._4449_ ),
    .B(\u_cpu.ALU.u_wallace._0629_ ),
    .Y(\u_cpu.ALU.u_wallace._2864_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8456_  (.A1(\u_cpu.ALU.u_wallace._2863_ ),
    .A2(\u_cpu.ALU.u_wallace._2864_ ),
    .B1(\u_cpu.ALU.u_wallace._2602_ ),
    .Y(\u_cpu.ALU.u_wallace._2865_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8457_  (.A1(\u_cpu.ALU.u_wallace._4444_ ),
    .A2(\u_cpu.ALU.u_wallace._0813_ ),
    .B1(\u_cpu.ALU.u_wallace._1270_ ),
    .B2(\u_cpu.ALU.u_wallace._3678_ ),
    .X(\u_cpu.ALU.u_wallace._2866_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8458_  (.A(\u_cpu.ALU.u_wallace._4645_ ),
    .B(\u_cpu.ALU.u_wallace._4562_ ),
    .C(\u_cpu.ALU.u_wallace._0639_ ),
    .D(\u_cpu.ALU.u_wallace._1270_ ),
    .Y(\u_cpu.ALU.u_wallace._2868_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8459_  (.A(\u_cpu.ALU.SrcA[26] ),
    .X(\u_cpu.ALU.u_wallace._2869_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8460_  (.A(\u_cpu.ALU.u_wallace._2866_ ),
    .B(\u_cpu.ALU.u_wallace._2868_ ),
    .C(\u_cpu.ALU.u_wallace._0873_ ),
    .D(\u_cpu.ALU.u_wallace._2869_ ),
    .Y(\u_cpu.ALU.u_wallace._2870_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._8461_  (.A(\u_cpu.ALU.SrcA[26] ),
    .Y(\u_cpu.ALU.u_wallace._2871_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8462_  (.A1(\u_cpu.ALU.u_wallace._4562_ ),
    .A2(\u_cpu.ALU.u_wallace._0639_ ),
    .B1(\u_cpu.ALU.u_wallace._1270_ ),
    .B2(\u_cpu.ALU.u_wallace._4645_ ),
    .Y(\u_cpu.ALU.u_wallace._2872_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8463_  (.A(\u_cpu.ALU.u_wallace._3678_ ),
    .B(\u_cpu.ALU.u_wallace._4444_ ),
    .C(\u_cpu.ALU.u_wallace._0813_ ),
    .D(\u_cpu.ALU.u_wallace._1270_ ),
    .X(\u_cpu.ALU.u_wallace._2873_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8464_  (.A1(\u_cpu.ALU.u_wallace._4923_ ),
    .A2(\u_cpu.ALU.u_wallace._2871_ ),
    .B1(\u_cpu.ALU.u_wallace._2872_ ),
    .B2(\u_cpu.ALU.u_wallace._2873_ ),
    .Y(\u_cpu.ALU.u_wallace._2874_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8465_  (.A1(\u_cpu.ALU.u_wallace._2583_ ),
    .A2(\u_cpu.ALU.u_wallace._2865_ ),
    .B1(\u_cpu.ALU.u_wallace._2870_ ),
    .C1(\u_cpu.ALU.u_wallace._2874_ ),
    .X(\u_cpu.ALU.u_wallace._2875_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8466_  (.A1(\u_cpu.ALU.u_wallace._0086_ ),
    .A2(\u_cpu.ALU.u_wallace._2869_ ),
    .B1(\u_cpu.ALU.u_wallace._2866_ ),
    .B2(\u_cpu.ALU.u_wallace._2868_ ),
    .Y(\u_cpu.ALU.u_wallace._2876_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8467_  (.A(\u_cpu.ALU.u_wallace._2757_ ),
    .B(\u_cpu.ALU.u_wallace._2869_ ),
    .Y(\u_cpu.ALU.u_wallace._2877_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._8468_  (.A(\u_cpu.ALU.u_wallace._2877_ ),
    .B(\u_cpu.ALU.u_wallace._2872_ ),
    .C(\u_cpu.ALU.u_wallace._2873_ ),
    .Y(\u_cpu.ALU.u_wallace._2879_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8469_  (.A1(\u_cpu.ALU.u_wallace._2602_ ),
    .A2(\u_cpu.ALU.u_wallace._2581_ ),
    .B1(\u_cpu.ALU.u_wallace._2577_ ),
    .Y(\u_cpu.ALU.u_wallace._2880_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._8470_  (.A1(\u_cpu.ALU.u_wallace._2876_ ),
    .A2(\u_cpu.ALU.u_wallace._2879_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2880_ ),
    .Y(\u_cpu.ALU.u_wallace._2881_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8471_  (.A(\u_cpu.ALU.u_wallace._2000_ ),
    .X(\u_cpu.ALU.u_wallace._2882_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8472_  (.A1(\u_cpu.ALU.u_wallace._1968_ ),
    .A2(\u_cpu.ALU.u_wallace._2226_ ),
    .B1(\u_cpu.ALU.SrcA[25] ),
    .B2(\u_cpu.ALU.u_wallace._4657_ ),
    .X(\u_cpu.ALU.u_wallace._2883_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8473_  (.A(\u_cpu.ALU.u_wallace._1158_ ),
    .B(\u_cpu.ALU.u_wallace._1169_ ),
    .C(\u_cpu.ALU.u_wallace._2226_ ),
    .D(\u_cpu.ALU.u_wallace._2578_ ),
    .Y(\u_cpu.ALU.u_wallace._2884_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8474_  (.A1(\u_cpu.ALU.u_wallace._4662_ ),
    .A2(\u_cpu.ALU.u_wallace._2882_ ),
    .B1(\u_cpu.ALU.u_wallace._2883_ ),
    .B2(\u_cpu.ALU.u_wallace._2884_ ),
    .Y(\u_cpu.ALU.u_wallace._2885_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8475_  (.A(\u_cpu.ALU.u_wallace._0840_ ),
    .B(\u_cpu.ALU.u_wallace._2002_ ),
    .Y(\u_cpu.ALU.u_wallace._2886_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8476_  (.A1(\u_cpu.ALU.u_wallace._1169_ ),
    .A2(\u_cpu.ALU.u_wallace._2226_ ),
    .B1(\u_cpu.ALU.u_wallace._2578_ ),
    .B2(\u_cpu.ALU.u_wallace._0523_ ),
    .Y(\u_cpu.ALU.u_wallace._2887_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8477_  (.A(\u_cpu.ALU.u_wallace._4657_ ),
    .B(\u_cpu.ALU.u_wallace._4658_ ),
    .C(\u_cpu.ALU.u_wallace._2226_ ),
    .D(\u_cpu.ALU.SrcA[25] ),
    .X(\u_cpu.ALU.u_wallace._2888_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._8478_  (.A(\u_cpu.ALU.u_wallace._2886_ ),
    .B(\u_cpu.ALU.u_wallace._2887_ ),
    .C(\u_cpu.ALU.u_wallace._2888_ ),
    .Y(\u_cpu.ALU.u_wallace._2890_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8479_  (.A(\u_cpu.ALU.u_wallace._2885_ ),
    .B(\u_cpu.ALU.u_wallace._2890_ ),
    .Y(\u_cpu.ALU.u_wallace._2891_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8480_  (.A(\u_cpu.ALU.u_wallace._2881_ ),
    .B(\u_cpu.ALU.u_wallace._2891_ ),
    .Y(\u_cpu.ALU.u_wallace._2892_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8481_  (.A1(\u_cpu.ALU.u_wallace._2874_ ),
    .A2(\u_cpu.ALU.u_wallace._2870_ ),
    .B1(\u_cpu.ALU.u_wallace._2880_ ),
    .Y(\u_cpu.ALU.u_wallace._2893_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8482_  (.A1(\u_cpu.ALU.u_wallace._2885_ ),
    .A2(\u_cpu.ALU.u_wallace._2890_ ),
    .B1(\u_cpu.ALU.u_wallace._2875_ ),
    .B2(\u_cpu.ALU.u_wallace._2893_ ),
    .Y(\u_cpu.ALU.u_wallace._2894_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._8483_  (.A1(\u_cpu.ALU.u_wallace._2585_ ),
    .A2(\u_cpu.ALU.u_wallace._2862_ ),
    .B1(\u_cpu.ALU.u_wallace._2875_ ),
    .B2(\u_cpu.ALU.u_wallace._2892_ ),
    .C1(\u_cpu.ALU.u_wallace._2894_ ),
    .Y(\u_cpu.ALU.u_wallace._2895_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8484_  (.A1(\u_cpu.ALU.u_wallace._2875_ ),
    .A2(\u_cpu.ALU.u_wallace._2893_ ),
    .B1(\u_cpu.ALU.u_wallace._2891_ ),
    .Y(\u_cpu.ALU.u_wallace._2896_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8485_  (.A1(\u_cpu.ALU.u_wallace._2583_ ),
    .A2(\u_cpu.ALU.u_wallace._2865_ ),
    .B1(\u_cpu.ALU.u_wallace._2870_ ),
    .C1(\u_cpu.ALU.u_wallace._2874_ ),
    .Y(\u_cpu.ALU.u_wallace._2897_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8486_  (.A1(\u_cpu.ALU.u_wallace._2885_ ),
    .A2(\u_cpu.ALU.u_wallace._2890_ ),
    .B1(\u_cpu.ALU.u_wallace._2897_ ),
    .C1(\u_cpu.ALU.u_wallace._2881_ ),
    .Y(\u_cpu.ALU.u_wallace._2898_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.ALU.u_wallace._8487_  (.A1(\u_cpu.ALU.u_wallace._2601_ ),
    .A2(\u_cpu.ALU.u_wallace._2603_ ),
    .A3(\u_cpu.ALU.u_wallace._2605_ ),
    .B1(\u_cpu.ALU.u_wallace._2861_ ),
    .B2(\u_cpu.ALU.u_wallace._2587_ ),
    .X(\u_cpu.ALU.u_wallace._2899_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8488_  (.A(\u_cpu.ALU.u_wallace._2896_ ),
    .B(\u_cpu.ALU.u_wallace._2898_ ),
    .C(\u_cpu.ALU.u_wallace._2899_ ),
    .Y(\u_cpu.ALU.u_wallace._2901_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8489_  (.A1(\u_cpu.ALU.u_wallace._2187_ ),
    .A2(\u_cpu.ALU.u_wallace._1531_ ),
    .B1(\u_cpu.ALU.u_wallace._1742_ ),
    .B2(\u_cpu.ALU.u_wallace._2155_ ),
    .Y(\u_cpu.ALU.u_wallace._2902_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8490_  (.A(\u_cpu.ALU.u_wallace._1530_ ),
    .B(\u_cpu.ALU.u_wallace._2056_ ),
    .C(\u_cpu.ALU.u_wallace._1535_ ),
    .D(\u_cpu.ALU.u_wallace._1734_ ),
    .X(\u_cpu.ALU.u_wallace._2903_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8491_  (.A1(\u_cpu.ALU.u_wallace._4539_ ),
    .A2(\u_cpu.ALU.u_wallace._1096_ ),
    .B1(\u_cpu.ALU.u_wallace._2902_ ),
    .B2(\u_cpu.ALU.u_wallace._2903_ ),
    .Y(\u_cpu.ALU.u_wallace._2904_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8492_  (.A1(\u_cpu.ALU.u_wallace._1552_ ),
    .A2(\u_cpu.ALU.u_wallace._1535_ ),
    .B1(\u_cpu.ALU.u_wallace._1742_ ),
    .B2(\u_cpu.ALU.u_wallace._2155_ ),
    .X(\u_cpu.ALU.u_wallace._2905_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8493_  (.A(\u_cpu.ALU.u_wallace._1476_ ),
    .B(\u_cpu.ALU.u_wallace._2187_ ),
    .C(\u_cpu.ALU.u_wallace._1531_ ),
    .D(\u_cpu.ALU.u_wallace._1742_ ),
    .Y(\u_cpu.ALU.u_wallace._2906_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8494_  (.A(\u_cpu.ALU.u_wallace._1101_ ),
    .X(\u_cpu.ALU.u_wallace._2907_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8495_  (.A(\u_cpu.ALU.u_wallace._2905_ ),
    .B(\u_cpu.ALU.u_wallace._2906_ ),
    .C(\u_cpu.ALU.u_wallace._3481_ ),
    .D(\u_cpu.ALU.u_wallace._2907_ ),
    .Y(\u_cpu.ALU.u_wallace._2908_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8496_  (.A1(\u_cpu.ALU.u_wallace._2589_ ),
    .A2(\u_cpu.ALU.u_wallace._2588_ ),
    .B1(\u_cpu.ALU.u_wallace._2597_ ),
    .Y(\u_cpu.ALU.u_wallace._2909_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8497_  (.A1(\u_cpu.ALU.u_wallace._2904_ ),
    .A2(\u_cpu.ALU.u_wallace._2908_ ),
    .B1(\u_cpu.ALU.u_wallace._2909_ ),
    .Y(\u_cpu.ALU.u_wallace._2910_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8498_  (.A(\u_cpu.ALU.u_wallace._2589_ ),
    .B(\u_cpu.ALU.u_wallace._2588_ ),
    .Y(\u_cpu.ALU.u_wallace._2912_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8499_  (.A1(\u_cpu.ALU.u_wallace._2591_ ),
    .A2(\u_cpu.ALU.u_wallace._2912_ ),
    .B1(\u_cpu.ALU.u_wallace._2908_ ),
    .C1(\u_cpu.ALU.u_wallace._2904_ ),
    .X(\u_cpu.ALU.u_wallace._2913_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._8500_  (.A1(\u_cpu.ALU.u_wallace._2284_ ),
    .A2(\u_cpu.ALU.u_wallace._0809_ ),
    .A3(\u_cpu.ALU.u_wallace._2613_ ),
    .B1(\u_cpu.ALU.u_wallace._2611_ ),
    .X(\u_cpu.ALU.u_wallace._2914_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8501_  (.A1(\u_cpu.ALU.u_wallace._2910_ ),
    .A2(\u_cpu.ALU.u_wallace._2913_ ),
    .B1(\u_cpu.ALU.u_wallace._2914_ ),
    .Y(\u_cpu.ALU.u_wallace._2915_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8502_  (.A(\u_cpu.ALU.u_wallace._0815_ ),
    .X(\u_cpu.ALU.u_wallace._2916_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8503_  (.A(\u_cpu.ALU.u_wallace._3481_ ),
    .X(\u_cpu.ALU.u_wallace._2917_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8504_  (.A1(\u_cpu.ALU.u_wallace._2610_ ),
    .A2(\u_cpu.ALU.u_wallace._2916_ ),
    .A3(\u_cpu.ALU.u_wallace._2917_ ),
    .B1(\u_cpu.ALU.u_wallace._2614_ ),
    .X(\u_cpu.ALU.u_wallace._2918_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8505_  (.A1(\u_cpu.ALU.u_wallace._2904_ ),
    .A2(\u_cpu.ALU.u_wallace._2908_ ),
    .B1(\u_cpu.ALU.u_wallace._2909_ ),
    .X(\u_cpu.ALU.u_wallace._2919_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8506_  (.A1(\u_cpu.ALU.u_wallace._2591_ ),
    .A2(\u_cpu.ALU.u_wallace._2912_ ),
    .B1(\u_cpu.ALU.u_wallace._2908_ ),
    .C1(\u_cpu.ALU.u_wallace._2904_ ),
    .Y(\u_cpu.ALU.u_wallace._2920_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8507_  (.A(\u_cpu.ALU.u_wallace._2918_ ),
    .B(\u_cpu.ALU.u_wallace._2919_ ),
    .C(\u_cpu.ALU.u_wallace._2920_ ),
    .Y(\u_cpu.ALU.u_wallace._2921_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8508_  (.A(\u_cpu.ALU.u_wallace._2915_ ),
    .B(\u_cpu.ALU.u_wallace._2921_ ),
    .Y(\u_cpu.ALU.u_wallace._2923_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8509_  (.A1(\u_cpu.ALU.u_wallace._2895_ ),
    .A2(\u_cpu.ALU.u_wallace._2901_ ),
    .B1(\u_cpu.ALU.u_wallace._2923_ ),
    .X(\u_cpu.ALU.u_wallace._2924_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8510_  (.A1(\u_cpu.ALU.u_wallace._2919_ ),
    .A2(\u_cpu.ALU.u_wallace._2920_ ),
    .B1(\u_cpu.ALU.u_wallace._2918_ ),
    .Y(\u_cpu.ALU.u_wallace._2925_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._8511_  (.A(\u_cpu.ALU.u_wallace._2914_ ),
    .B(\u_cpu.ALU.u_wallace._2910_ ),
    .C(\u_cpu.ALU.u_wallace._2913_ ),
    .Y(\u_cpu.ALU.u_wallace._2926_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8512_  (.A1(\u_cpu.ALU.u_wallace._2925_ ),
    .A2(\u_cpu.ALU.u_wallace._2926_ ),
    .B1(\u_cpu.ALU.u_wallace._2895_ ),
    .C1(\u_cpu.ALU.u_wallace._2901_ ),
    .Y(\u_cpu.ALU.u_wallace._2927_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8513_  (.A(\u_cpu.ALU.u_wallace._2682_ ),
    .B(\u_cpu.ALU.u_wallace._2683_ ),
    .Y(\u_cpu.ALU.u_wallace._2928_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8514_  (.A1(\u_cpu.ALU.u_wallace._2928_ ),
    .A2(\u_cpu.ALU.u_wallace._2630_ ),
    .B1(\u_cpu.ALU.u_wallace._2608_ ),
    .Y(\u_cpu.ALU.u_wallace._2929_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8515_  (.A(\u_cpu.ALU.u_wallace._2924_ ),
    .B(\u_cpu.ALU.u_wallace._2927_ ),
    .C(\u_cpu.ALU.u_wallace._2929_ ),
    .Y(\u_cpu.ALU.u_wallace._2930_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8516_  (.A(\u_cpu.ALU.u_wallace._2634_ ),
    .B(\u_cpu.ALU.u_wallace._2635_ ),
    .Y(\u_cpu.ALU.u_wallace._2931_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8517_  (.A1(\u_cpu.ALU.u_wallace._2682_ ),
    .A2(\u_cpu.ALU.u_wallace._2683_ ),
    .B1(\u_cpu.ALU.u_wallace._2931_ ),
    .B2(\u_cpu.ALU.u_wallace._2629_ ),
    .Y(\u_cpu.ALU.u_wallace._2932_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8518_  (.A(\u_cpu.ALU.u_wallace._2915_ ),
    .B(\u_cpu.ALU.u_wallace._2921_ ),
    .C(\u_cpu.ALU.u_wallace._2895_ ),
    .D(\u_cpu.ALU.u_wallace._2901_ ),
    .Y(\u_cpu.ALU.u_wallace._2934_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8519_  (.A(\u_cpu.ALU.u_wallace._2881_ ),
    .B(\u_cpu.ALU.u_wallace._2891_ ),
    .C(\u_cpu.ALU.u_wallace._2897_ ),
    .Y(\u_cpu.ALU.u_wallace._2935_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8520_  (.A1(\u_cpu.ALU.u_wallace._2585_ ),
    .A2(\u_cpu.ALU.u_wallace._2862_ ),
    .B1(\u_cpu.ALU.u_wallace._2935_ ),
    .C1(\u_cpu.ALU.u_wallace._2894_ ),
    .X(\u_cpu.ALU.u_wallace._2936_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._8521_  (.A1(\u_cpu.ALU.u_wallace._2584_ ),
    .A2(\u_cpu.ALU.u_wallace._2579_ ),
    .A3(\u_cpu.ALU.u_wallace._2586_ ),
    .B1(\u_cpu.ALU.u_wallace._2606_ ),
    .B2(\u_cpu.ALU.u_wallace._2594_ ),
    .X(\u_cpu.ALU.u_wallace._2937_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8522_  (.A1(\u_cpu.ALU.u_wallace._2935_ ),
    .A2(\u_cpu.ALU.u_wallace._2894_ ),
    .B1(\u_cpu.ALU.u_wallace._2937_ ),
    .Y(\u_cpu.ALU.u_wallace._2938_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8523_  (.A1(\u_cpu.ALU.u_wallace._2925_ ),
    .A2(\u_cpu.ALU.u_wallace._2926_ ),
    .B1(\u_cpu.ALU.u_wallace._2936_ ),
    .B2(\u_cpu.ALU.u_wallace._2938_ ),
    .Y(\u_cpu.ALU.u_wallace._2939_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8524_  (.A1(\u_cpu.ALU.u_wallace._2608_ ),
    .A2(\u_cpu.ALU.u_wallace._2932_ ),
    .B1(\u_cpu.ALU.u_wallace._2934_ ),
    .C1(\u_cpu.ALU.u_wallace._2939_ ),
    .Y(\u_cpu.ALU.u_wallace._2940_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._8525_  (.A1(\u_cpu.ALU.u_wallace._2850_ ),
    .A2(\u_cpu.ALU.u_wallace._2853_ ),
    .B1(\u_cpu.ALU.u_wallace._2859_ ),
    .C1(\u_cpu.ALU.u_wallace._2930_ ),
    .D1(\u_cpu.ALU.u_wallace._2940_ ),
    .Y(\u_cpu.ALU.u_wallace._2941_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8526_  (.A1(\u_cpu.ALU.u_wallace._2835_ ),
    .A2(\u_cpu.ALU.u_wallace._2854_ ),
    .B1(\u_cpu.ALU.u_wallace._2844_ ),
    .C1(\u_cpu.ALU.u_wallace._2836_ ),
    .X(\u_cpu.ALU.u_wallace._2942_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8527_  (.A1(\u_cpu.ALU.u_wallace._2646_ ),
    .A2(\u_cpu.ALU.u_wallace._2824_ ),
    .B1(\u_cpu.ALU.u_wallace._2827_ ),
    .C1(\u_cpu.ALU.u_wallace._2830_ ),
    .Y(\u_cpu.ALU.u_wallace._2943_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8528_  (.A1(\u_cpu.ALU.u_wallace._2943_ ),
    .A2(\u_cpu.ALU.u_wallace._2836_ ),
    .B1(\u_cpu.ALU.u_wallace._2844_ ),
    .Y(\u_cpu.ALU.u_wallace._2945_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8529_  (.A1(\u_cpu.ALU.u_wallace._2673_ ),
    .A2(\u_cpu.ALU.u_wallace._2662_ ),
    .B1(\u_cpu.ALU.u_wallace._2851_ ),
    .B2(\u_cpu.ALU.u_wallace._2852_ ),
    .Y(\u_cpu.ALU.u_wallace._2946_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._8530_  (.A1(\u_cpu.ALU.u_wallace._2852_ ),
    .A2(\u_cpu.ALU.u_wallace._2942_ ),
    .A3(\u_cpu.ALU.u_wallace._2945_ ),
    .B1(\u_cpu.ALU.u_wallace._2946_ ),
    .X(\u_cpu.ALU.u_wallace._2947_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._8531_  (.A1(\u_cpu.ALU.u_wallace._2654_ ),
    .A2(\u_cpu.ALU.u_wallace._2655_ ),
    .B1(\u_cpu.ALU.u_wallace._2850_ ),
    .B2(\u_cpu.ALU.u_wallace._2857_ ),
    .C1(\u_cpu.ALU.u_wallace._2662_ ),
    .X(\u_cpu.ALU.u_wallace._2948_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8532_  (.A1_N(\u_cpu.ALU.u_wallace._2940_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2930_ ),
    .B1(\u_cpu.ALU.u_wallace._2947_ ),
    .B2(\u_cpu.ALU.u_wallace._2948_ ),
    .Y(\u_cpu.ALU.u_wallace._2949_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8533_  (.A1(\u_cpu.ALU.u_wallace._2640_ ),
    .A2(\u_cpu.ALU.u_wallace._2821_ ),
    .B1(\u_cpu.ALU.u_wallace._2941_ ),
    .C1(\u_cpu.ALU.u_wallace._2949_ ),
    .Y(\u_cpu.ALU.u_wallace._2950_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8534_  (.A1(\u_cpu.ALU.u_wallace._2808_ ),
    .A2(\u_cpu.ALU.u_wallace._2810_ ),
    .B1(\u_cpu.ALU.u_wallace._2816_ ),
    .C1(\u_cpu.ALU.u_wallace._2950_ ),
    .Y(\u_cpu.ALU.u_wallace._2951_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8535_  (.A1(\u_cpu.ALU.u_wallace._2687_ ),
    .A2(\u_cpu.ALU.u_wallace._2820_ ),
    .B1(\u_cpu.ALU.u_wallace._2689_ ),
    .Y(\u_cpu.ALU.u_wallace._2952_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8536_  (.A1(\u_cpu.ALU.u_wallace._2941_ ),
    .A2(\u_cpu.ALU.u_wallace._2949_ ),
    .B1(\u_cpu.ALU.u_wallace._2952_ ),
    .Y(\u_cpu.ALU.u_wallace._2953_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8537_  (.A1(\u_cpu.ALU.u_wallace._2566_ ),
    .A2(\u_cpu.ALU.u_wallace._2562_ ),
    .B1(\u_cpu.ALU.u_wallace._2700_ ),
    .Y(\u_cpu.ALU.u_wallace._2954_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8538_  (.A1(\u_cpu.ALU.u_wallace._2701_ ),
    .A2(\u_cpu.ALU.u_wallace._2716_ ),
    .B1(\u_cpu.ALU.u_wallace._2954_ ),
    .B2(\u_cpu.ALU.u_wallace._2711_ ),
    .Y(\u_cpu.ALU.u_wallace._2956_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8539_  (.A1(\u_cpu.ALU.u_wallace._2805_ ),
    .A2(\u_cpu.ALU.u_wallace._2813_ ),
    .B1(\u_cpu.ALU.u_wallace._2809_ ),
    .X(\u_cpu.ALU.u_wallace._2957_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8540_  (.A1(\u_cpu.ALU.u_wallace._2775_ ),
    .A2(\u_cpu.ALU.u_wallace._2800_ ),
    .B1(\u_cpu.ALU.u_wallace._2805_ ),
    .C1(\u_cpu.ALU.u_wallace._2809_ ),
    .Y(\u_cpu.ALU.u_wallace._2958_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8541_  (.A1(\u_cpu.ALU.u_wallace._2957_ ),
    .A2(\u_cpu.ALU.u_wallace._2958_ ),
    .B1(\u_cpu.ALU.u_wallace._2815_ ),
    .Y(\u_cpu.ALU.u_wallace._2959_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8542_  (.A(\u_cpu.ALU.u_wallace._2957_ ),
    .B(\u_cpu.ALU.u_wallace._2958_ ),
    .C(\u_cpu.ALU.u_wallace._2815_ ),
    .X(\u_cpu.ALU.u_wallace._2960_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8543_  (.A1(\u_cpu.ALU.u_wallace._2640_ ),
    .A2(\u_cpu.ALU.u_wallace._2821_ ),
    .B1(\u_cpu.ALU.u_wallace._2941_ ),
    .C1(\u_cpu.ALU.u_wallace._2949_ ),
    .X(\u_cpu.ALU.u_wallace._2961_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8544_  (.A1(\u_cpu.ALU.u_wallace._2959_ ),
    .A2(\u_cpu.ALU.u_wallace._2960_ ),
    .B1(\u_cpu.ALU.u_wallace._2961_ ),
    .B2(\u_cpu.ALU.u_wallace._2953_ ),
    .Y(\u_cpu.ALU.u_wallace._2962_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8545_  (.A1(\u_cpu.ALU.u_wallace._2951_ ),
    .A2(\u_cpu.ALU.u_wallace._2953_ ),
    .B1(\u_cpu.ALU.u_wallace._2956_ ),
    .C1(\u_cpu.ALU.u_wallace._2962_ ),
    .Y(\u_cpu.ALU.u_wallace._2963_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._8546_  (.A1(\u_cpu.ALU.u_wallace._2701_ ),
    .A2(\u_cpu.ALU.u_wallace._2716_ ),
    .B1(\u_cpu.ALU.u_wallace._2954_ ),
    .B2(\u_cpu.ALU.u_wallace._2711_ ),
    .X(\u_cpu.ALU.u_wallace._2964_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8547_  (.A1(\u_cpu.ALU.u_wallace._2547_ ),
    .A2(\u_cpu.ALU.u_wallace._2565_ ),
    .B1(\u_cpu.ALU.u_wallace._2814_ ),
    .Y(\u_cpu.ALU.u_wallace._2965_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8548_  (.A1(\u_cpu.ALU.u_wallace._2958_ ),
    .A2(\u_cpu.ALU.u_wallace._2965_ ),
    .B1(\u_cpu.ALU.u_wallace._2959_ ),
    .Y(\u_cpu.ALU.u_wallace._2967_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8549_  (.A1(\u_cpu.ALU.u_wallace._2961_ ),
    .A2(\u_cpu.ALU.u_wallace._2953_ ),
    .B1(\u_cpu.ALU.u_wallace._2967_ ),
    .Y(\u_cpu.ALU.u_wallace._2968_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8550_  (.A1(\u_cpu.ALU.u_wallace._2941_ ),
    .A2(\u_cpu.ALU.u_wallace._2949_ ),
    .B1(\u_cpu.ALU.u_wallace._2952_ ),
    .X(\u_cpu.ALU.u_wallace._2969_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8551_  (.A1(\u_cpu.ALU.u_wallace._2959_ ),
    .A2(\u_cpu.ALU.u_wallace._2960_ ),
    .B1(\u_cpu.ALU.u_wallace._2950_ ),
    .C1(\u_cpu.ALU.u_wallace._2969_ ),
    .Y(\u_cpu.ALU.u_wallace._2970_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8552_  (.A(\u_cpu.ALU.u_wallace._2964_ ),
    .B(\u_cpu.ALU.u_wallace._2968_ ),
    .C(\u_cpu.ALU.u_wallace._2970_ ),
    .Y(\u_cpu.ALU.u_wallace._2971_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8553_  (.A1(\u_cpu.ALU.u_wallace._2511_ ),
    .A2(\u_cpu.ALU.u_wallace._2508_ ),
    .A3(\u_cpu.ALU.u_wallace._2509_ ),
    .B1(\u_cpu.ALU.u_wallace._2514_ ),
    .X(\u_cpu.ALU.u_wallace._2972_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8554_  (.A(\u_cpu.ALU.u_wallace._2514_ ),
    .B(\u_cpu.ALU.u_wallace._2509_ ),
    .C(\u_cpu.ALU.u_wallace._2508_ ),
    .D(\u_cpu.ALU.u_wallace._2511_ ),
    .Y(\u_cpu.ALU.u_wallace._2973_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8555_  (.A(\u_cpu.ALU.u_wallace._2972_ ),
    .B(\u_cpu.ALU.u_wallace._2973_ ),
    .Y(\u_cpu.ALU.u_wallace._2974_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8556_  (.A1(\u_cpu.ALU.u_wallace._2519_ ),
    .A2(\u_cpu.ALU.u_wallace._2974_ ),
    .B1(\u_cpu.ALU.u_wallace._2476_ ),
    .Y(\u_cpu.ALU.u_wallace._2975_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8557_  (.A(\u_cpu.ALU.u_wallace._2519_ ),
    .B(\u_cpu.ALU.u_wallace._2476_ ),
    .C(\u_cpu.ALU.u_wallace._2974_ ),
    .X(\u_cpu.ALU.u_wallace._2976_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8558_  (.A1(\u_cpu.ALU.u_wallace._0151_ ),
    .A2(\u_cpu.ALU.SrcB[25] ),
    .B1(\u_cpu.ALU.SrcB[26] ),
    .B2(\u_cpu.ALU.u_wallace._0021_ ),
    .Y(\u_cpu.ALU.u_wallace._2978_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8559_  (.A(\u_cpu.ALU.u_wallace._0994_ ),
    .B(\u_cpu.ALU.u_wallace._0261_ ),
    .C(\u_cpu.ALU.SrcB[25] ),
    .D(\u_cpu.ALU.SrcB[26] ),
    .Y(\u_cpu.ALU.u_wallace._2979_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._8560_  (.A(\u_cpu.ALU.u_wallace._1410_ ),
    .B(\u_cpu.ALU.SrcB[24] ),
    .X(\u_cpu.ALU.u_wallace._2980_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._8561_  (.A_N(\u_cpu.ALU.u_wallace._2978_ ),
    .B(\u_cpu.ALU.u_wallace._2979_ ),
    .C(\u_cpu.ALU.u_wallace._2980_ ),
    .Y(\u_cpu.ALU.u_wallace._2981_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8562_  (.A(\u_cpu.ALU.u_wallace._0021_ ),
    .B(\u_cpu.ALU.u_wallace._0151_ ),
    .C(\u_cpu.ALU.SrcB[25] ),
    .D(\u_cpu.ALU.SrcB[26] ),
    .X(\u_cpu.ALU.u_wallace._2982_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._8563_  (.A1(\u_cpu.ALU.u_wallace._2978_ ),
    .A2(\u_cpu.ALU.u_wallace._2982_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2980_ ),
    .Y(\u_cpu.ALU.u_wallace._2983_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8564_  (.A1(\u_cpu.ALU.u_wallace._2981_ ),
    .A2(\u_cpu.ALU.u_wallace._2983_ ),
    .B1(\u_cpu.ALU.u_wallace._2488_ ),
    .Y(\u_cpu.ALU.u_wallace._2984_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8565_  (.A(\u_cpu.ALU.u_wallace._2983_ ),
    .B(\u_cpu.ALU.u_wallace._2488_ ),
    .C(\u_cpu.ALU.u_wallace._2981_ ),
    .X(\u_cpu.ALU.u_wallace._2985_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8566_  (.A(\u_cpu.ALU.u_wallace._4541_ ),
    .X(\u_cpu.ALU.u_wallace._2986_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.ALU.u_wallace._8567_  (.A1_N(\u_cpu.ALU.u_wallace._2984_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2985_ ),
    .B1(\u_cpu.ALU.u_wallace._2986_ ),
    .B2(\u_cpu.ALU.u_wallace._2134_ ),
    .X(\u_cpu.ALU.u_wallace._2987_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.ALU.u_wallace._8568_  (.A1_N(\u_cpu.ALU.u_wallace._2482_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2484_ ),
    .B1(\u_cpu.ALU.u_wallace._2981_ ),
    .B2(\u_cpu.ALU.u_wallace._2983_ ),
    .X(\u_cpu.ALU.u_wallace._2989_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._8569_  (.A_N(\u_cpu.ALU.u_wallace._2985_ ),
    .B(\u_cpu.ALU.u_wallace._2134_ ),
    .C(\u_cpu.ALU.u_wallace._2986_ ),
    .D(\u_cpu.ALU.u_wallace._2989_ ),
    .Y(\u_cpu.ALU.u_wallace._2990_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._8570_  (.A(\u_cpu.ALU.u_wallace._2987_ ),
    .B(\u_cpu.ALU.u_wallace._2990_ ),
    .X(\u_cpu.ALU.u_wallace._2991_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8571_  (.A1(\u_cpu.ALU.u_wallace._2975_ ),
    .A2(\u_cpu.ALU.u_wallace._2976_ ),
    .B1(\u_cpu.ALU.u_wallace._2991_ ),
    .Y(\u_cpu.ALU.u_wallace._2992_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8572_  (.A1(\u_cpu.ALU.u_wallace._2556_ ),
    .A2(\u_cpu.ALU.u_wallace._2555_ ),
    .B1(\u_cpu.ALU.u_wallace._2476_ ),
    .C1(\u_cpu.ALU.u_wallace._2974_ ),
    .Y(\u_cpu.ALU.u_wallace._2993_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8573_  (.A(\u_cpu.ALU.u_wallace._2987_ ),
    .B(\u_cpu.ALU.u_wallace._2990_ ),
    .Y(\u_cpu.ALU.u_wallace._2994_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._8574_  (.A_N(\u_cpu.ALU.u_wallace._2975_ ),
    .B(\u_cpu.ALU.u_wallace._2993_ ),
    .C(\u_cpu.ALU.u_wallace._2994_ ),
    .Y(\u_cpu.ALU.u_wallace._2995_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8575_  (.A(\u_cpu.ALU.u_wallace._2699_ ),
    .B(\u_cpu.ALU.u_wallace._2992_ ),
    .C(\u_cpu.ALU.u_wallace._2995_ ),
    .Y(\u_cpu.ALU.u_wallace._2996_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8576_  (.A1(\u_cpu.ALU.u_wallace._2559_ ),
    .A2(\u_cpu.ALU.u_wallace._2699_ ),
    .A3(\u_cpu.ALU.u_wallace._2561_ ),
    .B1(\u_cpu.ALU.u_wallace._2996_ ),
    .X(\u_cpu.ALU.u_wallace._2997_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8577_  (.A(\u_cpu.ALU.u_wallace._2992_ ),
    .B(\u_cpu.ALU.u_wallace._2995_ ),
    .Y(\u_cpu.ALU.u_wallace._2998_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8578_  (.A1(\u_cpu.ALU.u_wallace._2566_ ),
    .A2(\u_cpu.ALU.u_wallace._2718_ ),
    .B1(\u_cpu.ALU.u_wallace._2998_ ),
    .Y(\u_cpu.ALU.u_wallace._3000_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._8579_  (.A1(\u_cpu.ALU.u_wallace._2479_ ),
    .A2(\u_cpu.ALU.u_wallace._2490_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2478_ ),
    .Y(\u_cpu.ALU.u_wallace._3001_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._8580_  (.A(\u_cpu.ALU.u_wallace._3001_ ),
    .Y(\u_cpu.ALU.u_wallace._3002_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8581_  (.A1(\u_cpu.ALU.u_wallace._2997_ ),
    .A2(\u_cpu.ALU.u_wallace._3000_ ),
    .B1(\u_cpu.ALU.u_wallace._3002_ ),
    .Y(\u_cpu.ALU.u_wallace._3003_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8582_  (.A1(\u_cpu.ALU.u_wallace._2996_ ),
    .A2(\u_cpu.ALU.u_wallace._2709_ ),
    .B1(\u_cpu.ALU.u_wallace._3002_ ),
    .C1(\u_cpu.ALU.u_wallace._3000_ ),
    .X(\u_cpu.ALU.u_wallace._3004_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8583_  (.A(\u_cpu.ALU.u_wallace._3003_ ),
    .B(\u_cpu.ALU.u_wallace._3004_ ),
    .Y(\u_cpu.ALU.u_wallace._3005_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8584_  (.A1(\u_cpu.ALU.u_wallace._2963_ ),
    .A2(\u_cpu.ALU.u_wallace._2971_ ),
    .B1(\u_cpu.ALU.u_wallace._3005_ ),
    .Y(\u_cpu.ALU.u_wallace._3006_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8585_  (.A(\u_cpu.ALU.u_wallace._2971_ ),
    .B(\u_cpu.ALU.u_wallace._3005_ ),
    .C(\u_cpu.ALU.u_wallace._2963_ ),
    .X(\u_cpu.ALU.u_wallace._3007_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU.u_wallace._8586_  (.A1_N(\u_cpu.ALU.u_wallace._2707_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2731_ ),
    .B1(\u_cpu.ALU.u_wallace._2732_ ),
    .B2(\u_cpu.ALU.u_wallace._2733_ ),
    .X(\u_cpu.ALU.u_wallace._3008_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8587_  (.A1(\u_cpu.ALU.u_wallace._3006_ ),
    .A2(\u_cpu.ALU.u_wallace._3007_ ),
    .B1(\u_cpu.ALU.u_wallace._3008_ ),
    .Y(\u_cpu.ALU.u_wallace._3009_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8588_  (.A(\u_cpu.ALU.u_wallace._2971_ ),
    .B(\u_cpu.ALU.u_wallace._3005_ ),
    .Y(\u_cpu.ALU.u_wallace._3011_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8589_  (.A1(\u_cpu.ALU.u_wallace._2951_ ),
    .A2(\u_cpu.ALU.u_wallace._2953_ ),
    .B1(\u_cpu.ALU.u_wallace._2956_ ),
    .C1(\u_cpu.ALU.u_wallace._2962_ ),
    .X(\u_cpu.ALU.u_wallace._3012_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8590_  (.A1(\u_cpu.ALU.u_wallace._2732_ ),
    .A2(\u_cpu.ALU.u_wallace._2733_ ),
    .B1(\u_cpu.ALU.u_wallace._2715_ ),
    .Y(\u_cpu.ALU.u_wallace._3013_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.ALU.u_wallace._8591_  (.A1_N(\u_cpu.ALU.u_wallace._3003_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3004_ ),
    .B1(\u_cpu.ALU.u_wallace._2963_ ),
    .B2(\u_cpu.ALU.u_wallace._2971_ ),
    .X(\u_cpu.ALU.u_wallace._3014_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8592_  (.A1(\u_cpu.ALU.u_wallace._3011_ ),
    .A2(\u_cpu.ALU.u_wallace._3012_ ),
    .B1(\u_cpu.ALU.u_wallace._3013_ ),
    .C1(\u_cpu.ALU.u_wallace._3014_ ),
    .Y(\u_cpu.ALU.u_wallace._3015_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU.u_wallace._8593_  (.A(\u_cpu.ALU.u_wallace._2498_ ),
    .B(\u_cpu.ALU.u_wallace._2727_ ),
    .X(\u_cpu.ALU.u_wallace._3016_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8594_  (.A1(\u_cpu.ALU.u_wallace._3009_ ),
    .A2(\u_cpu.ALU.u_wallace._3015_ ),
    .B1(\u_cpu.ALU.u_wallace._3016_ ),
    .X(\u_cpu.ALU.u_wallace._3017_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8595_  (.A1(\u_cpu.ALU.u_wallace._2498_ ),
    .A2(\u_cpu.ALU.u_wallace._2727_ ),
    .B1(\u_cpu.ALU.u_wallace._3009_ ),
    .C1(\u_cpu.ALU.u_wallace._3015_ ),
    .Y(\u_cpu.ALU.u_wallace._3018_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8596_  (.A(\u_cpu.ALU.u_wallace._2756_ ),
    .B(\u_cpu.ALU.u_wallace._3017_ ),
    .C(\u_cpu.ALU.u_wallace._3018_ ),
    .Y(\u_cpu.ALU.u_wallace._3019_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8597_  (.A1(\u_cpu.ALU.u_wallace._3009_ ),
    .A2(\u_cpu.ALU.u_wallace._3015_ ),
    .B1(\u_cpu.ALU.u_wallace._3016_ ),
    .Y(\u_cpu.ALU.u_wallace._3020_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8598_  (.A1(\u_cpu.ALU.u_wallace._2498_ ),
    .A2(\u_cpu.ALU.u_wallace._2727_ ),
    .B1(\u_cpu.ALU.u_wallace._3009_ ),
    .C1(\u_cpu.ALU.u_wallace._3015_ ),
    .X(\u_cpu.ALU.u_wallace._3022_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8599_  (.A1(\u_cpu.ALU.u_wallace._2742_ ),
    .A2(\u_cpu.ALU.u_wallace._2738_ ),
    .B1(\u_cpu.ALU.u_wallace._2740_ ),
    .Y(\u_cpu.ALU.u_wallace._3023_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8600_  (.A1(\u_cpu.ALU.u_wallace._3020_ ),
    .A2(\u_cpu.ALU.u_wallace._3022_ ),
    .B1(\u_cpu.ALU.u_wallace._3023_ ),
    .Y(\u_cpu.ALU.u_wallace._3024_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._8601_  (.A1_N(\u_cpu.ALU.u_wallace._2755_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2488_ ),
    .B1(\u_cpu.ALU.u_wallace._3019_ ),
    .B2(\u_cpu.ALU.u_wallace._3024_ ),
    .Y(\u_cpu.ALU.u_wallace._3025_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8602_  (.A(\u_cpu.ALU.u_wallace._2485_ ),
    .B(\u_cpu.ALU.u_wallace._2417_ ),
    .C(\u_cpu.ALU.u_wallace._0370_ ),
    .X(\u_cpu.ALU.u_wallace._3026_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._8603_  (.A1(\u_cpu.ALU.u_wallace._2482_ ),
    .A2(\u_cpu.ALU.u_wallace._2484_ ),
    .B1(\u_cpu.ALU.u_wallace._3019_ ),
    .C1(\u_cpu.ALU.u_wallace._3026_ ),
    .D1(\u_cpu.ALU.u_wallace._3024_ ),
    .X(\u_cpu.ALU.u_wallace._3027_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8604_  (.A(\u_cpu.ALU.u_wallace._2473_ ),
    .B(\u_cpu.ALU.u_wallace._2744_ ),
    .Y(\u_cpu.ALU.u_wallace._3028_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8605_  (.A1(\u_cpu.ALU.u_wallace._2739_ ),
    .A2(\u_cpu.ALU.u_wallace._2744_ ),
    .B1(\u_cpu.ALU.u_wallace._2473_ ),
    .Y(\u_cpu.ALU.u_wallace._3029_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._8606_  (.A1(\u_cpu.ALU.u_wallace._2746_ ),
    .A2(\u_cpu.ALU.u_wallace._3028_ ),
    .B1(\u_cpu.ALU.u_wallace._2401_ ),
    .B2(\u_cpu.ALU.u_wallace._3029_ ),
    .X(\u_cpu.ALU.u_wallace._3030_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8607_  (.A1(\u_cpu.ALU.u_wallace._3025_ ),
    .A2(\u_cpu.ALU.u_wallace._3027_ ),
    .B1(\u_cpu.ALU.u_wallace._3030_ ),
    .Y(\u_cpu.ALU.u_wallace._3031_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8608_  (.A1(\u_cpu.ALU.u_wallace._2746_ ),
    .A2(\u_cpu.ALU.u_wallace._3028_ ),
    .B1(\u_cpu.ALU.u_wallace._2401_ ),
    .B2(\u_cpu.ALU.u_wallace._3029_ ),
    .Y(\u_cpu.ALU.u_wallace._3033_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8609_  (.A1_N(\u_cpu.ALU.u_wallace._3024_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3019_ ),
    .B1(\u_cpu.ALU.u_wallace._2488_ ),
    .B2(\u_cpu.ALU.u_wallace._2755_ ),
    .Y(\u_cpu.ALU.u_wallace._3034_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._8610_  (.A1(\u_cpu.ALU.u_wallace._2482_ ),
    .A2(\u_cpu.ALU.u_wallace._2484_ ),
    .B1(\u_cpu.ALU.u_wallace._3019_ ),
    .C1(\u_cpu.ALU.u_wallace._3026_ ),
    .D1(\u_cpu.ALU.u_wallace._3024_ ),
    .Y(\u_cpu.ALU.u_wallace._3035_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8611_  (.A(\u_cpu.ALU.u_wallace._3033_ ),
    .B(\u_cpu.ALU.u_wallace._3034_ ),
    .C(\u_cpu.ALU.u_wallace._3035_ ),
    .Y(\u_cpu.ALU.u_wallace._3036_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._8612_  (.A(\u_cpu.ALU.u_wallace._3031_ ),
    .B(\u_cpu.ALU.u_wallace._3036_ ),
    .X(\u_cpu.ALU.u_wallace._3037_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8613_  (.A1(\u_cpu.ALU.u_wallace._2746_ ),
    .A2(\u_cpu.ALU.u_wallace._3028_ ),
    .B1(\u_cpu.ALU.u_wallace._2749_ ),
    .Y(\u_cpu.ALU.u_wallace._3038_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._8614_  (.A1_N(\u_cpu.ALU.u_wallace._2452_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2448_ ),
    .B1(\u_cpu.ALU.u_wallace._3038_ ),
    .B2(\u_cpu.ALU.u_wallace._2401_ ),
    .Y(\u_cpu.ALU.u_wallace._3039_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8615_  (.A1(\u_cpu.ALU.u_wallace._2752_ ),
    .A2(\u_cpu.ALU.u_wallace._2753_ ),
    .B1(\u_cpu.ALU.u_wallace._2455_ ),
    .Y(\u_cpu.ALU.u_wallace._3040_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8616_  (.A1(\u_cpu.ALU.u_wallace._2751_ ),
    .A2(\u_cpu.ALU.u_wallace._3039_ ),
    .B1(\u_cpu.ALU.u_wallace._3040_ ),
    .B2(\u_cpu.ALU.u_wallace._2468_ ),
    .Y(\u_cpu.ALU.u_wallace._3041_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu.ALU.u_wallace._8617_  (.A(\u_cpu.ALU.u_wallace._3037_ ),
    .B(\u_cpu.ALU.u_wallace._3041_ ),
    .Y(\u_cpu.ALU.Product_Wallace[26] ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.ALU.u_wallace._8618_  (.A1(\u_cpu.ALU.u_wallace._2959_ ),
    .A2(\u_cpu.ALU.u_wallace._2960_ ),
    .A3(\u_cpu.ALU.u_wallace._2953_ ),
    .B1(\u_cpu.ALU.u_wallace._2950_ ),
    .Y(\u_cpu.ALU.u_wallace._3043_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._8619_  (.A(\u_cpu.ALU.u_wallace._2934_ ),
    .Y(\u_cpu.ALU.u_wallace._3044_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8620_  (.A1(\u_cpu.ALU.u_wallace._2608_ ),
    .A2(\u_cpu.ALU.u_wallace._2932_ ),
    .B1(\u_cpu.ALU.u_wallace._2939_ ),
    .Y(\u_cpu.ALU.u_wallace._3045_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8621_  (.A(\u_cpu.ALU.u_wallace._2817_ ),
    .B(\u_cpu.ALU.u_wallace._2849_ ),
    .Y(\u_cpu.ALU.u_wallace._3046_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8622_  (.A1(\u_cpu.ALU.u_wallace._2942_ ),
    .A2(\u_cpu.ALU.u_wallace._2945_ ),
    .B1(\u_cpu.ALU.u_wallace._2852_ ),
    .Y(\u_cpu.ALU.u_wallace._3047_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8623_  (.A1(\u_cpu.ALU.u_wallace._2942_ ),
    .A2(\u_cpu.ALU.u_wallace._3046_ ),
    .B1(\u_cpu.ALU.u_wallace._3047_ ),
    .Y(\u_cpu.ALU.u_wallace._3048_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8624_  (.A1_N(\u_cpu.ALU.u_wallace._2858_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3048_ ),
    .B1(\u_cpu.ALU.u_wallace._2850_ ),
    .B2(\u_cpu.ALU.u_wallace._2853_ ),
    .Y(\u_cpu.ALU.u_wallace._3049_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._8625_  (.A1(\u_cpu.ALU.u_wallace._2934_ ),
    .A2(\u_cpu.ALU.u_wallace._2939_ ),
    .B1_N(\u_cpu.ALU.u_wallace._2929_ ),
    .Y(\u_cpu.ALU.u_wallace._3050_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._8626_  (.A1(\u_cpu.ALU.u_wallace._3044_ ),
    .A2(\u_cpu.ALU.u_wallace._3045_ ),
    .B1(\u_cpu.ALU.u_wallace._3049_ ),
    .B2(\u_cpu.ALU.u_wallace._3050_ ),
    .X(\u_cpu.ALU.u_wallace._3051_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8627_  (.A(\u_cpu.ALU.u_wallace._2779_ ),
    .B(\u_cpu.ALU.u_wallace._1275_ ),
    .Y(\u_cpu.ALU.u_wallace._3052_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8628_  (.A(\u_cpu.ALU.u_wallace._4783_ ),
    .B(\u_cpu.ALU.u_wallace._0629_ ),
    .Y(\u_cpu.ALU.u_wallace._3054_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8629_  (.A1(\u_cpu.ALU.u_wallace._3052_ ),
    .A2(\u_cpu.ALU.u_wallace._3054_ ),
    .B1(\u_cpu.ALU.u_wallace._2877_ ),
    .Y(\u_cpu.ALU.u_wallace._3055_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8630_  (.A1(\u_cpu.ALU.u_wallace._4642_ ),
    .A2(\u_cpu.ALU.u_wallace._1102_ ),
    .B1(\u_cpu.ALU.u_wallace._1730_ ),
    .B2(\u_cpu.ALU.u_wallace._1771_ ),
    .X(\u_cpu.ALU.u_wallace._3056_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8631_  (.A(\u_cpu.ALU.u_wallace._4431_ ),
    .B(\u_cpu.ALU.u_wallace._4642_ ),
    .C(\u_cpu.ALU.u_wallace._1102_ ),
    .D(\u_cpu.ALU.u_wallace._1730_ ),
    .Y(\u_cpu.ALU.u_wallace._3057_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8632_  (.A(\u_cpu.ALU.SrcA[27] ),
    .X(\u_cpu.ALU.u_wallace._3058_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8633_  (.A(\u_cpu.ALU.u_wallace._3056_ ),
    .B(\u_cpu.ALU.u_wallace._3057_ ),
    .C(\u_cpu.ALU.u_wallace._0086_ ),
    .D(\u_cpu.ALU.u_wallace._3058_ ),
    .Y(\u_cpu.ALU.u_wallace._3059_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._8634_  (.A(\u_cpu.ALU.SrcA[27] ),
    .Y(\u_cpu.ALU.u_wallace._3060_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8635_  (.A1(\u_cpu.ALU.u_wallace._4551_ ),
    .A2(\u_cpu.ALU.u_wallace._0629_ ),
    .B1(\u_cpu.ALU.u_wallace._1535_ ),
    .B2(\u_cpu.ALU.u_wallace._1826_ ),
    .Y(\u_cpu.ALU.u_wallace._3061_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8636_  (.A(\u_cpu.ALU.u_wallace._1771_ ),
    .B(\u_cpu.ALU.u_wallace._4557_ ),
    .C(\u_cpu.ALU.u_wallace._1102_ ),
    .D(\u_cpu.ALU.u_wallace._1730_ ),
    .X(\u_cpu.ALU.u_wallace._3062_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8637_  (.A1(\u_cpu.ALU.u_wallace._4923_ ),
    .A2(\u_cpu.ALU.u_wallace._3060_ ),
    .B1(\u_cpu.ALU.u_wallace._3061_ ),
    .B2(\u_cpu.ALU.u_wallace._3062_ ),
    .Y(\u_cpu.ALU.u_wallace._3063_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8638_  (.A1(\u_cpu.ALU.u_wallace._2873_ ),
    .A2(\u_cpu.ALU.u_wallace._3055_ ),
    .B1(\u_cpu.ALU.u_wallace._3059_ ),
    .C1(\u_cpu.ALU.u_wallace._3063_ ),
    .X(\u_cpu.ALU.u_wallace._3065_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8639_  (.A1(\u_cpu.ALU.u_wallace._2866_ ),
    .A2(\u_cpu.ALU.u_wallace._2869_ ),
    .A3(\u_cpu.ALU.u_wallace._0086_ ),
    .B1(\u_cpu.ALU.u_wallace._2873_ ),
    .X(\u_cpu.ALU.u_wallace._3066_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8640_  (.A1(\u_cpu.ALU.u_wallace._3063_ ),
    .A2(\u_cpu.ALU.u_wallace._3059_ ),
    .B1(\u_cpu.ALU.u_wallace._3066_ ),
    .Y(\u_cpu.ALU.u_wallace._3067_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8641_  (.A(\u_cpu.ALU.u_wallace._0187_ ),
    .B(\u_cpu.ALU.u_wallace._0304_ ),
    .C(\u_cpu.ALU.u_wallace._2578_ ),
    .D(\u_cpu.ALU.SrcA[26] ),
    .Y(\u_cpu.ALU.u_wallace._3068_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8642_  (.A1(\u_cpu.ALU.u_wallace._1169_ ),
    .A2(\u_cpu.ALU.u_wallace._2578_ ),
    .B1(\u_cpu.ALU.SrcA[26] ),
    .B2(\u_cpu.ALU.u_wallace._1158_ ),
    .X(\u_cpu.ALU.u_wallace._3069_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8643_  (.A1_N(\u_cpu.ALU.u_wallace._3068_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3069_ ),
    .B1(\u_cpu.ALU.u_wallace._4678_ ),
    .B2(\u_cpu.ALU.u_wallace._2215_ ),
    .Y(\u_cpu.ALU.u_wallace._3070_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8644_  (.A(\u_cpu.ALU.u_wallace._3069_ ),
    .B(\u_cpu.ALU.u_wallace._2569_ ),
    .C(\u_cpu.ALU.u_wallace._0983_ ),
    .D(\u_cpu.ALU.u_wallace._3068_ ),
    .Y(\u_cpu.ALU.u_wallace._3071_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8645_  (.A(\u_cpu.ALU.u_wallace._3070_ ),
    .B(\u_cpu.ALU.u_wallace._3071_ ),
    .Y(\u_cpu.ALU.u_wallace._3072_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._8646_  (.A1(\u_cpu.ALU.u_wallace._3065_ ),
    .A2(\u_cpu.ALU.u_wallace._3067_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3072_ ),
    .Y(\u_cpu.ALU.u_wallace._3073_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU.u_wallace._8647_  (.A1_N(\u_cpu.ALU.u_wallace._3068_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3069_ ),
    .B1(\u_cpu.ALU.u_wallace._4678_ ),
    .B2(\u_cpu.ALU.u_wallace._2215_ ),
    .X(\u_cpu.ALU.u_wallace._3074_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8648_  (.A(\u_cpu.ALU.u_wallace._3069_ ),
    .B(\u_cpu.ALU.u_wallace._2569_ ),
    .C(\u_cpu.ALU.u_wallace._0983_ ),
    .D(\u_cpu.ALU.u_wallace._3068_ ),
    .X(\u_cpu.ALU.u_wallace._3076_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8649_  (.A1(\u_cpu.ALU.u_wallace._2873_ ),
    .A2(\u_cpu.ALU.u_wallace._3055_ ),
    .B1(\u_cpu.ALU.u_wallace._3059_ ),
    .C1(\u_cpu.ALU.u_wallace._3063_ ),
    .Y(\u_cpu.ALU.u_wallace._3077_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8650_  (.A1(\u_cpu.ALU.u_wallace._0884_ ),
    .A2(\u_cpu.ALU.u_wallace._3058_ ),
    .B1(\u_cpu.ALU.u_wallace._3056_ ),
    .B2(\u_cpu.ALU.u_wallace._3057_ ),
    .Y(\u_cpu.ALU.u_wallace._3078_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8651_  (.A(\u_cpu.ALU.u_wallace._2757_ ),
    .B(\u_cpu.ALU.u_wallace._3058_ ),
    .Y(\u_cpu.ALU.u_wallace._3079_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._8652_  (.A(\u_cpu.ALU.u_wallace._3079_ ),
    .B(\u_cpu.ALU.u_wallace._3061_ ),
    .C(\u_cpu.ALU.u_wallace._3062_ ),
    .Y(\u_cpu.ALU.u_wallace._3080_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._8653_  (.A1(\u_cpu.ALU.u_wallace._4934_ ),
    .A2(\u_cpu.ALU.u_wallace._2871_ ),
    .A3(\u_cpu.ALU.u_wallace._2872_ ),
    .B1(\u_cpu.ALU.u_wallace._2868_ ),
    .X(\u_cpu.ALU.u_wallace._3081_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8654_  (.A1(\u_cpu.ALU.u_wallace._3078_ ),
    .A2(\u_cpu.ALU.u_wallace._3080_ ),
    .B1(\u_cpu.ALU.u_wallace._3081_ ),
    .Y(\u_cpu.ALU.u_wallace._3082_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8655_  (.A1(\u_cpu.ALU.u_wallace._3074_ ),
    .A2(\u_cpu.ALU.u_wallace._3076_ ),
    .B1(\u_cpu.ALU.u_wallace._3077_ ),
    .C1(\u_cpu.ALU.u_wallace._3082_ ),
    .Y(\u_cpu.ALU.u_wallace._3083_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8656_  (.A1(\u_cpu.ALU.u_wallace._2897_ ),
    .A2(\u_cpu.ALU.u_wallace._2892_ ),
    .B1(\u_cpu.ALU.u_wallace._3073_ ),
    .B2(\u_cpu.ALU.u_wallace._3083_ ),
    .Y(\u_cpu.ALU.u_wallace._3084_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8657_  (.A1(\u_cpu.ALU.u_wallace._2883_ ),
    .A2(\u_cpu.ALU.u_wallace._2882_ ),
    .A3(\u_cpu.ALU.u_wallace._0983_ ),
    .B1(\u_cpu.ALU.u_wallace._2888_ ),
    .X(\u_cpu.ALU.u_wallace._3085_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8658_  (.A1(\u_cpu.ALU.u_wallace._2187_ ),
    .A2(\u_cpu.ALU.u_wallace._1742_ ),
    .B1(\u_cpu.ALU.u_wallace._2002_ ),
    .B2(\u_cpu.ALU.u_wallace._2155_ ),
    .X(\u_cpu.ALU.u_wallace._3087_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8659_  (.A(\u_cpu.ALU.u_wallace._1543_ ),
    .X(\u_cpu.ALU.u_wallace._3088_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8660_  (.A(\u_cpu.ALU.u_wallace._1476_ ),
    .B(\u_cpu.ALU.u_wallace._2187_ ),
    .C(\u_cpu.ALU.u_wallace._1742_ ),
    .D(\u_cpu.ALU.u_wallace._2002_ ),
    .Y(\u_cpu.ALU.u_wallace._3089_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8661_  (.A(\u_cpu.ALU.u_wallace._3087_ ),
    .B(\u_cpu.ALU.u_wallace._3088_ ),
    .C(\u_cpu.ALU.u_wallace._4542_ ),
    .D(\u_cpu.ALU.u_wallace._3089_ ),
    .Y(\u_cpu.ALU.u_wallace._3090_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8662_  (.A1(\u_cpu.ALU.u_wallace._4542_ ),
    .A2(\u_cpu.ALU.u_wallace._3088_ ),
    .B1(\u_cpu.ALU.u_wallace._3089_ ),
    .B2(\u_cpu.ALU.u_wallace._3087_ ),
    .X(\u_cpu.ALU.u_wallace._3091_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8663_  (.A(\u_cpu.ALU.u_wallace._3085_ ),
    .B(\u_cpu.ALU.u_wallace._3090_ ),
    .C(\u_cpu.ALU.u_wallace._3091_ ),
    .Y(\u_cpu.ALU.u_wallace._3092_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.ALU.u_wallace._8664_  (.A1_N(\u_cpu.ALU.u_wallace._4539_ ),
    .A2_N(\u_cpu.ALU.u_wallace._1271_ ),
    .B1(\u_cpu.ALU.u_wallace._3089_ ),
    .B2(\u_cpu.ALU.u_wallace._3087_ ),
    .Y(\u_cpu.ALU.u_wallace._3093_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8665_  (.A1(\u_cpu.ALU.u_wallace._1508_ ),
    .A2(\u_cpu.ALU.u_wallace._1742_ ),
    .B1(\u_cpu.ALU.u_wallace._2882_ ),
    .B2(\u_cpu.ALU.u_wallace._1476_ ),
    .Y(\u_cpu.ALU.u_wallace._3094_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8666_  (.A(\u_cpu.ALU.u_wallace._2604_ ),
    .B(\u_cpu.ALU.u_wallace._1275_ ),
    .Y(\u_cpu.ALU.u_wallace._3095_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8667_  (.A(\u_cpu.ALU.u_wallace._2155_ ),
    .B(\u_cpu.ALU.u_wallace._2187_ ),
    .C(\u_cpu.ALU.u_wallace._1742_ ),
    .D(\u_cpu.ALU.u_wallace._2000_ ),
    .X(\u_cpu.ALU.u_wallace._3096_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._8668_  (.A(\u_cpu.ALU.u_wallace._3094_ ),
    .B(\u_cpu.ALU.u_wallace._3095_ ),
    .C(\u_cpu.ALU.u_wallace._3096_ ),
    .Y(\u_cpu.ALU.u_wallace._3098_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._8669_  (.A1(\u_cpu.ALU.u_wallace._2887_ ),
    .A2(\u_cpu.ALU.u_wallace._2886_ ),
    .B1(\u_cpu.ALU.u_wallace._3093_ ),
    .B2(\u_cpu.ALU.u_wallace._3098_ ),
    .C1(\u_cpu.ALU.u_wallace._2884_ ),
    .Y(\u_cpu.ALU.u_wallace._3099_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._8670_  (.A1(\u_cpu.ALU.u_wallace._2284_ ),
    .A2(\u_cpu.ALU.u_wallace._1096_ ),
    .A3(\u_cpu.ALU.u_wallace._2902_ ),
    .B1(\u_cpu.ALU.u_wallace._2906_ ),
    .X(\u_cpu.ALU.u_wallace._3100_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8671_  (.A1(\u_cpu.ALU.u_wallace._3092_ ),
    .A2(\u_cpu.ALU.u_wallace._3099_ ),
    .B1(\u_cpu.ALU.u_wallace._3100_ ),
    .Y(\u_cpu.ALU.u_wallace._3101_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8672_  (.A(\u_cpu.ALU.u_wallace._3099_ ),
    .B(\u_cpu.ALU.u_wallace._3100_ ),
    .C(\u_cpu.ALU.u_wallace._3092_ ),
    .X(\u_cpu.ALU.u_wallace._3102_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8673_  (.A1(\u_cpu.ALU.u_wallace._2881_ ),
    .A2(\u_cpu.ALU.u_wallace._2891_ ),
    .B1(\u_cpu.ALU.u_wallace._2875_ ),
    .Y(\u_cpu.ALU.u_wallace._3103_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8674_  (.A(\u_cpu.ALU.u_wallace._3073_ ),
    .B(\u_cpu.ALU.u_wallace._3083_ ),
    .C(\u_cpu.ALU.u_wallace._3103_ ),
    .Y(\u_cpu.ALU.u_wallace._3104_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8675_  (.A1(\u_cpu.ALU.u_wallace._3101_ ),
    .A2(\u_cpu.ALU.u_wallace._3102_ ),
    .B1(\u_cpu.ALU.u_wallace._3104_ ),
    .Y(\u_cpu.ALU.u_wallace._3105_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._8676_  (.A1(\u_cpu.ALU.u_wallace._2899_ ),
    .A2(\u_cpu.ALU.u_wallace._2896_ ),
    .A3(\u_cpu.ALU.u_wallace._2898_ ),
    .B1(\u_cpu.ALU.u_wallace._2923_ ),
    .Y(\u_cpu.ALU.u_wallace._3106_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8677_  (.A(\u_cpu.ALU.u_wallace._2905_ ),
    .B(\u_cpu.ALU.u_wallace._2907_ ),
    .C(\u_cpu.ALU.u_wallace._2917_ ),
    .X(\u_cpu.ALU.u_wallace._3107_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8678_  (.A1(\u_cpu.ALU.u_wallace._2903_ ),
    .A2(\u_cpu.ALU.u_wallace._3107_ ),
    .B1(\u_cpu.ALU.u_wallace._3092_ ),
    .C1(\u_cpu.ALU.u_wallace._3099_ ),
    .X(\u_cpu.ALU.u_wallace._3109_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8679_  (.A1(\u_cpu.ALU.u_wallace._2905_ ),
    .A2(\u_cpu.ALU.u_wallace._2907_ ),
    .A3(\u_cpu.ALU.u_wallace._2917_ ),
    .B1(\u_cpu.ALU.u_wallace._2903_ ),
    .X(\u_cpu.ALU.u_wallace._3110_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8680_  (.A1(\u_cpu.ALU.u_wallace._3092_ ),
    .A2(\u_cpu.ALU.u_wallace._3099_ ),
    .B1(\u_cpu.ALU.u_wallace._3110_ ),
    .Y(\u_cpu.ALU.u_wallace._3111_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8681_  (.A(\u_cpu.ALU.u_wallace._3070_ ),
    .B(\u_cpu.ALU.u_wallace._3071_ ),
    .C(\u_cpu.ALU.u_wallace._3077_ ),
    .D(\u_cpu.ALU.u_wallace._3082_ ),
    .Y(\u_cpu.ALU.u_wallace._3112_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8682_  (.A1(\u_cpu.ALU.u_wallace._3074_ ),
    .A2(\u_cpu.ALU.u_wallace._3076_ ),
    .B1(\u_cpu.ALU.u_wallace._3065_ ),
    .B2(\u_cpu.ALU.u_wallace._3067_ ),
    .Y(\u_cpu.ALU.u_wallace._3113_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._8683_  (.A1(\u_cpu.ALU.u_wallace._2874_ ),
    .A2(\u_cpu.ALU.u_wallace._2870_ ),
    .A3(\u_cpu.ALU.u_wallace._2880_ ),
    .B1(\u_cpu.ALU.u_wallace._2881_ ),
    .B2(\u_cpu.ALU.u_wallace._2891_ ),
    .X(\u_cpu.ALU.u_wallace._3114_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8684_  (.A1(\u_cpu.ALU.u_wallace._3112_ ),
    .A2(\u_cpu.ALU.u_wallace._3113_ ),
    .B1(\u_cpu.ALU.u_wallace._3114_ ),
    .Y(\u_cpu.ALU.u_wallace._3115_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8685_  (.A1(\u_cpu.ALU.u_wallace._3109_ ),
    .A2(\u_cpu.ALU.u_wallace._3111_ ),
    .B1(\u_cpu.ALU.u_wallace._3084_ ),
    .B2(\u_cpu.ALU.u_wallace._3115_ ),
    .Y(\u_cpu.ALU.u_wallace._3116_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._8686_  (.A1(\u_cpu.ALU.u_wallace._3084_ ),
    .A2(\u_cpu.ALU.u_wallace._3105_ ),
    .B1(\u_cpu.ALU.u_wallace._2936_ ),
    .B2(\u_cpu.ALU.u_wallace._3106_ ),
    .C1(\u_cpu.ALU.u_wallace._3116_ ),
    .X(\u_cpu.ALU.u_wallace._3117_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8687_  (.A(\u_cpu.ALU.u_wallace._2925_ ),
    .B(\u_cpu.ALU.u_wallace._2926_ ),
    .Y(\u_cpu.ALU.u_wallace._3118_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8688_  (.A1(\u_cpu.ALU.u_wallace._3118_ ),
    .A2(\u_cpu.ALU.u_wallace._2901_ ),
    .B1(\u_cpu.ALU.u_wallace._2936_ ),
    .Y(\u_cpu.ALU.u_wallace._3120_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8689_  (.A1(\u_cpu.ALU.u_wallace._3101_ ),
    .A2(\u_cpu.ALU.u_wallace._3102_ ),
    .B1(\u_cpu.ALU.u_wallace._3084_ ),
    .B2(\u_cpu.ALU.u_wallace._3115_ ),
    .Y(\u_cpu.ALU.u_wallace._3121_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8690_  (.A(\u_cpu.ALU.u_wallace._3114_ ),
    .B(\u_cpu.ALU.u_wallace._3112_ ),
    .C(\u_cpu.ALU.u_wallace._3113_ ),
    .Y(\u_cpu.ALU.u_wallace._3122_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8691_  (.A1(\u_cpu.ALU.u_wallace._3109_ ),
    .A2(\u_cpu.ALU.u_wallace._3111_ ),
    .B1(\u_cpu.ALU.u_wallace._3122_ ),
    .C1(\u_cpu.ALU.u_wallace._3104_ ),
    .Y(\u_cpu.ALU.u_wallace._3123_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8692_  (.A(\u_cpu.ALU.u_wallace._3120_ ),
    .B(\u_cpu.ALU.u_wallace._3121_ ),
    .C(\u_cpu.ALU.u_wallace._3123_ ),
    .Y(\u_cpu.ALU.u_wallace._3124_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8693_  (.A1(\u_cpu.ALU.u_wallace._4599_ ),
    .A2(\u_cpu.ALU.u_wallace._0815_ ),
    .B1(\u_cpu.ALU.u_wallace._1101_ ),
    .B2(\u_cpu.ALU.u_wallace._4717_ ),
    .Y(\u_cpu.ALU.u_wallace._3125_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8694_  (.A(\u_cpu.ALU.u_wallace._4594_ ),
    .B(\u_cpu.ALU.u_wallace._4595_ ),
    .C(\u_cpu.ALU.u_wallace._0802_ ),
    .D(\u_cpu.ALU.u_wallace._1090_ ),
    .X(\u_cpu.ALU.u_wallace._3126_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8695_  (.A1(\u_cpu.ALU.u_wallace._4602_ ),
    .A2(\u_cpu.ALU.u_wallace._0635_ ),
    .B1(\u_cpu.ALU.u_wallace._3125_ ),
    .B2(\u_cpu.ALU.u_wallace._3126_ ),
    .Y(\u_cpu.ALU.u_wallace._3127_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8696_  (.A1(\u_cpu.ALU.u_wallace._4302_ ),
    .A2(\u_cpu.ALU.u_wallace._0802_ ),
    .B1(\u_cpu.ALU.u_wallace._1101_ ),
    .B2(\u_cpu.ALU.u_wallace._4018_ ),
    .X(\u_cpu.ALU.u_wallace._3128_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8697_  (.A(\u_cpu.ALU.u_wallace._4717_ ),
    .B(\u_cpu.ALU.u_wallace._4599_ ),
    .C(\u_cpu.ALU.u_wallace._0815_ ),
    .D(\u_cpu.ALU.u_wallace._1101_ ),
    .Y(\u_cpu.ALU.u_wallace._3129_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8698_  (.A(\u_cpu.ALU.u_wallace._3128_ ),
    .B(\u_cpu.ALU.u_wallace._3129_ ),
    .C(\u_cpu.ALU.u_wallace._4610_ ),
    .D(\u_cpu.ALU.u_wallace._1286_ ),
    .Y(\u_cpu.ALU.u_wallace._3131_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8699_  (.A1(\u_cpu.ALU.u_wallace._2833_ ),
    .A2(\u_cpu.ALU.u_wallace._2829_ ),
    .B1(\u_cpu.ALU.u_wallace._2826_ ),
    .Y(\u_cpu.ALU.u_wallace._3132_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8700_  (.A(\u_cpu.ALU.u_wallace._4732_ ),
    .B(\u_cpu.ALU.u_wallace._4842_ ),
    .C(\u_cpu.ALU.u_wallace._0826_ ),
    .D(\u_cpu.ALU.u_wallace._1075_ ),
    .Y(\u_cpu.ALU.u_wallace._3133_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8701_  (.A1(\u_cpu.ALU.u_wallace._4842_ ),
    .A2(\u_cpu.ALU.u_wallace._0826_ ),
    .B1(\u_cpu.ALU.u_wallace._1075_ ),
    .B2(\u_cpu.ALU.u_wallace._4732_ ),
    .X(\u_cpu.ALU.u_wallace._3134_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8702_  (.A1(\u_cpu.ALU.u_wallace._0037_ ),
    .A2(\u_cpu.ALU.u_wallace._1323_ ),
    .B1(\u_cpu.ALU.u_wallace._3133_ ),
    .C1(\u_cpu.ALU.u_wallace._3134_ ),
    .Y(\u_cpu.ALU.u_wallace._3135_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8703_  (.A(\u_cpu.ALU.u_wallace._4840_ ),
    .B(\u_cpu.ALU.u_wallace._4842_ ),
    .C(\u_cpu.ALU.u_wallace._0325_ ),
    .D(\u_cpu.ALU.u_wallace._0850_ ),
    .X(\u_cpu.ALU.u_wallace._3136_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8704_  (.A1(\u_cpu.ALU.u_wallace._4842_ ),
    .A2(\u_cpu.ALU.u_wallace._0325_ ),
    .B1(\u_cpu.ALU.u_wallace._1075_ ),
    .B2(\u_cpu.ALU.u_wallace._4840_ ),
    .Y(\u_cpu.ALU.u_wallace._3137_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8705_  (.A(\u_cpu.ALU.u_wallace._0363_ ),
    .B(\u_cpu.ALU.u_wallace._0320_ ),
    .Y(\u_cpu.ALU.u_wallace._3138_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._8706_  (.A1(\u_cpu.ALU.u_wallace._3136_ ),
    .A2(\u_cpu.ALU.u_wallace._3137_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3138_ ),
    .Y(\u_cpu.ALU.u_wallace._3139_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._8707_  (.A1(\u_cpu.ALU.u_wallace._3127_ ),
    .A2(\u_cpu.ALU.u_wallace._3131_ ),
    .A3(\u_cpu.ALU.u_wallace._3132_ ),
    .B1(\u_cpu.ALU.u_wallace._3135_ ),
    .B2(\u_cpu.ALU.u_wallace._3139_ ),
    .X(\u_cpu.ALU.u_wallace._3140_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8708_  (.A1(\u_cpu.ALU.u_wallace._3127_ ),
    .A2(\u_cpu.ALU.u_wallace._3131_ ),
    .B1(\u_cpu.ALU.u_wallace._3132_ ),
    .Y(\u_cpu.ALU.u_wallace._3142_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8709_  (.A1(\u_cpu.ALU.u_wallace._2914_ ),
    .A2(\u_cpu.ALU.u_wallace._2910_ ),
    .B1(\u_cpu.ALU.u_wallace._2920_ ),
    .Y(\u_cpu.ALU.u_wallace._3143_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8710_  (.A(\u_cpu.ALU.u_wallace._4599_ ),
    .B(\u_cpu.ALU.u_wallace._1286_ ),
    .Y(\u_cpu.ALU.u_wallace._3144_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8711_  (.A(\u_cpu.ALU.u_wallace._4717_ ),
    .B(\u_cpu.ALU.u_wallace._0815_ ),
    .Y(\u_cpu.ALU.u_wallace._3145_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8712_  (.A1(\u_cpu.ALU.u_wallace._3144_ ),
    .A2(\u_cpu.ALU.u_wallace._3145_ ),
    .B1(\u_cpu.ALU.u_wallace._2833_ ),
    .Y(\u_cpu.ALU.u_wallace._3146_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8713_  (.A1(\u_cpu.ALU.u_wallace._2828_ ),
    .A2(\u_cpu.ALU.u_wallace._3146_ ),
    .B1(\u_cpu.ALU.u_wallace._3131_ ),
    .C1(\u_cpu.ALU.u_wallace._3127_ ),
    .X(\u_cpu.ALU.u_wallace._3147_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._8714_  (.A(\u_cpu.ALU.u_wallace._3139_ ),
    .B(\u_cpu.ALU.u_wallace._3135_ ),
    .X(\u_cpu.ALU.u_wallace._3148_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8715_  (.A1(\u_cpu.ALU.u_wallace._3147_ ),
    .A2(\u_cpu.ALU.u_wallace._3142_ ),
    .B1(\u_cpu.ALU.u_wallace._3148_ ),
    .Y(\u_cpu.ALU.u_wallace._3149_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8716_  (.A1(\u_cpu.ALU.u_wallace._3140_ ),
    .A2(\u_cpu.ALU.u_wallace._3142_ ),
    .B1(\u_cpu.ALU.u_wallace._3143_ ),
    .C1(\u_cpu.ALU.u_wallace._3149_ ),
    .Y(\u_cpu.ALU.u_wallace._3150_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._8717_  (.A1(\u_cpu.ALU.u_wallace._2914_ ),
    .A2(\u_cpu.ALU.u_wallace._2910_ ),
    .B1(\u_cpu.ALU.u_wallace._2920_ ),
    .X(\u_cpu.ALU.u_wallace._3151_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8718_  (.A(\u_cpu.ALU.u_wallace._3139_ ),
    .B(\u_cpu.ALU.u_wallace._3135_ ),
    .Y(\u_cpu.ALU.u_wallace._3153_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8719_  (.A1(\u_cpu.ALU.u_wallace._3147_ ),
    .A2(\u_cpu.ALU.u_wallace._3142_ ),
    .B1(\u_cpu.ALU.u_wallace._3153_ ),
    .Y(\u_cpu.ALU.u_wallace._3154_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8720_  (.A1(\u_cpu.ALU.u_wallace._2828_ ),
    .A2(\u_cpu.ALU.u_wallace._3146_ ),
    .B1(\u_cpu.ALU.u_wallace._3131_ ),
    .C1(\u_cpu.ALU.u_wallace._3127_ ),
    .Y(\u_cpu.ALU.u_wallace._3155_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8721_  (.A1(\u_cpu.ALU.u_wallace._3127_ ),
    .A2(\u_cpu.ALU.u_wallace._3131_ ),
    .B1(\u_cpu.ALU.u_wallace._3132_ ),
    .X(\u_cpu.ALU.u_wallace._3156_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8722_  (.A(\u_cpu.ALU.u_wallace._3148_ ),
    .B(\u_cpu.ALU.u_wallace._3155_ ),
    .C(\u_cpu.ALU.u_wallace._3156_ ),
    .Y(\u_cpu.ALU.u_wallace._3157_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8723_  (.A(\u_cpu.ALU.u_wallace._3151_ ),
    .B(\u_cpu.ALU.u_wallace._3154_ ),
    .C(\u_cpu.ALU.u_wallace._3157_ ),
    .Y(\u_cpu.ALU.u_wallace._3158_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._8724_  (.A1(\u_cpu.ALU.u_wallace._2831_ ),
    .A2(\u_cpu.ALU.u_wallace._2942_ ),
    .B1(\u_cpu.ALU.u_wallace._3158_ ),
    .X(\u_cpu.ALU.u_wallace._3159_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8725_  (.A1(\u_cpu.ALU.u_wallace._1578_ ),
    .A2(\u_cpu.ALU.u_wallace._0117_ ),
    .B1(\u_cpu.ALU.u_wallace._2837_ ),
    .B2(\u_cpu.ALU.u_wallace._2838_ ),
    .X(\u_cpu.ALU.u_wallace._3160_ ));
 sky130_fd_sc_hd__or4_2 \u_cpu.ALU.u_wallace._8726_  (.A(\u_cpu.ALU.u_wallace._0458_ ),
    .B(\u_cpu.ALU.u_wallace._0124_ ),
    .C(\u_cpu.ALU.u_wallace._2841_ ),
    .D(\u_cpu.ALU.u_wallace._2842_ ),
    .X(\u_cpu.ALU.u_wallace._3161_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8727_  (.A1(\u_cpu.ALU.u_wallace._2836_ ),
    .A2(\u_cpu.ALU.u_wallace._3160_ ),
    .A3(\u_cpu.ALU.u_wallace._3161_ ),
    .B1(\u_cpu.ALU.u_wallace._2831_ ),
    .X(\u_cpu.ALU.u_wallace._3162_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8728_  (.A1(\u_cpu.ALU.u_wallace._3158_ ),
    .A2(\u_cpu.ALU.u_wallace._3150_ ),
    .B1(\u_cpu.ALU.u_wallace._3162_ ),
    .Y(\u_cpu.ALU.u_wallace._3164_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8729_  (.A1(\u_cpu.ALU.u_wallace._3150_ ),
    .A2(\u_cpu.ALU.u_wallace._3159_ ),
    .B1(\u_cpu.ALU.u_wallace._3164_ ),
    .Y(\u_cpu.ALU.u_wallace._3165_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8730_  (.A(\u_cpu.ALU.u_wallace._3124_ ),
    .B(\u_cpu.ALU.u_wallace._3165_ ),
    .Y(\u_cpu.ALU.u_wallace._3166_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._8731_  (.A1(\u_cpu.ALU.u_wallace._3084_ ),
    .A2(\u_cpu.ALU.u_wallace._3105_ ),
    .B1(\u_cpu.ALU.u_wallace._2936_ ),
    .B2(\u_cpu.ALU.u_wallace._3106_ ),
    .C1(\u_cpu.ALU.u_wallace._3116_ ),
    .Y(\u_cpu.ALU.u_wallace._3167_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8732_  (.A1(\u_cpu.ALU.u_wallace._2831_ ),
    .A2(\u_cpu.ALU.u_wallace._2942_ ),
    .B1(\u_cpu.ALU.u_wallace._3158_ ),
    .C1(\u_cpu.ALU.u_wallace._3150_ ),
    .Y(\u_cpu.ALU.u_wallace._3168_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._8733_  (.A(\u_cpu.ALU.u_wallace._3168_ ),
    .Y(\u_cpu.ALU.u_wallace._3169_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8734_  (.A1_N(\u_cpu.ALU.u_wallace._3167_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3124_ ),
    .B1(\u_cpu.ALU.u_wallace._3164_ ),
    .B2(\u_cpu.ALU.u_wallace._3169_ ),
    .Y(\u_cpu.ALU.u_wallace._3170_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8735_  (.A1(\u_cpu.ALU.u_wallace._3117_ ),
    .A2(\u_cpu.ALU.u_wallace._3166_ ),
    .B1(\u_cpu.ALU.u_wallace._3170_ ),
    .Y(\u_cpu.ALU.u_wallace._3171_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8736_  (.A(\u_cpu.ALU.u_wallace._4669_ ),
    .B(\u_cpu.ALU.u_wallace._4698_ ),
    .C(\u_cpu.ALU.u_wallace._0958_ ),
    .D(\u_cpu.ALU.u_wallace._1208_ ),
    .X(\u_cpu.ALU.u_wallace._3172_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8737_  (.A(\u_cpu.ALU.u_wallace._4452_ ),
    .B(\u_cpu.ALU.u_wallace._1386_ ),
    .Y(\u_cpu.ALU.u_wallace._3173_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8738_  (.A1(\u_cpu.ALU.u_wallace._4669_ ),
    .A2(\u_cpu.ALU.u_wallace._0958_ ),
    .B1(\u_cpu.ALU.u_wallace._1208_ ),
    .B2(\u_cpu.ALU.u_wallace._2801_ ),
    .Y(\u_cpu.ALU.u_wallace._3175_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8739_  (.A(\u_cpu.ALU.u_wallace._3173_ ),
    .B(\u_cpu.ALU.u_wallace._3175_ ),
    .Y(\u_cpu.ALU.u_wallace._3176_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8740_  (.A1(\u_cpu.ALU.u_wallace._4783_ ),
    .A2(\u_cpu.ALU.u_wallace._2050_ ),
    .B1(\u_cpu.ALU.u_wallace._1175_ ),
    .B2(\u_cpu.ALU.u_wallace._4660_ ),
    .X(\u_cpu.ALU.u_wallace._3177_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8741_  (.A(\u_cpu.ALU.u_wallace._4669_ ),
    .B(\u_cpu.ALU.u_wallace._4783_ ),
    .C(\u_cpu.ALU.u_wallace._2050_ ),
    .D(\u_cpu.ALU.u_wallace._1208_ ),
    .Y(\u_cpu.ALU.u_wallace._3178_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8742_  (.A(\u_cpu.ALU.u_wallace._3177_ ),
    .B(\u_cpu.ALU.u_wallace._3178_ ),
    .C(\u_cpu.ALU.u_wallace._4698_ ),
    .D(\u_cpu.ALU.u_wallace._1615_ ),
    .Y(\u_cpu.ALU.u_wallace._3179_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8743_  (.A1(\u_cpu.ALU.u_wallace._4783_ ),
    .A2(\u_cpu.ALU.u_wallace._2050_ ),
    .B1(\u_cpu.ALU.u_wallace._1208_ ),
    .B2(\u_cpu.ALU.u_wallace._4660_ ),
    .Y(\u_cpu.ALU.u_wallace._3180_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8744_  (.A(\u_cpu.ALU.u_wallace._4660_ ),
    .B(\u_cpu.ALU.u_wallace._4567_ ),
    .C(\u_cpu.ALU.u_wallace._1387_ ),
    .D(\u_cpu.ALU.u_wallace._1175_ ),
    .X(\u_cpu.ALU.u_wallace._3181_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8745_  (.A1(\u_cpu.ALU.u_wallace._0203_ ),
    .A2(\u_cpu.ALU.u_wallace._2053_ ),
    .B1(\u_cpu.ALU.u_wallace._3180_ ),
    .B2(\u_cpu.ALU.u_wallace._3181_ ),
    .Y(\u_cpu.ALU.u_wallace._3182_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8746_  (.A1(\u_cpu.ALU.u_wallace._3172_ ),
    .A2(\u_cpu.ALU.u_wallace._3176_ ),
    .B1(\u_cpu.ALU.u_wallace._3179_ ),
    .C1(\u_cpu.ALU.u_wallace._3182_ ),
    .X(\u_cpu.ALU.u_wallace._3183_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8747_  (.A1(\u_cpu.ALU.u_wallace._3173_ ),
    .A2(\u_cpu.ALU.u_wallace._3175_ ),
    .B1(\u_cpu.ALU.u_wallace._2784_ ),
    .Y(\u_cpu.ALU.u_wallace._3184_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8748_  (.A1(\u_cpu.ALU.u_wallace._3179_ ),
    .A2(\u_cpu.ALU.u_wallace._3182_ ),
    .B1(\u_cpu.ALU.u_wallace._3184_ ),
    .Y(\u_cpu.ALU.u_wallace._3186_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8749_  (.A(\u_cpu.ALU.u_wallace._4452_ ),
    .B(\u_cpu.ALU.u_wallace._1322_ ),
    .C(\u_cpu.ALU.SrcB[21] ),
    .D(\u_cpu.ALU.SrcB[22] ),
    .X(\u_cpu.ALU.u_wallace._3187_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8750_  (.A1(\u_cpu.ALU.u_wallace._4452_ ),
    .A2(\u_cpu.ALU.SrcB[21] ),
    .B1(\u_cpu.ALU.SrcB[22] ),
    .B2(\u_cpu.ALU.u_wallace._1136_ ),
    .Y(\u_cpu.ALU.u_wallace._3188_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._8751_  (.A1(\u_cpu.ALU.u_wallace._3183_ ),
    .A2(\u_cpu.ALU.u_wallace._3186_ ),
    .B1(\u_cpu.ALU.u_wallace._3187_ ),
    .B2(\u_cpu.ALU.u_wallace._3188_ ),
    .X(\u_cpu.ALU.u_wallace._3189_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU.u_wallace._8752_  (.A(\u_cpu.ALU.u_wallace._3187_ ),
    .B(\u_cpu.ALU.u_wallace._3188_ ),
    .X(\u_cpu.ALU.u_wallace._3190_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8753_  (.A1(\u_cpu.ALU.u_wallace._3184_ ),
    .A2(\u_cpu.ALU.u_wallace._3179_ ),
    .A3(\u_cpu.ALU.u_wallace._3182_ ),
    .B1(\u_cpu.ALU.u_wallace._3190_ ),
    .X(\u_cpu.ALU.u_wallace._3191_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8754_  (.A(\u_cpu.ALU.u_wallace._3186_ ),
    .B(\u_cpu.ALU.u_wallace._3191_ ),
    .Y(\u_cpu.ALU.u_wallace._3192_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8755_  (.A1(\u_cpu.ALU.u_wallace._0188_ ),
    .A2(\u_cpu.ALU.u_wallace._0546_ ),
    .B1(\u_cpu.ALU.u_wallace._0279_ ),
    .B2(\u_cpu.ALU.u_wallace._4917_ ),
    .Y(\u_cpu.ALU.u_wallace._3193_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8756_  (.A(\u_cpu.ALU.u_wallace._4785_ ),
    .B(\u_cpu.ALU.u_wallace._4907_ ),
    .C(\u_cpu.ALU.u_wallace._0730_ ),
    .D(\u_cpu.ALU.u_wallace._0732_ ),
    .X(\u_cpu.ALU.u_wallace._3194_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8757_  (.A1(\u_cpu.ALU.u_wallace._0169_ ),
    .A2(\u_cpu.ALU.u_wallace._0941_ ),
    .B1(\u_cpu.ALU.u_wallace._3193_ ),
    .B2(\u_cpu.ALU.u_wallace._3194_ ),
    .Y(\u_cpu.ALU.u_wallace._3195_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8758_  (.A1(\u_cpu.ALU.u_wallace._4921_ ),
    .A2(\u_cpu.ALU.u_wallace._0730_ ),
    .B1(\u_cpu.ALU.u_wallace._0547_ ),
    .B2(\u_cpu.ALU.u_wallace._4787_ ),
    .X(\u_cpu.ALU.u_wallace._3197_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8759_  (.A(\u_cpu.ALU.u_wallace._4917_ ),
    .B(\u_cpu.ALU.u_wallace._0188_ ),
    .C(\u_cpu.ALU.u_wallace._0546_ ),
    .D(\u_cpu.ALU.u_wallace._0547_ ),
    .Y(\u_cpu.ALU.u_wallace._3198_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8760_  (.A(\u_cpu.ALU.u_wallace._3197_ ),
    .B(\u_cpu.ALU.u_wallace._3198_ ),
    .C(\u_cpu.ALU.u_wallace._4798_ ),
    .D(\u_cpu.ALU.u_wallace._0735_ ),
    .Y(\u_cpu.ALU.u_wallace._3199_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8761_  (.A1(\u_cpu.ALU.u_wallace._2839_ ),
    .A2(\u_cpu.ALU.u_wallace._2841_ ),
    .B1(\u_cpu.ALU.u_wallace._2838_ ),
    .Y(\u_cpu.ALU.u_wallace._3200_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8762_  (.A1(\u_cpu.ALU.u_wallace._3195_ ),
    .A2(\u_cpu.ALU.u_wallace._3199_ ),
    .B1(\u_cpu.ALU.u_wallace._3200_ ),
    .Y(\u_cpu.ALU.u_wallace._3201_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8763_  (.A(\u_cpu.ALU.u_wallace._2839_ ),
    .B(\u_cpu.ALU.u_wallace._2841_ ),
    .Y(\u_cpu.ALU.u_wallace._3202_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8764_  (.A1(\u_cpu.ALU.u_wallace._2842_ ),
    .A2(\u_cpu.ALU.u_wallace._3202_ ),
    .B1(\u_cpu.ALU.u_wallace._3199_ ),
    .C1(\u_cpu.ALU.u_wallace._3195_ ),
    .X(\u_cpu.ALU.u_wallace._3203_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8765_  (.A(\u_cpu.ALU.u_wallace._0551_ ),
    .X(\u_cpu.ALU.u_wallace._3204_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8766_  (.A(\u_cpu.ALU.u_wallace._4798_ ),
    .B(\u_cpu.ALU.u_wallace._0475_ ),
    .C(\u_cpu.ALU.u_wallace._0121_ ),
    .D(\u_cpu.ALU.u_wallace._0279_ ),
    .X(\u_cpu.ALU.u_wallace._3205_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._8767_  (.A1(\u_cpu.ALU.u_wallace._2760_ ),
    .A2(\u_cpu.ALU.u_wallace._3204_ ),
    .A3(\u_cpu.ALU.u_wallace._0847_ ),
    .B1(\u_cpu.ALU.u_wallace._3205_ ),
    .Y(\u_cpu.ALU.u_wallace._3206_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8768_  (.A1(\u_cpu.ALU.u_wallace._3201_ ),
    .A2(\u_cpu.ALU.u_wallace._3203_ ),
    .B1(\u_cpu.ALU.u_wallace._3206_ ),
    .Y(\u_cpu.ALU.u_wallace._3208_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8769_  (.A1(\u_cpu.ALU.u_wallace._3195_ ),
    .A2(\u_cpu.ALU.u_wallace._3199_ ),
    .B1(\u_cpu.ALU.u_wallace._3200_ ),
    .X(\u_cpu.ALU.u_wallace._3209_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8770_  (.A1(\u_cpu.ALU.u_wallace._2842_ ),
    .A2(\u_cpu.ALU.u_wallace._3202_ ),
    .B1(\u_cpu.ALU.u_wallace._3199_ ),
    .C1(\u_cpu.ALU.u_wallace._3195_ ),
    .Y(\u_cpu.ALU.u_wallace._3210_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8771_  (.A1(\u_cpu.ALU.u_wallace._2760_ ),
    .A2(\u_cpu.ALU.u_wallace._3204_ ),
    .A3(\u_cpu.ALU.u_wallace._0847_ ),
    .B1(\u_cpu.ALU.u_wallace._3205_ ),
    .X(\u_cpu.ALU.u_wallace._3211_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8772_  (.A(\u_cpu.ALU.u_wallace._3209_ ),
    .B(\u_cpu.ALU.u_wallace._3210_ ),
    .C(\u_cpu.ALU.u_wallace._3211_ ),
    .Y(\u_cpu.ALU.u_wallace._3212_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8773_  (.A1(\u_cpu.ALU.u_wallace._2769_ ),
    .A2(\u_cpu.ALU.u_wallace._2766_ ),
    .B1(\u_cpu.ALU.u_wallace._2772_ ),
    .Y(\u_cpu.ALU.u_wallace._3213_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8774_  (.A1(\u_cpu.ALU.u_wallace._3208_ ),
    .A2(\u_cpu.ALU.u_wallace._3212_ ),
    .B1(\u_cpu.ALU.u_wallace._3213_ ),
    .Y(\u_cpu.ALU.u_wallace._3214_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8775_  (.A(\u_cpu.ALU.u_wallace._3209_ ),
    .B(\u_cpu.ALU.u_wallace._3211_ ),
    .Y(\u_cpu.ALU.u_wallace._3215_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8776_  (.A1(\u_cpu.ALU.u_wallace._3203_ ),
    .A2(\u_cpu.ALU.u_wallace._3215_ ),
    .B1(\u_cpu.ALU.u_wallace._3208_ ),
    .C1(\u_cpu.ALU.u_wallace._3213_ ),
    .X(\u_cpu.ALU.u_wallace._3216_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8777_  (.A1(\u_cpu.ALU.u_wallace._3189_ ),
    .A2(\u_cpu.ALU.u_wallace._3192_ ),
    .B1(\u_cpu.ALU.u_wallace._3214_ ),
    .B2(\u_cpu.ALU.u_wallace._3216_ ),
    .Y(\u_cpu.ALU.u_wallace._3217_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8778_  (.A1(\u_cpu.ALU.u_wallace._3208_ ),
    .A2(\u_cpu.ALU.u_wallace._3212_ ),
    .B1(\u_cpu.ALU.u_wallace._3213_ ),
    .X(\u_cpu.ALU.u_wallace._3219_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8779_  (.A1(\u_cpu.ALU.u_wallace._3203_ ),
    .A2(\u_cpu.ALU.u_wallace._3215_ ),
    .B1(\u_cpu.ALU.u_wallace._3208_ ),
    .C1(\u_cpu.ALU.u_wallace._3213_ ),
    .Y(\u_cpu.ALU.u_wallace._3220_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8780_  (.A1(\u_cpu.ALU.u_wallace._3183_ ),
    .A2(\u_cpu.ALU.u_wallace._3186_ ),
    .B1(\u_cpu.ALU.u_wallace._3190_ ),
    .Y(\u_cpu.ALU.u_wallace._3221_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._8781_  (.A1(\u_cpu.ALU.u_wallace._3186_ ),
    .A2(\u_cpu.ALU.u_wallace._3191_ ),
    .B1(\u_cpu.ALU.u_wallace._3221_ ),
    .X(\u_cpu.ALU.u_wallace._3222_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8782_  (.A(\u_cpu.ALU.u_wallace._3219_ ),
    .B(\u_cpu.ALU.u_wallace._3220_ ),
    .C(\u_cpu.ALU.u_wallace._3222_ ),
    .Y(\u_cpu.ALU.u_wallace._3223_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8783_  (.A1(\u_cpu.ALU.u_wallace._2850_ ),
    .A2(\u_cpu.ALU.u_wallace._2946_ ),
    .B1(\u_cpu.ALU.u_wallace._3217_ ),
    .C1(\u_cpu.ALU.u_wallace._3223_ ),
    .X(\u_cpu.ALU.u_wallace._3224_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._8784_  (.A1(\u_cpu.ALU.u_wallace._3046_ ),
    .A2(\u_cpu.ALU.u_wallace._2942_ ),
    .B1(\u_cpu.ALU.u_wallace._2858_ ),
    .B2(\u_cpu.ALU.u_wallace._2857_ ),
    .X(\u_cpu.ALU.u_wallace._3225_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8785_  (.A(\u_cpu.ALU.u_wallace._3217_ ),
    .B(\u_cpu.ALU.u_wallace._3223_ ),
    .Y(\u_cpu.ALU.u_wallace._3226_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8786_  (.A1(\u_cpu.ALU.u_wallace._2776_ ),
    .A2(\u_cpu.ALU.u_wallace._2778_ ),
    .B1(\u_cpu.ALU.u_wallace._2799_ ),
    .C1(\u_cpu.ALU.u_wallace._2811_ ),
    .X(\u_cpu.ALU.u_wallace._3227_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8787_  (.A1_N(\u_cpu.ALU.u_wallace._3225_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3226_ ),
    .B1(\u_cpu.ALU.u_wallace._2804_ ),
    .B2(\u_cpu.ALU.u_wallace._3227_ ),
    .Y(\u_cpu.ALU.u_wallace._3228_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8788_  (.A1(\u_cpu.ALU.u_wallace._3046_ ),
    .A2(\u_cpu.ALU.u_wallace._2942_ ),
    .B1(\u_cpu.ALU.u_wallace._2858_ ),
    .B2(\u_cpu.ALU.u_wallace._2857_ ),
    .Y(\u_cpu.ALU.u_wallace._3230_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8789_  (.A1(\u_cpu.ALU.u_wallace._3217_ ),
    .A2(\u_cpu.ALU.u_wallace._3223_ ),
    .B1(\u_cpu.ALU.u_wallace._3230_ ),
    .Y(\u_cpu.ALU.u_wallace._3231_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.ALU.u_wallace._8790_  (.A1(\u_cpu.ALU.u_wallace._2802_ ),
    .A2(\u_cpu.ALU.u_wallace._2803_ ),
    .A3(\u_cpu.ALU.u_wallace._2775_ ),
    .B1(\u_cpu.ALU.u_wallace._2778_ ),
    .B2(\u_cpu.ALU.u_wallace._2776_ ),
    .X(\u_cpu.ALU.u_wallace._3232_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8791_  (.A1(\u_cpu.ALU.u_wallace._3231_ ),
    .A2(\u_cpu.ALU.u_wallace._3224_ ),
    .B1(\u_cpu.ALU.u_wallace._3232_ ),
    .Y(\u_cpu.ALU.u_wallace._3233_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8792_  (.A1(\u_cpu.ALU.u_wallace._3224_ ),
    .A2(\u_cpu.ALU.u_wallace._3228_ ),
    .B1(\u_cpu.ALU.u_wallace._3233_ ),
    .Y(\u_cpu.ALU.u_wallace._3234_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8793_  (.A1(\u_cpu.ALU.u_wallace._3051_ ),
    .A2(\u_cpu.ALU.u_wallace._3171_ ),
    .B1(\u_cpu.ALU.u_wallace._3234_ ),
    .Y(\u_cpu.ALU.u_wallace._3235_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8794_  (.A1(\u_cpu.ALU.u_wallace._3044_ ),
    .A2(\u_cpu.ALU.u_wallace._3045_ ),
    .B1(\u_cpu.ALU.u_wallace._3049_ ),
    .B2(\u_cpu.ALU.u_wallace._3050_ ),
    .Y(\u_cpu.ALU.u_wallace._3236_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8795_  (.A1(\u_cpu.ALU.u_wallace._3117_ ),
    .A2(\u_cpu.ALU.u_wallace._3166_ ),
    .B1(\u_cpu.ALU.u_wallace._3170_ ),
    .C1(\u_cpu.ALU.u_wallace._3236_ ),
    .Y(\u_cpu.ALU.u_wallace._3237_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8796_  (.A(\u_cpu.ALU.u_wallace._3165_ ),
    .B(\u_cpu.ALU.u_wallace._3124_ ),
    .C(\u_cpu.ALU.u_wallace._3167_ ),
    .X(\u_cpu.ALU.u_wallace._3238_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8797_  (.A(\u_cpu.ALU.u_wallace._3236_ ),
    .B(\u_cpu.ALU.u_wallace._3170_ ),
    .Y(\u_cpu.ALU.u_wallace._3239_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8798_  (.A(\u_cpu.ALU.u_wallace._3165_ ),
    .B(\u_cpu.ALU.u_wallace._3124_ ),
    .C(\u_cpu.ALU.u_wallace._3167_ ),
    .Y(\u_cpu.ALU.u_wallace._3241_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8799_  (.A1(\u_cpu.ALU.u_wallace._3241_ ),
    .A2(\u_cpu.ALU.u_wallace._3170_ ),
    .B1(\u_cpu.ALU.u_wallace._3236_ ),
    .X(\u_cpu.ALU.u_wallace._3242_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8800_  (.A1(\u_cpu.ALU.u_wallace._3238_ ),
    .A2(\u_cpu.ALU.u_wallace._3239_ ),
    .B1(\u_cpu.ALU.u_wallace._3242_ ),
    .Y(\u_cpu.ALU.u_wallace._3243_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8801_  (.A1(\u_cpu.ALU.u_wallace._3235_ ),
    .A2(\u_cpu.ALU.u_wallace._3237_ ),
    .B1(\u_cpu.ALU.u_wallace._3234_ ),
    .B2(\u_cpu.ALU.u_wallace._3243_ ),
    .Y(\u_cpu.ALU.u_wallace._3244_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8802_  (.A(\u_cpu.ALU.u_wallace._3236_ ),
    .B(\u_cpu.ALU.u_wallace._3241_ ),
    .C(\u_cpu.ALU.u_wallace._3170_ ),
    .X(\u_cpu.ALU.u_wallace._3245_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8803_  (.A1(\u_cpu.ALU.u_wallace._3051_ ),
    .A2(\u_cpu.ALU.u_wallace._3171_ ),
    .B1(\u_cpu.ALU.u_wallace._3234_ ),
    .X(\u_cpu.ALU.u_wallace._3246_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._8804_  (.A1(\u_cpu.ALU.u_wallace._2776_ ),
    .A2(\u_cpu.ALU.u_wallace._2778_ ),
    .B1(\u_cpu.ALU.u_wallace._3231_ ),
    .B2(\u_cpu.ALU.u_wallace._3224_ ),
    .C1(\u_cpu.ALU.u_wallace._2813_ ),
    .X(\u_cpu.ALU.u_wallace._3247_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8805_  (.A1(\u_cpu.ALU.u_wallace._3226_ ),
    .A2(\u_cpu.ALU.u_wallace._3225_ ),
    .B1(\u_cpu.ALU.u_wallace._3232_ ),
    .Y(\u_cpu.ALU.u_wallace._3248_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._8806_  (.A1(\u_cpu.ALU.u_wallace._3225_ ),
    .A2(\u_cpu.ALU.u_wallace._3226_ ),
    .B1(\u_cpu.ALU.u_wallace._3248_ ),
    .X(\u_cpu.ALU.u_wallace._3249_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8807_  (.A1_N(\u_cpu.ALU.u_wallace._3237_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3242_ ),
    .B1(\u_cpu.ALU.u_wallace._3247_ ),
    .B2(\u_cpu.ALU.u_wallace._3249_ ),
    .Y(\u_cpu.ALU.u_wallace._3250_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8808_  (.A1(\u_cpu.ALU.u_wallace._3245_ ),
    .A2(\u_cpu.ALU.u_wallace._3246_ ),
    .B1(\u_cpu.ALU.u_wallace._3250_ ),
    .C1(\u_cpu.ALU.u_wallace._3043_ ),
    .Y(\u_cpu.ALU.u_wallace._3252_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8809_  (.A(\u_cpu.ALU.u_wallace._0917_ ),
    .X(\u_cpu.ALU.u_wallace._3253_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8810_  (.A(\u_cpu.ALU.SrcB[27] ),
    .X(\u_cpu.ALU.u_wallace._3254_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8811_  (.A1(\u_cpu.ALU.u_wallace._0261_ ),
    .A2(\u_cpu.ALU.SrcB[26] ),
    .B1(\u_cpu.ALU.u_wallace._3254_ ),
    .B2(\u_cpu.ALU.u_wallace._0994_ ),
    .Y(\u_cpu.ALU.u_wallace._3255_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8812_  (.A(\u_cpu.ALU.u_wallace._0446_ ),
    .B(\u_cpu.ALU.u_wallace._0261_ ),
    .C(\u_cpu.ALU.SrcB[26] ),
    .D(\u_cpu.ALU.SrcB[27] ),
    .X(\u_cpu.ALU.u_wallace._3256_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8813_  (.A1(\u_cpu.ALU.u_wallace._0414_ ),
    .A2(\u_cpu.ALU.u_wallace._2481_ ),
    .B1(\u_cpu.ALU.u_wallace._3255_ ),
    .B2(\u_cpu.ALU.u_wallace._3256_ ),
    .Y(\u_cpu.ALU.u_wallace._3257_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8814_  (.A(\u_cpu.ALU.SrcB[26] ),
    .X(\u_cpu.ALU.u_wallace._3258_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8815_  (.A1(\u_cpu.ALU.u_wallace._4463_ ),
    .A2(\u_cpu.ALU.u_wallace._3258_ ),
    .B1(\u_cpu.ALU.u_wallace._3254_ ),
    .B2(\u_cpu.ALU.u_wallace._0994_ ),
    .X(\u_cpu.ALU.u_wallace._3259_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8816_  (.A(\u_cpu.ALU.u_wallace._0994_ ),
    .B(\u_cpu.ALU.u_wallace._4463_ ),
    .C(\u_cpu.ALU.u_wallace._3258_ ),
    .D(\u_cpu.ALU.u_wallace._3254_ ),
    .Y(\u_cpu.ALU.u_wallace._3260_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8817_  (.A(\u_cpu.ALU.u_wallace._3259_ ),
    .B(\u_cpu.ALU.u_wallace._3260_ ),
    .C(\u_cpu.ALU.u_wallace._0370_ ),
    .D(\u_cpu.ALU.u_wallace._2480_ ),
    .Y(\u_cpu.ALU.u_wallace._3261_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._8818_  (.A(\u_cpu.ALU.u_wallace._3258_ ),
    .Y(\u_cpu.ALU.u_wallace._3263_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8819_  (.A(\u_cpu.ALU.u_wallace._0118_ ),
    .B(\u_cpu.ALU.u_wallace._0173_ ),
    .C(\u_cpu.ALU.u_wallace._2480_ ),
    .Y(\u_cpu.ALU.u_wallace._3264_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8820_  (.A1_N(\u_cpu.ALU.u_wallace._3257_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3261_ ),
    .B1(\u_cpu.ALU.u_wallace._3263_ ),
    .B2(\u_cpu.ALU.u_wallace._3264_ ),
    .Y(\u_cpu.ALU.u_wallace._3265_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8821_  (.A(\u_cpu.ALU.u_wallace._3257_ ),
    .B(\u_cpu.ALU.u_wallace._3261_ ),
    .C(\u_cpu.ALU.u_wallace._2982_ ),
    .Y(\u_cpu.ALU.u_wallace._3266_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8822_  (.A1(\u_cpu.ALU.u_wallace._2986_ ),
    .A2(\u_cpu.ALU.u_wallace._2397_ ),
    .B1(\u_cpu.ALU.u_wallace._3265_ ),
    .B2(\u_cpu.ALU.u_wallace._3266_ ),
    .Y(\u_cpu.ALU.u_wallace._3267_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8823_  (.A(\u_cpu.ALU.u_wallace._2986_ ),
    .B(\u_cpu.ALU.u_wallace._2397_ ),
    .Y(\u_cpu.ALU.u_wallace._3268_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8824_  (.A1(\u_cpu.ALU.u_wallace._3257_ ),
    .A2(\u_cpu.ALU.u_wallace._3261_ ),
    .B1(\u_cpu.ALU.u_wallace._2982_ ),
    .Y(\u_cpu.ALU.u_wallace._3269_ ));
 sky130_fd_sc_hd__nor3b_2 \u_cpu.ALU.u_wallace._8825_  (.A(\u_cpu.ALU.u_wallace._3268_ ),
    .B(\u_cpu.ALU.u_wallace._3269_ ),
    .C_N(\u_cpu.ALU.u_wallace._3266_ ),
    .Y(\u_cpu.ALU.u_wallace._3270_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8826_  (.A1(\u_cpu.ALU.u_wallace._3267_ ),
    .A2(\u_cpu.ALU.u_wallace._3270_ ),
    .B1(\u_cpu.ALU.u_wallace._2981_ ),
    .Y(\u_cpu.ALU.u_wallace._3271_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8827_  (.A1(\u_cpu.ALU.u_wallace._2986_ ),
    .A2(\u_cpu.ALU.u_wallace._2397_ ),
    .B1(\u_cpu.ALU.u_wallace._3265_ ),
    .B2(\u_cpu.ALU.u_wallace._3266_ ),
    .X(\u_cpu.ALU.u_wallace._3272_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8828_  (.A(\u_cpu.ALU.u_wallace._3265_ ),
    .B(\u_cpu.ALU.u_wallace._3266_ ),
    .C(\u_cpu.ALU.u_wallace._2986_ ),
    .D(\u_cpu.ALU.u_wallace._2402_ ),
    .Y(\u_cpu.ALU.u_wallace._3274_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._8829_  (.A_N(\u_cpu.ALU.u_wallace._2981_ ),
    .B(\u_cpu.ALU.u_wallace._3272_ ),
    .C(\u_cpu.ALU.u_wallace._3274_ ),
    .Y(\u_cpu.ALU.u_wallace._3275_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8830_  (.A1(\u_cpu.ALU.u_wallace._3253_ ),
    .A2(\u_cpu.ALU.u_wallace._2134_ ),
    .B1(\u_cpu.ALU.u_wallace._3271_ ),
    .B2(\u_cpu.ALU.u_wallace._3275_ ),
    .X(\u_cpu.ALU.u_wallace._3276_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8831_  (.A(\u_cpu.ALU.u_wallace._3271_ ),
    .B(\u_cpu.ALU.u_wallace._3275_ ),
    .C(\u_cpu.ALU.u_wallace._3253_ ),
    .D(\u_cpu.ALU.u_wallace._2134_ ),
    .Y(\u_cpu.ALU.u_wallace._3277_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._8832_  (.A1(\u_cpu.ALU.u_wallace._2787_ ),
    .A2(\u_cpu.ALU.u_wallace._2789_ ),
    .A3(\u_cpu.ALU.u_wallace._2791_ ),
    .B1(\u_cpu.ALU.u_wallace._2794_ ),
    .Y(\u_cpu.ALU.u_wallace._3278_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8833_  (.A(\u_cpu.ALU.u_wallace._2794_ ),
    .B(\u_cpu.ALU.u_wallace._2791_ ),
    .C(\u_cpu.ALU.u_wallace._2789_ ),
    .D(\u_cpu.ALU.u_wallace._2787_ ),
    .X(\u_cpu.ALU.u_wallace._3279_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8834_  (.A1(\u_cpu.ALU.u_wallace._3278_ ),
    .A2(\u_cpu.ALU.u_wallace._3279_ ),
    .B1(\u_cpu.ALU.u_wallace._2798_ ),
    .Y(\u_cpu.ALU.u_wallace._3280_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8835_  (.A1(\u_cpu.ALU.u_wallace._3278_ ),
    .A2(\u_cpu.ALU.u_wallace._3279_ ),
    .B1(\u_cpu.ALU.u_wallace._2973_ ),
    .C1(\u_cpu.ALU.u_wallace._2798_ ),
    .X(\u_cpu.ALU.u_wallace._3281_ ));
 sky130_fd_sc_hd__a41oi_2 \u_cpu.ALU.u_wallace._8836_  (.A1(\u_cpu.ALU.u_wallace._2554_ ),
    .A2(\u_cpu.ALU.u_wallace._3280_ ),
    .A3(\u_cpu.ALU.u_wallace._2514_ ),
    .A4(\u_cpu.ALU.u_wallace._2511_ ),
    .B1(\u_cpu.ALU.u_wallace._3281_ ),
    .Y(\u_cpu.ALU.u_wallace._3282_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8837_  (.A1(\u_cpu.ALU.u_wallace._3276_ ),
    .A2(\u_cpu.ALU.u_wallace._3277_ ),
    .B1(\u_cpu.ALU.u_wallace._3282_ ),
    .X(\u_cpu.ALU.u_wallace._3283_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8838_  (.A(\u_cpu.ALU.u_wallace._3276_ ),
    .B(\u_cpu.ALU.u_wallace._3277_ ),
    .C(\u_cpu.ALU.u_wallace._3282_ ),
    .Y(\u_cpu.ALU.u_wallace._3285_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8839_  (.A(\u_cpu.ALU.u_wallace._3283_ ),
    .B(\u_cpu.ALU.u_wallace._3285_ ),
    .Y(\u_cpu.ALU.u_wallace._3286_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8840_  (.A(\u_cpu.ALU.u_wallace._2958_ ),
    .B(\u_cpu.ALU.u_wallace._2808_ ),
    .C(\u_cpu.ALU.u_wallace._3286_ ),
    .Y(\u_cpu.ALU.u_wallace._3287_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._8841_  (.A(\u_cpu.ALU.u_wallace._3276_ ),
    .B(\u_cpu.ALU.u_wallace._3282_ ),
    .X(\u_cpu.ALU.u_wallace._3288_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8842_  (.A1(\u_cpu.ALU.u_wallace._3276_ ),
    .A2(\u_cpu.ALU.u_wallace._3277_ ),
    .B1(\u_cpu.ALU.u_wallace._3282_ ),
    .Y(\u_cpu.ALU.u_wallace._3289_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8843_  (.A1(\u_cpu.ALU.u_wallace._3288_ ),
    .A2(\u_cpu.ALU.u_wallace._3277_ ),
    .B1(\u_cpu.ALU.u_wallace._3289_ ),
    .Y(\u_cpu.ALU.u_wallace._3290_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8844_  (.A1(\u_cpu.ALU.u_wallace._2810_ ),
    .A2(\u_cpu.ALU.u_wallace._2965_ ),
    .B1(\u_cpu.ALU.u_wallace._3290_ ),
    .Y(\u_cpu.ALU.u_wallace._3291_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8845_  (.A1(\u_cpu.ALU.u_wallace._2991_ ),
    .A2(\u_cpu.ALU.u_wallace._2993_ ),
    .B1(\u_cpu.ALU.u_wallace._2975_ ),
    .Y(\u_cpu.ALU.u_wallace._3292_ ));
 sky130_fd_sc_hd__a21bo_2 \u_cpu.ALU.u_wallace._8846_  (.A1(\u_cpu.ALU.u_wallace._3287_ ),
    .A2(\u_cpu.ALU.u_wallace._3291_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3292_ ),
    .X(\u_cpu.ALU.u_wallace._3293_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._8847_  (.A_N(\u_cpu.ALU.u_wallace._3292_ ),
    .B(\u_cpu.ALU.u_wallace._3287_ ),
    .C(\u_cpu.ALU.u_wallace._3291_ ),
    .Y(\u_cpu.ALU.u_wallace._3294_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._8848_  (.A1(\u_cpu.ALU.u_wallace._3043_ ),
    .A2(\u_cpu.ALU.u_wallace._3244_ ),
    .B1(\u_cpu.ALU.u_wallace._3252_ ),
    .C1(\u_cpu.ALU.u_wallace._3293_ ),
    .D1(\u_cpu.ALU.u_wallace._3294_ ),
    .Y(\u_cpu.ALU.u_wallace._3296_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.ALU.u_wallace._8849_  (.A1(\u_cpu.ALU.u_wallace._2991_ ),
    .A2(\u_cpu.ALU.u_wallace._2993_ ),
    .B1(\u_cpu.ALU.u_wallace._3291_ ),
    .B2(\u_cpu.ALU.u_wallace._3287_ ),
    .C1(\u_cpu.ALU.u_wallace._2975_ ),
    .Y(\u_cpu.ALU.u_wallace._3297_ ));
 sky130_fd_sc_hd__and3b_2 \u_cpu.ALU.u_wallace._8850_  (.A_N(\u_cpu.ALU.u_wallace._3292_ ),
    .B(\u_cpu.ALU.u_wallace._3287_ ),
    .C(\u_cpu.ALU.u_wallace._3291_ ),
    .X(\u_cpu.ALU.u_wallace._3298_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._8851_  (.A1(\u_cpu.ALU.u_wallace._3224_ ),
    .A2(\u_cpu.ALU.u_wallace._3228_ ),
    .B1(\u_cpu.ALU.u_wallace._3233_ ),
    .C1(\u_cpu.ALU.u_wallace._3237_ ),
    .D1(\u_cpu.ALU.u_wallace._3242_ ),
    .Y(\u_cpu.ALU.u_wallace._3299_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8852_  (.A1(\u_cpu.ALU.u_wallace._3299_ ),
    .A2(\u_cpu.ALU.u_wallace._3250_ ),
    .B1(\u_cpu.ALU.u_wallace._3043_ ),
    .Y(\u_cpu.ALU.u_wallace._3300_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8853_  (.A1(\u_cpu.ALU.u_wallace._3245_ ),
    .A2(\u_cpu.ALU.u_wallace._3246_ ),
    .B1(\u_cpu.ALU.u_wallace._3250_ ),
    .C1(\u_cpu.ALU.u_wallace._3043_ ),
    .X(\u_cpu.ALU.u_wallace._3301_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8854_  (.A1(\u_cpu.ALU.u_wallace._3297_ ),
    .A2(\u_cpu.ALU.u_wallace._3298_ ),
    .B1(\u_cpu.ALU.u_wallace._3300_ ),
    .B2(\u_cpu.ALU.u_wallace._3301_ ),
    .Y(\u_cpu.ALU.u_wallace._3302_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8855_  (.A1(\u_cpu.ALU.u_wallace._2971_ ),
    .A2(\u_cpu.ALU.u_wallace._3005_ ),
    .B1(\u_cpu.ALU.u_wallace._3012_ ),
    .X(\u_cpu.ALU.u_wallace._3303_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8856_  (.A1(\u_cpu.ALU.u_wallace._3296_ ),
    .A2(\u_cpu.ALU.u_wallace._3302_ ),
    .B1(\u_cpu.ALU.u_wallace._3303_ ),
    .Y(\u_cpu.ALU.u_wallace._3304_ ));
 sky130_fd_sc_hd__a311oi_2 \u_cpu.ALU.u_wallace._8857_  (.A1(\u_cpu.ALU.u_wallace._2964_ ),
    .A2(\u_cpu.ALU.u_wallace._2968_ ),
    .A3(\u_cpu.ALU.u_wallace._2970_ ),
    .B1(\u_cpu.ALU.u_wallace._3004_ ),
    .C1(\u_cpu.ALU.u_wallace._3003_ ),
    .Y(\u_cpu.ALU.u_wallace._3305_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8858_  (.A1(\u_cpu.ALU.u_wallace._3012_ ),
    .A2(\u_cpu.ALU.u_wallace._3305_ ),
    .B1(\u_cpu.ALU.u_wallace._3296_ ),
    .C1(\u_cpu.ALU.u_wallace._3302_ ),
    .X(\u_cpu.ALU.u_wallace._3307_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._8859_  (.A1(\u_cpu.ALU.u_wallace._3002_ ),
    .A2(\u_cpu.ALU.u_wallace._2997_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3000_ ),
    .Y(\u_cpu.ALU.u_wallace._3308_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8860_  (.A1(\u_cpu.ALU.u_wallace._3304_ ),
    .A2(\u_cpu.ALU.u_wallace._3307_ ),
    .B1(\u_cpu.ALU.u_wallace._3308_ ),
    .Y(\u_cpu.ALU.u_wallace._3309_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._8861_  (.A(\u_cpu.ALU.u_wallace._3308_ ),
    .Y(\u_cpu.ALU.u_wallace._3310_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8862_  (.A1(\u_cpu.ALU.u_wallace._3296_ ),
    .A2(\u_cpu.ALU.u_wallace._3302_ ),
    .B1(\u_cpu.ALU.u_wallace._3303_ ),
    .X(\u_cpu.ALU.u_wallace._3311_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8863_  (.A1(\u_cpu.ALU.u_wallace._3012_ ),
    .A2(\u_cpu.ALU.u_wallace._3305_ ),
    .B1(\u_cpu.ALU.u_wallace._3296_ ),
    .C1(\u_cpu.ALU.u_wallace._3302_ ),
    .Y(\u_cpu.ALU.u_wallace._3312_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8864_  (.A(\u_cpu.ALU.u_wallace._3310_ ),
    .B(\u_cpu.ALU.u_wallace._3311_ ),
    .C(\u_cpu.ALU.u_wallace._3312_ ),
    .Y(\u_cpu.ALU.u_wallace._3313_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8865_  (.A1(\u_cpu.ALU.u_wallace._2498_ ),
    .A2(\u_cpu.ALU.u_wallace._2727_ ),
    .B1(\u_cpu.ALU.u_wallace._3009_ ),
    .Y(\u_cpu.ALU.u_wallace._3314_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8866_  (.A(\u_cpu.ALU.u_wallace._3015_ ),
    .B(\u_cpu.ALU.u_wallace._3314_ ),
    .Y(\u_cpu.ALU.u_wallace._3315_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8867_  (.A1(\u_cpu.ALU.u_wallace._3309_ ),
    .A2(\u_cpu.ALU.u_wallace._3313_ ),
    .B1(\u_cpu.ALU.u_wallace._3315_ ),
    .Y(\u_cpu.ALU.u_wallace._3316_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8868_  (.A(\u_cpu.ALU.u_wallace._3308_ ),
    .B(\u_cpu.ALU.u_wallace._3304_ ),
    .Y(\u_cpu.ALU.u_wallace._3318_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8869_  (.A1(\u_cpu.ALU.u_wallace._3311_ ),
    .A2(\u_cpu.ALU.u_wallace._3312_ ),
    .B1(\u_cpu.ALU.u_wallace._3310_ ),
    .Y(\u_cpu.ALU.u_wallace._3319_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.ALU.u_wallace._8870_  (.A1(\u_cpu.ALU.u_wallace._3015_ ),
    .A2(\u_cpu.ALU.u_wallace._3314_ ),
    .B1(\u_cpu.ALU.u_wallace._3318_ ),
    .B2(\u_cpu.ALU.u_wallace._3312_ ),
    .C1(\u_cpu.ALU.u_wallace._3319_ ),
    .Y(\u_cpu.ALU.u_wallace._3320_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.ALU.u_wallace._8871_  (.A_N(\u_cpu.ALU.u_wallace._2985_ ),
    .B(\u_cpu.ALU.u_wallace._2417_ ),
    .C(\u_cpu.ALU.u_wallace._2986_ ),
    .D(\u_cpu.ALU.u_wallace._2989_ ),
    .X(\u_cpu.ALU.u_wallace._3321_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8872_  (.A(\u_cpu.ALU.u_wallace._2985_ ),
    .B(\u_cpu.ALU.u_wallace._3321_ ),
    .Y(\u_cpu.ALU.u_wallace._3322_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8873_  (.A1(\u_cpu.ALU.u_wallace._3316_ ),
    .A2(\u_cpu.ALU.u_wallace._3320_ ),
    .B1(\u_cpu.ALU.u_wallace._3322_ ),
    .Y(\u_cpu.ALU.u_wallace._3323_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8874_  (.A1(\u_cpu.ALU.u_wallace._3309_ ),
    .A2(\u_cpu.ALU.u_wallace._3313_ ),
    .B1(\u_cpu.ALU.u_wallace._3315_ ),
    .X(\u_cpu.ALU.u_wallace._3324_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8875_  (.A(\u_cpu.ALU.u_wallace._3315_ ),
    .B(\u_cpu.ALU.u_wallace._3309_ ),
    .C(\u_cpu.ALU.u_wallace._3313_ ),
    .Y(\u_cpu.ALU.u_wallace._3325_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8876_  (.A1(\u_cpu.ALU.u_wallace._2985_ ),
    .A2(\u_cpu.ALU.u_wallace._3321_ ),
    .B1(\u_cpu.ALU.u_wallace._3324_ ),
    .C1(\u_cpu.ALU.u_wallace._3325_ ),
    .Y(\u_cpu.ALU.u_wallace._3326_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._8877_  (.A1(\u_cpu.ALU.u_wallace._2756_ ),
    .A2(\u_cpu.ALU.u_wallace._3017_ ),
    .A3(\u_cpu.ALU.u_wallace._3018_ ),
    .B1(\u_cpu.ALU.u_wallace._3024_ ),
    .B2(\u_cpu.ALU.u_wallace._2486_ ),
    .X(\u_cpu.ALU.u_wallace._3327_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8878_  (.A1(\u_cpu.ALU.u_wallace._3323_ ),
    .A2(\u_cpu.ALU.u_wallace._3326_ ),
    .B1(\u_cpu.ALU.u_wallace._3327_ ),
    .Y(\u_cpu.ALU.u_wallace._3329_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8879_  (.A1(\u_cpu.ALU.u_wallace._2985_ ),
    .A2(\u_cpu.ALU.u_wallace._3321_ ),
    .B1(\u_cpu.ALU.u_wallace._3324_ ),
    .Y(\u_cpu.ALU.u_wallace._3330_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8880_  (.A1(\u_cpu.ALU.u_wallace._3320_ ),
    .A2(\u_cpu.ALU.u_wallace._3330_ ),
    .B1(\u_cpu.ALU.u_wallace._3323_ ),
    .C1(\u_cpu.ALU.u_wallace._3327_ ),
    .X(\u_cpu.ALU.u_wallace._3331_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8881_  (.A(\u_cpu.ALU.u_wallace._3329_ ),
    .B(\u_cpu.ALU.u_wallace._3331_ ),
    .Y(\u_cpu.ALU.u_wallace._3332_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._8882_  (.A1(\u_cpu.ALU.u_wallace._2401_ ),
    .A2(\u_cpu.ALU.u_wallace._3029_ ),
    .B1(\u_cpu.ALU.u_wallace._3025_ ),
    .B2(\u_cpu.ALU.u_wallace._3027_ ),
    .C1(\u_cpu.ALU.u_wallace._2745_ ),
    .X(\u_cpu.ALU.u_wallace._3333_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8883_  (.A1(\u_cpu.ALU.u_wallace._3333_ ),
    .A2(\u_cpu.ALU.u_wallace._3041_ ),
    .B1(\u_cpu.ALU.u_wallace._3036_ ),
    .Y(\u_cpu.ALU.u_wallace._3334_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._8884_  (.A(\u_cpu.ALU.u_wallace._3332_ ),
    .B(\u_cpu.ALU.u_wallace._3334_ ),
    .X(\u_cpu.ALU.Product_Wallace[27] ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._8885_  (.A1(\u_cpu.ALU.u_wallace._3322_ ),
    .A2(\u_cpu.ALU.u_wallace._3316_ ),
    .B1(\u_cpu.ALU.u_wallace._3325_ ),
    .X(\u_cpu.ALU.u_wallace._3335_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.ALU.u_wallace._8886_  (.A_N(\u_cpu.ALU.u_wallace._2978_ ),
    .B(\u_cpu.ALU.u_wallace._2979_ ),
    .C(\u_cpu.ALU.u_wallace._3272_ ),
    .D(\u_cpu.ALU.u_wallace._2980_ ),
    .X(\u_cpu.ALU.u_wallace._3336_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._8887_  (.A1(\u_cpu.ALU.u_wallace._3271_ ),
    .A2(\u_cpu.ALU.u_wallace._2417_ ),
    .A3(\u_cpu.ALU.u_wallace._3253_ ),
    .B1(\u_cpu.ALU.u_wallace._3274_ ),
    .B2(\u_cpu.ALU.u_wallace._3336_ ),
    .X(\u_cpu.ALU.u_wallace._3337_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._8888_  (.A(\u_cpu.ALU.u_wallace._3337_ ),
    .Y(\u_cpu.ALU.u_wallace._3339_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8889_  (.A(\u_cpu.ALU.u_wallace._3293_ ),
    .B(\u_cpu.ALU.u_wallace._3294_ ),
    .Y(\u_cpu.ALU.u_wallace._3340_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8890_  (.A(\u_cpu.ALU.u_wallace._3340_ ),
    .B(\u_cpu.ALU.u_wallace._3300_ ),
    .Y(\u_cpu.ALU.u_wallace._3341_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8891_  (.A(\u_cpu.ALU.u_wallace._3201_ ),
    .B(\u_cpu.ALU.u_wallace._3206_ ),
    .Y(\u_cpu.ALU.u_wallace._3342_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8892_  (.A(\u_cpu.ALU.u_wallace._0319_ ),
    .B(\u_cpu.ALU.u_wallace._0320_ ),
    .C(\u_cpu.ALU.u_wallace._0121_ ),
    .D(\u_cpu.ALU.u_wallace._0279_ ),
    .Y(\u_cpu.ALU.u_wallace._3343_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8893_  (.A1(\u_cpu.ALU.u_wallace._0179_ ),
    .A2(\u_cpu.ALU.u_wallace._0546_ ),
    .B1(\u_cpu.ALU.u_wallace._0547_ ),
    .B2(\u_cpu.ALU.u_wallace._0188_ ),
    .X(\u_cpu.ALU.u_wallace._3344_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8894_  (.A1_N(\u_cpu.ALU.u_wallace._3343_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3344_ ),
    .B1(\u_cpu.ALU.u_wallace._4913_ ),
    .B2(\u_cpu.ALU.u_wallace._0554_ ),
    .Y(\u_cpu.ALU.u_wallace._3345_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8895_  (.A(\u_cpu.ALU.u_wallace._3344_ ),
    .B(\u_cpu.ALU.u_wallace._0551_ ),
    .C(\u_cpu.ALU.u_wallace._0475_ ),
    .D(\u_cpu.ALU.u_wallace._3343_ ),
    .Y(\u_cpu.ALU.u_wallace._3346_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8896_  (.A1(\u_cpu.ALU.u_wallace._3138_ ),
    .A2(\u_cpu.ALU.u_wallace._3137_ ),
    .B1(\u_cpu.ALU.u_wallace._3133_ ),
    .Y(\u_cpu.ALU.u_wallace._3347_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8897_  (.A1(\u_cpu.ALU.u_wallace._3345_ ),
    .A2(\u_cpu.ALU.u_wallace._3346_ ),
    .B1(\u_cpu.ALU.u_wallace._3347_ ),
    .Y(\u_cpu.ALU.u_wallace._3348_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8898_  (.A(\u_cpu.ALU.u_wallace._3347_ ),
    .B(\u_cpu.ALU.u_wallace._3345_ ),
    .C(\u_cpu.ALU.u_wallace._3346_ ),
    .X(\u_cpu.ALU.u_wallace._3350_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8899_  (.A1(\u_cpu.ALU.u_wallace._3197_ ),
    .A2(\u_cpu.ALU.u_wallace._0551_ ),
    .A3(\u_cpu.ALU.u_wallace._1129_ ),
    .B1(\u_cpu.ALU.u_wallace._3194_ ),
    .X(\u_cpu.ALU.u_wallace._3351_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._8900_  (.A1(\u_cpu.ALU.u_wallace._3348_ ),
    .A2(\u_cpu.ALU.u_wallace._3350_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3351_ ),
    .Y(\u_cpu.ALU.u_wallace._3352_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8901_  (.A(\u_cpu.ALU.u_wallace._3347_ ),
    .B(\u_cpu.ALU.u_wallace._3345_ ),
    .Y(\u_cpu.ALU.u_wallace._3353_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8902_  (.A(\u_cpu.ALU.u_wallace._3344_ ),
    .B(\u_cpu.ALU.u_wallace._3204_ ),
    .C(\u_cpu.ALU.u_wallace._2658_ ),
    .D(\u_cpu.ALU.u_wallace._3343_ ),
    .X(\u_cpu.ALU.u_wallace._3354_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8903_  (.A1(\u_cpu.ALU.u_wallace._3345_ ),
    .A2(\u_cpu.ALU.u_wallace._3346_ ),
    .B1(\u_cpu.ALU.u_wallace._3347_ ),
    .X(\u_cpu.ALU.u_wallace._3355_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8904_  (.A1(\u_cpu.ALU.u_wallace._3353_ ),
    .A2(\u_cpu.ALU.u_wallace._3354_ ),
    .B1(\u_cpu.ALU.u_wallace._3351_ ),
    .C1(\u_cpu.ALU.u_wallace._3355_ ),
    .Y(\u_cpu.ALU.u_wallace._3356_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8905_  (.A1(\u_cpu.ALU.u_wallace._3203_ ),
    .A2(\u_cpu.ALU.u_wallace._3342_ ),
    .B1(\u_cpu.ALU.u_wallace._3352_ ),
    .C1(\u_cpu.ALU.u_wallace._3356_ ),
    .X(\u_cpu.ALU.u_wallace._3357_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8906_  (.A1(\u_cpu.ALU.u_wallace._3201_ ),
    .A2(\u_cpu.ALU.u_wallace._3206_ ),
    .B1(\u_cpu.ALU.u_wallace._3210_ ),
    .Y(\u_cpu.ALU.u_wallace._3358_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8907_  (.A1(\u_cpu.ALU.u_wallace._3352_ ),
    .A2(\u_cpu.ALU.u_wallace._3356_ ),
    .B1(\u_cpu.ALU.u_wallace._3358_ ),
    .Y(\u_cpu.ALU.u_wallace._3359_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8908_  (.A1(\u_cpu.ALU.u_wallace._2343_ ),
    .A2(\u_cpu.ALU.u_wallace._1610_ ),
    .B1(\u_cpu.ALU.u_wallace._1824_ ),
    .B2(\u_cpu.ALU.u_wallace._0198_ ),
    .Y(\u_cpu.ALU.u_wallace._3361_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8909_  (.A(\u_cpu.ALU.u_wallace._4698_ ),
    .B(\u_cpu.ALU.u_wallace._0198_ ),
    .C(\u_cpu.ALU.u_wallace._1610_ ),
    .D(\u_cpu.ALU.u_wallace._1824_ ),
    .X(\u_cpu.ALU.u_wallace._3362_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU.u_wallace._8910_  (.A(\u_cpu.ALU.u_wallace._3361_ ),
    .B(\u_cpu.ALU.u_wallace._3362_ ),
    .X(\u_cpu.ALU.u_wallace._3363_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8911_  (.A1(\u_cpu.ALU.u_wallace._4554_ ),
    .A2(\u_cpu.ALU.u_wallace._1387_ ),
    .B1(\u_cpu.ALU.u_wallace._1175_ ),
    .B2(\u_cpu.ALU.u_wallace._4567_ ),
    .Y(\u_cpu.ALU.u_wallace._3364_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8912_  (.A(\u_cpu.ALU.u_wallace._4783_ ),
    .B(\u_cpu.ALU.u_wallace._4643_ ),
    .C(\u_cpu.ALU.u_wallace._0958_ ),
    .D(\u_cpu.ALU.u_wallace._1208_ ),
    .Y(\u_cpu.ALU.u_wallace._3365_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._8913_  (.A_N(\u_cpu.ALU.u_wallace._3364_ ),
    .B(\u_cpu.ALU.u_wallace._3365_ ),
    .C(\u_cpu.ALU.u_wallace._4661_ ),
    .D(\u_cpu.ALU.u_wallace._1615_ ),
    .Y(\u_cpu.ALU.u_wallace._3366_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8914_  (.A(\u_cpu.ALU.u_wallace._4567_ ),
    .B(\u_cpu.ALU.u_wallace._4554_ ),
    .C(\u_cpu.ALU.u_wallace._2050_ ),
    .D(\u_cpu.ALU.u_wallace._1175_ ),
    .X(\u_cpu.ALU.u_wallace._3367_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8915_  (.A1(\u_cpu.ALU.u_wallace._4677_ ),
    .A2(\u_cpu.ALU.u_wallace._2053_ ),
    .B1(\u_cpu.ALU.u_wallace._3364_ ),
    .B2(\u_cpu.ALU.u_wallace._3367_ ),
    .Y(\u_cpu.ALU.u_wallace._3368_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.ALU.u_wallace._8916_  (.A1(\u_cpu.ALU.u_wallace._0203_ ),
    .A2(\u_cpu.ALU.u_wallace._2053_ ),
    .A3(\u_cpu.ALU.u_wallace._3180_ ),
    .B1(\u_cpu.ALU.u_wallace._3178_ ),
    .Y(\u_cpu.ALU.u_wallace._3369_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8917_  (.A1(\u_cpu.ALU.u_wallace._3366_ ),
    .A2(\u_cpu.ALU.u_wallace._3368_ ),
    .B1(\u_cpu.ALU.u_wallace._3369_ ),
    .X(\u_cpu.ALU.u_wallace._3370_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8918_  (.A(\u_cpu.ALU.u_wallace._3369_ ),
    .B(\u_cpu.ALU.u_wallace._3366_ ),
    .C(\u_cpu.ALU.u_wallace._3368_ ),
    .Y(\u_cpu.ALU.u_wallace._3372_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8919_  (.A(\u_cpu.ALU.u_wallace._3370_ ),
    .B(\u_cpu.ALU.u_wallace._3372_ ),
    .Y(\u_cpu.ALU.u_wallace._3373_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8920_  (.A(\u_cpu.ALU.u_wallace._3363_ ),
    .B(\u_cpu.ALU.u_wallace._3373_ ),
    .Y(\u_cpu.ALU.u_wallace._3374_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._8921_  (.A1(\u_cpu.ALU.u_wallace._3361_ ),
    .A2(\u_cpu.ALU.u_wallace._3362_ ),
    .B1(\u_cpu.ALU.u_wallace._3373_ ),
    .X(\u_cpu.ALU.u_wallace._3375_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8922_  (.A(\u_cpu.ALU.u_wallace._3374_ ),
    .B(\u_cpu.ALU.u_wallace._3375_ ),
    .Y(\u_cpu.ALU.u_wallace._3376_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8923_  (.A1(\u_cpu.ALU.u_wallace._3357_ ),
    .A2(\u_cpu.ALU.u_wallace._3359_ ),
    .B1(\u_cpu.ALU.u_wallace._3376_ ),
    .Y(\u_cpu.ALU.u_wallace._3377_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8924_  (.A1(\u_cpu.ALU.u_wallace._3203_ ),
    .A2(\u_cpu.ALU.u_wallace._3342_ ),
    .B1(\u_cpu.ALU.u_wallace._3352_ ),
    .C1(\u_cpu.ALU.u_wallace._3356_ ),
    .Y(\u_cpu.ALU.u_wallace._3378_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8925_  (.A1(\u_cpu.ALU.u_wallace._3352_ ),
    .A2(\u_cpu.ALU.u_wallace._3356_ ),
    .B1(\u_cpu.ALU.u_wallace._3358_ ),
    .X(\u_cpu.ALU.u_wallace._3379_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8926_  (.A1(\u_cpu.ALU.u_wallace._3374_ ),
    .A2(\u_cpu.ALU.u_wallace._3375_ ),
    .B1(\u_cpu.ALU.u_wallace._3378_ ),
    .C1(\u_cpu.ALU.u_wallace._3379_ ),
    .Y(\u_cpu.ALU.u_wallace._3380_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8927_  (.A1(\u_cpu.ALU.u_wallace._3140_ ),
    .A2(\u_cpu.ALU.u_wallace._3142_ ),
    .B1(\u_cpu.ALU.u_wallace._3143_ ),
    .C1(\u_cpu.ALU.u_wallace._3149_ ),
    .X(\u_cpu.ALU.u_wallace._3381_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8928_  (.A1(\u_cpu.ALU.u_wallace._3162_ ),
    .A2(\u_cpu.ALU.u_wallace._3158_ ),
    .B1(\u_cpu.ALU.u_wallace._3381_ ),
    .Y(\u_cpu.ALU.u_wallace._3383_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._8929_  (.A1(\u_cpu.ALU.u_wallace._3377_ ),
    .A2(\u_cpu.ALU.u_wallace._3380_ ),
    .A3(\u_cpu.ALU.u_wallace._3383_ ),
    .B1(\u_cpu.ALU.u_wallace._3223_ ),
    .B2(\u_cpu.ALU.u_wallace._3220_ ),
    .X(\u_cpu.ALU.u_wallace._3384_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8930_  (.A(\u_cpu.ALU.u_wallace._3376_ ),
    .B(\u_cpu.ALU.u_wallace._3378_ ),
    .C(\u_cpu.ALU.u_wallace._3379_ ),
    .Y(\u_cpu.ALU.u_wallace._3385_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8931_  (.A1(\u_cpu.ALU.u_wallace._3374_ ),
    .A2(\u_cpu.ALU.u_wallace._3375_ ),
    .B1(\u_cpu.ALU.u_wallace._3357_ ),
    .B2(\u_cpu.ALU.u_wallace._3359_ ),
    .Y(\u_cpu.ALU.u_wallace._3386_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8932_  (.A1(\u_cpu.ALU.u_wallace._3381_ ),
    .A2(\u_cpu.ALU.u_wallace._3159_ ),
    .B1(\u_cpu.ALU.u_wallace._3385_ ),
    .C1(\u_cpu.ALU.u_wallace._3386_ ),
    .X(\u_cpu.ALU.u_wallace._3387_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8933_  (.A(\u_cpu.ALU.u_wallace._3377_ ),
    .B(\u_cpu.ALU.u_wallace._3380_ ),
    .C(\u_cpu.ALU.u_wallace._3383_ ),
    .Y(\u_cpu.ALU.u_wallace._3388_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8934_  (.A1(\u_cpu.ALU.u_wallace._3381_ ),
    .A2(\u_cpu.ALU.u_wallace._3159_ ),
    .B1(\u_cpu.ALU.u_wallace._3385_ ),
    .C1(\u_cpu.ALU.u_wallace._3386_ ),
    .Y(\u_cpu.ALU.u_wallace._3389_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8935_  (.A1(\u_cpu.ALU.u_wallace._3219_ ),
    .A2(\u_cpu.ALU.u_wallace._3222_ ),
    .B1(\u_cpu.ALU.u_wallace._3216_ ),
    .X(\u_cpu.ALU.u_wallace._3390_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8936_  (.A1(\u_cpu.ALU.u_wallace._3388_ ),
    .A2(\u_cpu.ALU.u_wallace._3389_ ),
    .B1(\u_cpu.ALU.u_wallace._3390_ ),
    .X(\u_cpu.ALU.u_wallace._3391_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._8937_  (.A1(\u_cpu.ALU.u_wallace._3101_ ),
    .A2(\u_cpu.ALU.u_wallace._3102_ ),
    .B1(\u_cpu.ALU.u_wallace._3104_ ),
    .X(\u_cpu.ALU.u_wallace._3392_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._8938_  (.A1(\u_cpu.ALU.u_wallace._4934_ ),
    .A2(\u_cpu.ALU.u_wallace._3060_ ),
    .A3(\u_cpu.ALU.u_wallace._3061_ ),
    .B1(\u_cpu.ALU.u_wallace._3057_ ),
    .X(\u_cpu.ALU.u_wallace._3394_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8939_  (.A(\u_cpu.ALU.u_wallace._1826_ ),
    .B(\u_cpu.ALU.u_wallace._4653_ ),
    .C(\u_cpu.ALU.u_wallace._0629_ ),
    .Y(\u_cpu.ALU.u_wallace._3395_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._8940_  (.A(\u_cpu.ALU.u_wallace._0075_ ),
    .B(\u_cpu.ALU.SrcA[28] ),
    .X(\u_cpu.ALU.u_wallace._3396_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8941_  (.A1(\u_cpu.ALU.u_wallace._4647_ ),
    .A2(\u_cpu.ALU.u_wallace._1102_ ),
    .B1(\u_cpu.ALU.u_wallace._1734_ ),
    .B2(\u_cpu.ALU.u_wallace._1771_ ),
    .X(\u_cpu.ALU.u_wallace._3397_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8942_  (.A1(\u_cpu.ALU.u_wallace._1737_ ),
    .A2(\u_cpu.ALU.u_wallace._3395_ ),
    .B1(\u_cpu.ALU.u_wallace._3396_ ),
    .C1(\u_cpu.ALU.u_wallace._3397_ ),
    .Y(\u_cpu.ALU.u_wallace._3398_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8943_  (.A(\u_cpu.ALU.SrcA[28] ),
    .X(\u_cpu.ALU.u_wallace._3399_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._8944_  (.A(\u_cpu.ALU.u_wallace._3399_ ),
    .Y(\u_cpu.ALU.u_wallace._3400_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8945_  (.A1(\u_cpu.ALU.u_wallace._4653_ ),
    .A2(\u_cpu.ALU.u_wallace._0629_ ),
    .B1(\u_cpu.ALU.u_wallace._1734_ ),
    .B2(\u_cpu.ALU.u_wallace._1826_ ),
    .Y(\u_cpu.ALU.u_wallace._3401_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8946_  (.A(\u_cpu.ALU.u_wallace._4645_ ),
    .B(\u_cpu.ALU.u_wallace._4797_ ),
    .C(\u_cpu.ALU.u_wallace._0639_ ),
    .D(\u_cpu.ALU.SrcA[22] ),
    .X(\u_cpu.ALU.u_wallace._3402_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8947_  (.A1(\u_cpu.ALU.u_wallace._4923_ ),
    .A2(\u_cpu.ALU.u_wallace._3400_ ),
    .B1(\u_cpu.ALU.u_wallace._3401_ ),
    .B2(\u_cpu.ALU.u_wallace._3402_ ),
    .Y(\u_cpu.ALU.u_wallace._3403_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8948_  (.A(\u_cpu.ALU.u_wallace._3398_ ),
    .B(\u_cpu.ALU.u_wallace._3403_ ),
    .Y(\u_cpu.ALU.u_wallace._3405_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8949_  (.A(\u_cpu.ALU.u_wallace._0187_ ),
    .B(\u_cpu.ALU.u_wallace._0304_ ),
    .C(\u_cpu.ALU.SrcA[26] ),
    .D(\u_cpu.ALU.SrcA[27] ),
    .Y(\u_cpu.ALU.u_wallace._3406_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8950_  (.A1(\u_cpu.ALU.u_wallace._1169_ ),
    .A2(\u_cpu.ALU.SrcA[26] ),
    .B1(\u_cpu.ALU.SrcA[27] ),
    .B2(\u_cpu.ALU.u_wallace._1158_ ),
    .X(\u_cpu.ALU.u_wallace._3407_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8951_  (.A(\u_cpu.ALU.u_wallace._0468_ ),
    .B(\u_cpu.ALU.u_wallace._2578_ ),
    .Y(\u_cpu.ALU.u_wallace._3408_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8952_  (.A1(\u_cpu.ALU.u_wallace._3406_ ),
    .A2(\u_cpu.ALU.u_wallace._3407_ ),
    .B1(\u_cpu.ALU.u_wallace._3408_ ),
    .X(\u_cpu.ALU.u_wallace._3409_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._8953_  (.A1(\u_cpu.ALU.u_wallace._4678_ ),
    .A2(\u_cpu.ALU.u_wallace._2580_ ),
    .B1(\u_cpu.ALU.u_wallace._3406_ ),
    .C1(\u_cpu.ALU.u_wallace._3407_ ),
    .Y(\u_cpu.ALU.u_wallace._3410_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8954_  (.A1(\u_cpu.ALU.u_wallace._3409_ ),
    .A2(\u_cpu.ALU.u_wallace._3410_ ),
    .B1(\u_cpu.ALU.u_wallace._3405_ ),
    .B2(\u_cpu.ALU.u_wallace._3394_ ),
    .Y(\u_cpu.ALU.u_wallace._3411_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8955_  (.A1(\u_cpu.ALU.u_wallace._3394_ ),
    .A2(\u_cpu.ALU.u_wallace._3405_ ),
    .B1(\u_cpu.ALU.u_wallace._3411_ ),
    .Y(\u_cpu.ALU.u_wallace._3412_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8956_  (.A(\u_cpu.ALU.u_wallace._2779_ ),
    .B(\u_cpu.ALU.u_wallace._1531_ ),
    .Y(\u_cpu.ALU.u_wallace._3413_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8957_  (.A(\u_cpu.ALU.u_wallace._4554_ ),
    .B(\u_cpu.ALU.u_wallace._0629_ ),
    .Y(\u_cpu.ALU.u_wallace._3414_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8958_  (.A1(\u_cpu.ALU.u_wallace._3413_ ),
    .A2(\u_cpu.ALU.u_wallace._3414_ ),
    .B1(\u_cpu.ALU.u_wallace._3079_ ),
    .Y(\u_cpu.ALU.u_wallace._3416_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8959_  (.A1(\u_cpu.ALU.u_wallace._3062_ ),
    .A2(\u_cpu.ALU.u_wallace._3416_ ),
    .B1(\u_cpu.ALU.u_wallace._3398_ ),
    .C1(\u_cpu.ALU.u_wallace._3403_ ),
    .X(\u_cpu.ALU.u_wallace._3417_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8960_  (.A1(\u_cpu.ALU.u_wallace._3056_ ),
    .A2(\u_cpu.ALU.u_wallace._3058_ ),
    .A3(\u_cpu.ALU.u_wallace._0884_ ),
    .B1(\u_cpu.ALU.u_wallace._3062_ ),
    .X(\u_cpu.ALU.u_wallace._3418_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8961_  (.A1(\u_cpu.ALU.u_wallace._3398_ ),
    .A2(\u_cpu.ALU.u_wallace._3403_ ),
    .B1(\u_cpu.ALU.u_wallace._3418_ ),
    .Y(\u_cpu.ALU.u_wallace._3419_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8962_  (.A(\u_cpu.ALU.u_wallace._3409_ ),
    .B(\u_cpu.ALU.u_wallace._3410_ ),
    .Y(\u_cpu.ALU.u_wallace._3420_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._8963_  (.A1(\u_cpu.ALU.u_wallace._3417_ ),
    .A2(\u_cpu.ALU.u_wallace._3419_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3420_ ),
    .Y(\u_cpu.ALU.u_wallace._3421_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8964_  (.A1(\u_cpu.ALU.u_wallace._3072_ ),
    .A2(\u_cpu.ALU.u_wallace._3067_ ),
    .B1(\u_cpu.ALU.u_wallace._3077_ ),
    .Y(\u_cpu.ALU.u_wallace._3422_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._8965_  (.A1(\u_cpu.ALU.u_wallace._3412_ ),
    .A2(\u_cpu.ALU.u_wallace._3421_ ),
    .B1(\u_cpu.ALU.u_wallace._3422_ ),
    .X(\u_cpu.ALU.u_wallace._3423_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8966_  (.A1(\u_cpu.ALU.u_wallace._2187_ ),
    .A2(\u_cpu.ALU.u_wallace._2002_ ),
    .B1(\u_cpu.ALU.u_wallace._2222_ ),
    .B2(\u_cpu.ALU.u_wallace._2155_ ),
    .X(\u_cpu.ALU.u_wallace._3424_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8967_  (.A(\u_cpu.ALU.u_wallace._1476_ ),
    .B(\u_cpu.ALU.u_wallace._1508_ ),
    .C(\u_cpu.ALU.u_wallace._2002_ ),
    .D(\u_cpu.ALU.u_wallace._2222_ ),
    .Y(\u_cpu.ALU.u_wallace._3425_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8968_  (.A1(\u_cpu.ALU.u_wallace._4542_ ),
    .A2(\u_cpu.ALU.u_wallace._2618_ ),
    .B1(\u_cpu.ALU.u_wallace._3424_ ),
    .B2(\u_cpu.ALU.u_wallace._3425_ ),
    .Y(\u_cpu.ALU.u_wallace._3427_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8969_  (.A1(\u_cpu.ALU.u_wallace._1508_ ),
    .A2(\u_cpu.ALU.u_wallace._2002_ ),
    .B1(\u_cpu.ALU.u_wallace._2222_ ),
    .B2(\u_cpu.ALU.u_wallace._1476_ ),
    .Y(\u_cpu.ALU.u_wallace._3428_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8970_  (.A(\u_cpu.ALU.u_wallace._2604_ ),
    .B(\u_cpu.ALU.u_wallace._1531_ ),
    .Y(\u_cpu.ALU.u_wallace._3429_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8971_  (.A(\u_cpu.ALU.u_wallace._2155_ ),
    .B(\u_cpu.ALU.u_wallace._1552_ ),
    .C(\u_cpu.ALU.u_wallace._2000_ ),
    .D(\u_cpu.ALU.u_wallace._2226_ ),
    .X(\u_cpu.ALU.u_wallace._3430_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._8972_  (.A(\u_cpu.ALU.u_wallace._3428_ ),
    .B(\u_cpu.ALU.u_wallace._3429_ ),
    .C(\u_cpu.ALU.u_wallace._3430_ ),
    .Y(\u_cpu.ALU.u_wallace._3431_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8973_  (.A(\u_cpu.ALU.u_wallace._0578_ ),
    .B(\u_cpu.ALU.u_wallace._2222_ ),
    .Y(\u_cpu.ALU.u_wallace._3432_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8974_  (.A1(\u_cpu.ALU.u_wallace._4796_ ),
    .A2(\u_cpu.ALU.u_wallace._2578_ ),
    .B1(\u_cpu.ALU.u_wallace._2869_ ),
    .B2(\u_cpu.ALU.u_wallace._0217_ ),
    .Y(\u_cpu.ALU.u_wallace._3433_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._8975_  (.A1(\u_cpu.ALU.u_wallace._3432_ ),
    .A2(\u_cpu.ALU.u_wallace._3433_ ),
    .B1(\u_cpu.ALU.u_wallace._3068_ ),
    .Y(\u_cpu.ALU.u_wallace._3434_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._8976_  (.A1(\u_cpu.ALU.u_wallace._3427_ ),
    .A2(\u_cpu.ALU.u_wallace._3431_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3434_ ),
    .Y(\u_cpu.ALU.u_wallace._3435_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._8977_  (.A1(\u_cpu.ALU.u_wallace._4542_ ),
    .A2(\u_cpu.ALU.u_wallace._2618_ ),
    .B1(\u_cpu.ALU.u_wallace._3424_ ),
    .B2(\u_cpu.ALU.u_wallace._3425_ ),
    .X(\u_cpu.ALU.u_wallace._3436_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._8978_  (.A(\u_cpu.ALU.u_wallace._3424_ ),
    .B(\u_cpu.ALU.u_wallace._3425_ ),
    .C(\u_cpu.ALU.u_wallace._0015_ ),
    .D(\u_cpu.ALU.u_wallace._2618_ ),
    .Y(\u_cpu.ALU.u_wallace._3438_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8979_  (.A(\u_cpu.ALU.u_wallace._3434_ ),
    .B(\u_cpu.ALU.u_wallace._3436_ ),
    .C(\u_cpu.ALU.u_wallace._3438_ ),
    .Y(\u_cpu.ALU.u_wallace._3439_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._8980_  (.A1(\u_cpu.ALU.u_wallace._3087_ ),
    .A2(\u_cpu.ALU.u_wallace._3088_ ),
    .A3(\u_cpu.ALU.u_wallace._0015_ ),
    .B1(\u_cpu.ALU.u_wallace._3096_ ),
    .X(\u_cpu.ALU.u_wallace._3440_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8981_  (.A1(\u_cpu.ALU.u_wallace._3435_ ),
    .A2(\u_cpu.ALU.u_wallace._3439_ ),
    .B1(\u_cpu.ALU.u_wallace._3440_ ),
    .Y(\u_cpu.ALU.u_wallace._3441_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8982_  (.A(\u_cpu.ALU.u_wallace._3440_ ),
    .B(\u_cpu.ALU.u_wallace._3435_ ),
    .C(\u_cpu.ALU.u_wallace._3439_ ),
    .X(\u_cpu.ALU.u_wallace._3442_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._8983_  (.A(\u_cpu.ALU.u_wallace._3441_ ),
    .B(\u_cpu.ALU.u_wallace._3442_ ),
    .Y(\u_cpu.ALU.u_wallace._3443_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8984_  (.A(\u_cpu.ALU.u_wallace._3063_ ),
    .B(\u_cpu.ALU.u_wallace._3059_ ),
    .Y(\u_cpu.ALU.u_wallace._3444_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8985_  (.A1(\u_cpu.ALU.u_wallace._3444_ ),
    .A2(\u_cpu.ALU.u_wallace._3081_ ),
    .B1(\u_cpu.ALU.u_wallace._3072_ ),
    .Y(\u_cpu.ALU.u_wallace._3445_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._8986_  (.A(\u_cpu.ALU.u_wallace._0187_ ),
    .B(\u_cpu.ALU.u_wallace._4796_ ),
    .C(\u_cpu.ALU.SrcA[26] ),
    .D(\u_cpu.ALU.SrcA[27] ),
    .X(\u_cpu.ALU.u_wallace._3446_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._8987_  (.A1(\u_cpu.ALU.u_wallace._4796_ ),
    .A2(\u_cpu.ALU.u_wallace._2869_ ),
    .B1(\u_cpu.ALU.u_wallace._3058_ ),
    .B2(\u_cpu.ALU.u_wallace._0217_ ),
    .Y(\u_cpu.ALU.u_wallace._3447_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._8988_  (.A(\u_cpu.ALU.u_wallace._2578_ ),
    .X(\u_cpu.ALU.u_wallace._3449_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8989_  (.A1(\u_cpu.ALU.u_wallace._3446_ ),
    .A2(\u_cpu.ALU.u_wallace._3447_ ),
    .B1(\u_cpu.ALU.u_wallace._4663_ ),
    .C1(\u_cpu.ALU.u_wallace._3449_ ),
    .X(\u_cpu.ALU.u_wallace._3450_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._8990_  (.A(\u_cpu.ALU.u_wallace._3408_ ),
    .B(\u_cpu.ALU.u_wallace._3406_ ),
    .C(\u_cpu.ALU.u_wallace._3407_ ),
    .X(\u_cpu.ALU.u_wallace._3451_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._8991_  (.A1_N(\u_cpu.ALU.u_wallace._3394_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3405_ ),
    .B1(\u_cpu.ALU.u_wallace._3450_ ),
    .B2(\u_cpu.ALU.u_wallace._3451_ ),
    .Y(\u_cpu.ALU.u_wallace._3452_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._8992_  (.A1(\u_cpu.ALU.u_wallace._3065_ ),
    .A2(\u_cpu.ALU.u_wallace._3445_ ),
    .B1(\u_cpu.ALU.u_wallace._3417_ ),
    .B2(\u_cpu.ALU.u_wallace._3452_ ),
    .C1(\u_cpu.ALU.u_wallace._3421_ ),
    .Y(\u_cpu.ALU.u_wallace._3453_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._8993_  (.A(\u_cpu.ALU.u_wallace._3423_ ),
    .B(\u_cpu.ALU.u_wallace._3443_ ),
    .C(\u_cpu.ALU.u_wallace._3453_ ),
    .Y(\u_cpu.ALU.u_wallace._3454_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._8994_  (.A1(\u_cpu.ALU.u_wallace._3065_ ),
    .A2(\u_cpu.ALU.u_wallace._3445_ ),
    .B1(\u_cpu.ALU.u_wallace._3417_ ),
    .B2(\u_cpu.ALU.u_wallace._3452_ ),
    .C1(\u_cpu.ALU.u_wallace._3421_ ),
    .X(\u_cpu.ALU.u_wallace._3455_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._8995_  (.A1(\u_cpu.ALU.u_wallace._3412_ ),
    .A2(\u_cpu.ALU.u_wallace._3421_ ),
    .B1(\u_cpu.ALU.u_wallace._3422_ ),
    .Y(\u_cpu.ALU.u_wallace._3456_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._8996_  (.A1(\u_cpu.ALU.u_wallace._3441_ ),
    .A2(\u_cpu.ALU.u_wallace._3442_ ),
    .B1(\u_cpu.ALU.u_wallace._3455_ ),
    .B2(\u_cpu.ALU.u_wallace._3456_ ),
    .Y(\u_cpu.ALU.u_wallace._3457_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._8997_  (.A1(\u_cpu.ALU.u_wallace._3084_ ),
    .A2(\u_cpu.ALU.u_wallace._3392_ ),
    .B1(\u_cpu.ALU.u_wallace._3454_ ),
    .C1(\u_cpu.ALU.u_wallace._3457_ ),
    .X(\u_cpu.ALU.u_wallace._3458_ ));
 sky130_fd_sc_hd__a32oi_2 \u_cpu.ALU.u_wallace._8998_  (.A1(\u_cpu.ALU.u_wallace._3085_ ),
    .A2(\u_cpu.ALU.u_wallace._3090_ ),
    .A3(\u_cpu.ALU.u_wallace._3091_ ),
    .B1(\u_cpu.ALU.u_wallace._3099_ ),
    .B2(\u_cpu.ALU.u_wallace._3110_ ),
    .Y(\u_cpu.ALU.u_wallace._3460_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._8999_  (.A(\u_cpu.ALU.u_wallace._4610_ ),
    .B(\u_cpu.ALU.u_wallace._1286_ ),
    .Y(\u_cpu.ALU.u_wallace._3461_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9000_  (.A(\u_cpu.ALU.u_wallace._3461_ ),
    .B(\u_cpu.ALU.u_wallace._3125_ ),
    .Y(\u_cpu.ALU.u_wallace._3462_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9001_  (.A1(\u_cpu.ALU.u_wallace._4302_ ),
    .A2(\u_cpu.ALU.u_wallace._1101_ ),
    .B1(\u_cpu.ALU.u_wallace._1275_ ),
    .B2(\u_cpu.ALU.u_wallace._4018_ ),
    .X(\u_cpu.ALU.u_wallace._3463_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9002_  (.A(\u_cpu.ALU.u_wallace._4717_ ),
    .B(\u_cpu.ALU.u_wallace._4599_ ),
    .C(\u_cpu.ALU.u_wallace._1101_ ),
    .D(\u_cpu.ALU.u_wallace._1275_ ),
    .Y(\u_cpu.ALU.u_wallace._3464_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9003_  (.A(\u_cpu.ALU.u_wallace._3463_ ),
    .B(\u_cpu.ALU.u_wallace._3464_ ),
    .C(\u_cpu.ALU.u_wallace._4610_ ),
    .D(\u_cpu.ALU.u_wallace._2916_ ),
    .Y(\u_cpu.ALU.u_wallace._3465_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._9004_  (.A1_N(\u_cpu.ALU.u_wallace._3463_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3464_ ),
    .B1(\u_cpu.ALU.u_wallace._4602_ ),
    .B2(\u_cpu.ALU.u_wallace._0809_ ),
    .Y(\u_cpu.ALU.u_wallace._3466_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9005_  (.A1(\u_cpu.ALU.u_wallace._3126_ ),
    .A2(\u_cpu.ALU.u_wallace._3462_ ),
    .B1(\u_cpu.ALU.u_wallace._3465_ ),
    .C1(\u_cpu.ALU.u_wallace._3466_ ),
    .X(\u_cpu.ALU.u_wallace._3467_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._9006_  (.A1(\u_cpu.ALU.u_wallace._3128_ ),
    .A2(\u_cpu.ALU.u_wallace._2621_ ),
    .A3(\u_cpu.ALU.u_wallace._4605_ ),
    .B1(\u_cpu.ALU.u_wallace._3126_ ),
    .X(\u_cpu.ALU.u_wallace._3468_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9007_  (.A1(\u_cpu.ALU.u_wallace._3465_ ),
    .A2(\u_cpu.ALU.u_wallace._3466_ ),
    .B1(\u_cpu.ALU.u_wallace._3468_ ),
    .Y(\u_cpu.ALU.u_wallace._3469_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9008_  (.A1(\u_cpu.ALU.u_wallace._4842_ ),
    .A2(\u_cpu.ALU.u_wallace._0850_ ),
    .B1(\u_cpu.ALU.u_wallace._1286_ ),
    .B2(\u_cpu.ALU.u_wallace._4732_ ),
    .Y(\u_cpu.ALU.u_wallace._3471_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9009_  (.A(\u_cpu.ALU.u_wallace._4840_ ),
    .B(\u_cpu.ALU.u_wallace._4838_ ),
    .C(\u_cpu.ALU.u_wallace._0850_ ),
    .D(\u_cpu.ALU.u_wallace._0642_ ),
    .X(\u_cpu.ALU.u_wallace._3472_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9010_  (.A1(\u_cpu.ALU.u_wallace._3471_ ),
    .A2(\u_cpu.ALU.u_wallace._3472_ ),
    .B1(\u_cpu.ALU.u_wallace._0034_ ),
    .C1(\u_cpu.ALU.u_wallace._1974_ ),
    .Y(\u_cpu.ALU.u_wallace._3473_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._9011_  (.A1(\u_cpu.ALU.u_wallace._0034_ ),
    .A2(\u_cpu.ALU.u_wallace._1974_ ),
    .B1(\u_cpu.ALU.u_wallace._3471_ ),
    .C1(\u_cpu.ALU.u_wallace._3472_ ),
    .X(\u_cpu.ALU.u_wallace._3474_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9012_  (.A(\u_cpu.ALU.u_wallace._3473_ ),
    .B(\u_cpu.ALU.u_wallace._3474_ ),
    .Y(\u_cpu.ALU.u_wallace._3475_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9013_  (.A1(\u_cpu.ALU.u_wallace._3467_ ),
    .A2(\u_cpu.ALU.u_wallace._3469_ ),
    .B1(\u_cpu.ALU.u_wallace._3475_ ),
    .Y(\u_cpu.ALU.u_wallace._3476_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9014_  (.A1(\u_cpu.ALU.u_wallace._3126_ ),
    .A2(\u_cpu.ALU.u_wallace._3462_ ),
    .B1(\u_cpu.ALU.u_wallace._3465_ ),
    .C1(\u_cpu.ALU.u_wallace._3466_ ),
    .Y(\u_cpu.ALU.u_wallace._3477_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9015_  (.A1(\u_cpu.ALU.u_wallace._3465_ ),
    .A2(\u_cpu.ALU.u_wallace._3466_ ),
    .B1(\u_cpu.ALU.u_wallace._3468_ ),
    .X(\u_cpu.ALU.u_wallace._3478_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._9016_  (.A_N(\u_cpu.ALU.u_wallace._3475_ ),
    .B(\u_cpu.ALU.u_wallace._3477_ ),
    .C(\u_cpu.ALU.u_wallace._3478_ ),
    .Y(\u_cpu.ALU.u_wallace._3479_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9017_  (.A(\u_cpu.ALU.u_wallace._3460_ ),
    .B(\u_cpu.ALU.u_wallace._3476_ ),
    .C(\u_cpu.ALU.u_wallace._3479_ ),
    .Y(\u_cpu.ALU.u_wallace._3480_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._9018_  (.A1(\u_cpu.ALU.u_wallace._3085_ ),
    .A2(\u_cpu.ALU.u_wallace._3090_ ),
    .A3(\u_cpu.ALU.u_wallace._3091_ ),
    .B1(\u_cpu.ALU.u_wallace._3099_ ),
    .B2(\u_cpu.ALU.u_wallace._3110_ ),
    .X(\u_cpu.ALU.u_wallace._3482_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9019_  (.A(\u_cpu.ALU.u_wallace._3475_ ),
    .B(\u_cpu.ALU.u_wallace._3477_ ),
    .C(\u_cpu.ALU.u_wallace._3478_ ),
    .Y(\u_cpu.ALU.u_wallace._3483_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9020_  (.A1(\u_cpu.ALU.u_wallace._3467_ ),
    .A2(\u_cpu.ALU.u_wallace._3469_ ),
    .B1(\u_cpu.ALU.u_wallace._3473_ ),
    .C1(\u_cpu.ALU.u_wallace._3474_ ),
    .Y(\u_cpu.ALU.u_wallace._3484_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9021_  (.A1(\u_cpu.ALU.u_wallace._3153_ ),
    .A2(\u_cpu.ALU.u_wallace._3156_ ),
    .B1(\u_cpu.ALU.u_wallace._3147_ ),
    .Y(\u_cpu.ALU.u_wallace._3485_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._9022_  (.A1(\u_cpu.ALU.u_wallace._3482_ ),
    .A2(\u_cpu.ALU.u_wallace._3483_ ),
    .A3(\u_cpu.ALU.u_wallace._3484_ ),
    .B1(\u_cpu.ALU.u_wallace._3485_ ),
    .Y(\u_cpu.ALU.u_wallace._3486_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9023_  (.A(\u_cpu.ALU.u_wallace._3482_ ),
    .B(\u_cpu.ALU.u_wallace._3483_ ),
    .C(\u_cpu.ALU.u_wallace._3484_ ),
    .Y(\u_cpu.ALU.u_wallace._3487_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._9024_  (.A1(\u_cpu.ALU.u_wallace._3127_ ),
    .A2(\u_cpu.ALU.u_wallace._3131_ ),
    .A3(\u_cpu.ALU.u_wallace._3132_ ),
    .B1(\u_cpu.ALU.u_wallace._3156_ ),
    .B2(\u_cpu.ALU.u_wallace._3153_ ),
    .X(\u_cpu.ALU.u_wallace._3488_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9025_  (.A1(\u_cpu.ALU.u_wallace._3487_ ),
    .A2(\u_cpu.ALU.u_wallace._3480_ ),
    .B1(\u_cpu.ALU.u_wallace._3488_ ),
    .Y(\u_cpu.ALU.u_wallace._3489_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9026_  (.A1(\u_cpu.ALU.u_wallace._3480_ ),
    .A2(\u_cpu.ALU.u_wallace._3486_ ),
    .B1(\u_cpu.ALU.u_wallace._3489_ ),
    .Y(\u_cpu.ALU.u_wallace._3490_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9027_  (.A1(\u_cpu.ALU.u_wallace._3455_ ),
    .A2(\u_cpu.ALU.u_wallace._3456_ ),
    .B1(\u_cpu.ALU.u_wallace._3443_ ),
    .Y(\u_cpu.ALU.u_wallace._3491_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9028_  (.A1(\u_cpu.ALU.u_wallace._3441_ ),
    .A2(\u_cpu.ALU.u_wallace._3442_ ),
    .B1(\u_cpu.ALU.u_wallace._3453_ ),
    .C1(\u_cpu.ALU.u_wallace._3423_ ),
    .Y(\u_cpu.ALU.u_wallace._3493_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9029_  (.A(\u_cpu.ALU.u_wallace._3092_ ),
    .B(\u_cpu.ALU.u_wallace._3099_ ),
    .Y(\u_cpu.ALU.u_wallace._3494_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9030_  (.A1(\u_cpu.ALU.u_wallace._3100_ ),
    .A2(\u_cpu.ALU.u_wallace._3494_ ),
    .B1(\u_cpu.ALU.u_wallace._3109_ ),
    .Y(\u_cpu.ALU.u_wallace._3495_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9031_  (.A1(\u_cpu.ALU.u_wallace._3495_ ),
    .A2(\u_cpu.ALU.u_wallace._3104_ ),
    .B1(\u_cpu.ALU.u_wallace._3084_ ),
    .Y(\u_cpu.ALU.u_wallace._3496_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9032_  (.A(\u_cpu.ALU.u_wallace._3491_ ),
    .B(\u_cpu.ALU.u_wallace._3493_ ),
    .C(\u_cpu.ALU.u_wallace._3496_ ),
    .Y(\u_cpu.ALU.u_wallace._3497_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9033_  (.A(\u_cpu.ALU.u_wallace._3490_ ),
    .B(\u_cpu.ALU.u_wallace._3497_ ),
    .Y(\u_cpu.ALU.u_wallace._3498_ ));
 sky130_fd_sc_hd__a311oi_2 \u_cpu.ALU.u_wallace._9034_  (.A1(\u_cpu.ALU.u_wallace._3120_ ),
    .A2(\u_cpu.ALU.u_wallace._3121_ ),
    .A3(\u_cpu.ALU.u_wallace._3123_ ),
    .B1(\u_cpu.ALU.u_wallace._3164_ ),
    .C1(\u_cpu.ALU.u_wallace._3169_ ),
    .Y(\u_cpu.ALU.u_wallace._3499_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9035_  (.A1(\u_cpu.ALU.u_wallace._3487_ ),
    .A2(\u_cpu.ALU.u_wallace._3480_ ),
    .B1(\u_cpu.ALU.u_wallace._3488_ ),
    .X(\u_cpu.ALU.u_wallace._3500_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9036_  (.A(\u_cpu.ALU.u_wallace._3488_ ),
    .B(\u_cpu.ALU.u_wallace._3487_ ),
    .C(\u_cpu.ALU.u_wallace._3480_ ),
    .Y(\u_cpu.ALU.u_wallace._3501_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9037_  (.A1(\u_cpu.ALU.u_wallace._3084_ ),
    .A2(\u_cpu.ALU.u_wallace._3392_ ),
    .B1(\u_cpu.ALU.u_wallace._3454_ ),
    .C1(\u_cpu.ALU.u_wallace._3457_ ),
    .Y(\u_cpu.ALU.u_wallace._3502_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9038_  (.A1(\u_cpu.ALU.u_wallace._3500_ ),
    .A2(\u_cpu.ALU.u_wallace._3501_ ),
    .B1(\u_cpu.ALU.u_wallace._3502_ ),
    .B2(\u_cpu.ALU.u_wallace._3497_ ),
    .X(\u_cpu.ALU.u_wallace._3504_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._9039_  (.A1(\u_cpu.ALU.u_wallace._3458_ ),
    .A2(\u_cpu.ALU.u_wallace._3498_ ),
    .B1(\u_cpu.ALU.u_wallace._3117_ ),
    .B2(\u_cpu.ALU.u_wallace._3499_ ),
    .C1(\u_cpu.ALU.u_wallace._3504_ ),
    .Y(\u_cpu.ALU.u_wallace._3505_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9040_  (.A(\u_cpu.ALU.u_wallace._3500_ ),
    .B(\u_cpu.ALU.u_wallace._3501_ ),
    .Y(\u_cpu.ALU.u_wallace._3506_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9041_  (.A1(\u_cpu.ALU.u_wallace._3502_ ),
    .A2(\u_cpu.ALU.u_wallace._3497_ ),
    .B1(\u_cpu.ALU.u_wallace._3506_ ),
    .X(\u_cpu.ALU.u_wallace._3507_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9042_  (.A(\u_cpu.ALU.u_wallace._3506_ ),
    .B(\u_cpu.ALU.u_wallace._3502_ ),
    .C(\u_cpu.ALU.u_wallace._3497_ ),
    .Y(\u_cpu.ALU.u_wallace._3508_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9043_  (.A1(\u_cpu.ALU.u_wallace._3124_ ),
    .A2(\u_cpu.ALU.u_wallace._3165_ ),
    .B1(\u_cpu.ALU.u_wallace._3117_ ),
    .Y(\u_cpu.ALU.u_wallace._3509_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9044_  (.A(\u_cpu.ALU.u_wallace._3507_ ),
    .B(\u_cpu.ALU.u_wallace._3508_ ),
    .C(\u_cpu.ALU.u_wallace._3509_ ),
    .Y(\u_cpu.ALU.u_wallace._3510_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._9045_  (.A1(\u_cpu.ALU.u_wallace._3384_ ),
    .A2(\u_cpu.ALU.u_wallace._3387_ ),
    .B1(\u_cpu.ALU.u_wallace._3391_ ),
    .C1(\u_cpu.ALU.u_wallace._3505_ ),
    .D1(\u_cpu.ALU.u_wallace._3510_ ),
    .Y(\u_cpu.ALU.u_wallace._3511_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9046_  (.A(\u_cpu.ALU.u_wallace._3390_ ),
    .B(\u_cpu.ALU.u_wallace._3388_ ),
    .C(\u_cpu.ALU.u_wallace._3389_ ),
    .Y(\u_cpu.ALU.u_wallace._3512_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9047_  (.A1(\u_cpu.ALU.u_wallace._3391_ ),
    .A2(\u_cpu.ALU.u_wallace._3512_ ),
    .B1(\u_cpu.ALU.u_wallace._3505_ ),
    .B2(\u_cpu.ALU.u_wallace._3510_ ),
    .X(\u_cpu.ALU.u_wallace._3513_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9048_  (.A1(\u_cpu.ALU.u_wallace._3245_ ),
    .A2(\u_cpu.ALU.u_wallace._3235_ ),
    .B1(\u_cpu.ALU.u_wallace._3511_ ),
    .C1(\u_cpu.ALU.u_wallace._3513_ ),
    .Y(\u_cpu.ALU.u_wallace._3515_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9049_  (.A1(\u_cpu.ALU.u_wallace._3241_ ),
    .A2(\u_cpu.ALU.u_wallace._3170_ ),
    .B1(\u_cpu.ALU.u_wallace._3236_ ),
    .Y(\u_cpu.ALU.u_wallace._3516_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9050_  (.A1(\u_cpu.ALU.u_wallace._3238_ ),
    .A2(\u_cpu.ALU.u_wallace._3239_ ),
    .B1(\u_cpu.ALU.u_wallace._3234_ ),
    .B2(\u_cpu.ALU.u_wallace._3516_ ),
    .Y(\u_cpu.ALU.u_wallace._3517_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9051_  (.A1(\u_cpu.ALU.u_wallace._3387_ ),
    .A2(\u_cpu.ALU.u_wallace._3384_ ),
    .B1(\u_cpu.ALU.u_wallace._3391_ ),
    .Y(\u_cpu.ALU.u_wallace._3518_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9052_  (.A1(\u_cpu.ALU.u_wallace._3505_ ),
    .A2(\u_cpu.ALU.u_wallace._3510_ ),
    .B1(\u_cpu.ALU.u_wallace._3518_ ),
    .X(\u_cpu.ALU.u_wallace._3519_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9053_  (.A(\u_cpu.ALU.u_wallace._3518_ ),
    .B(\u_cpu.ALU.u_wallace._3505_ ),
    .C(\u_cpu.ALU.u_wallace._3510_ ),
    .Y(\u_cpu.ALU.u_wallace._3520_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._9054_  (.A_N(\u_cpu.ALU.u_wallace._3517_ ),
    .B(\u_cpu.ALU.u_wallace._3519_ ),
    .C(\u_cpu.ALU.u_wallace._3520_ ),
    .Y(\u_cpu.ALU.u_wallace._3521_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._9055_  (.A1(\u_cpu.ALU.u_wallace._0414_ ),
    .A2(\u_cpu.ALU.u_wallace._2482_ ),
    .A3(\u_cpu.ALU.u_wallace._3255_ ),
    .B1(\u_cpu.ALU.u_wallace._3260_ ),
    .X(\u_cpu.ALU.u_wallace._3522_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9056_  (.A1(\u_cpu.ALU.u_wallace._4597_ ),
    .A2(\u_cpu.ALU.SrcB[26] ),
    .B1(\u_cpu.ALU.SrcB[27] ),
    .B2(\u_cpu.ALU.u_wallace._0261_ ),
    .Y(\u_cpu.ALU.u_wallace._3523_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9057_  (.A(\u_cpu.ALU.u_wallace._0359_ ),
    .B(\u_cpu.ALU.u_wallace._1454_ ),
    .C(\u_cpu.ALU.SrcB[26] ),
    .D(\u_cpu.ALU.SrcB[27] ),
    .X(\u_cpu.ALU.u_wallace._3524_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9058_  (.A1(\u_cpu.ALU.u_wallace._0621_ ),
    .A2(\u_cpu.ALU.u_wallace._2481_ ),
    .B1(\u_cpu.ALU.u_wallace._3523_ ),
    .B2(\u_cpu.ALU.u_wallace._3524_ ),
    .Y(\u_cpu.ALU.u_wallace._3526_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9059_  (.A(\u_cpu.ALU.u_wallace._4545_ ),
    .B(\u_cpu.ALU.u_wallace._4463_ ),
    .C(\u_cpu.ALU.u_wallace._3258_ ),
    .D(\u_cpu.ALU.u_wallace._3254_ ),
    .Y(\u_cpu.ALU.u_wallace._3527_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._9060_  (.A_N(\u_cpu.ALU.u_wallace._3523_ ),
    .B(\u_cpu.ALU.u_wallace._3527_ ),
    .C(\u_cpu.ALU.u_wallace._4541_ ),
    .D(\u_cpu.ALU.u_wallace._2480_ ),
    .Y(\u_cpu.ALU.u_wallace._3528_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9061_  (.A(\u_cpu.ALU.u_wallace._3526_ ),
    .B(\u_cpu.ALU.u_wallace._3528_ ),
    .Y(\u_cpu.ALU.u_wallace._3529_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.ALU.u_wallace._9062_  (.A1(\u_cpu.ALU.u_wallace._0414_ ),
    .A2(\u_cpu.ALU.u_wallace._2481_ ),
    .A3(\u_cpu.ALU.u_wallace._3255_ ),
    .B1(\u_cpu.ALU.u_wallace._3260_ ),
    .Y(\u_cpu.ALU.u_wallace._3530_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9063_  (.A(\u_cpu.ALU.u_wallace._3253_ ),
    .B(\u_cpu.ALU.u_wallace._2397_ ),
    .Y(\u_cpu.ALU.u_wallace._3531_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._9064_  (.A1(\u_cpu.ALU.u_wallace._3530_ ),
    .A2(\u_cpu.ALU.u_wallace._3526_ ),
    .A3(\u_cpu.ALU.u_wallace._3528_ ),
    .B1(\u_cpu.ALU.u_wallace._3531_ ),
    .X(\u_cpu.ALU.u_wallace._3532_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9065_  (.A1(\u_cpu.ALU.u_wallace._3522_ ),
    .A2(\u_cpu.ALU.u_wallace._3529_ ),
    .B1(\u_cpu.ALU.u_wallace._3532_ ),
    .Y(\u_cpu.ALU.u_wallace._3533_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9066_  (.A(\u_cpu.ALU.u_wallace._3530_ ),
    .B(\u_cpu.ALU.u_wallace._3526_ ),
    .C(\u_cpu.ALU.u_wallace._3528_ ),
    .Y(\u_cpu.ALU.u_wallace._3534_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9067_  (.A1(\u_cpu.ALU.u_wallace._3526_ ),
    .A2(\u_cpu.ALU.u_wallace._3528_ ),
    .B1(\u_cpu.ALU.u_wallace._3530_ ),
    .X(\u_cpu.ALU.u_wallace._3535_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9068_  (.A1(\u_cpu.ALU.u_wallace._3253_ ),
    .A2(\u_cpu.ALU.u_wallace._2397_ ),
    .B1(\u_cpu.ALU.u_wallace._3534_ ),
    .B2(\u_cpu.ALU.u_wallace._3535_ ),
    .Y(\u_cpu.ALU.u_wallace._3537_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9069_  (.A1(\u_cpu.ALU.u_wallace._3268_ ),
    .A2(\u_cpu.ALU.u_wallace._3269_ ),
    .B1(\u_cpu.ALU.u_wallace._3266_ ),
    .Y(\u_cpu.ALU.u_wallace._3538_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._9070_  (.A1(\u_cpu.ALU.u_wallace._3533_ ),
    .A2(\u_cpu.ALU.u_wallace._3537_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3538_ ),
    .Y(\u_cpu.ALU.u_wallace._3539_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU.u_wallace._9071_  (.A1(\u_cpu.ALU.u_wallace._0414_ ),
    .A2(\u_cpu.ALU.u_wallace._2482_ ),
    .A3(\u_cpu.ALU.u_wallace._3255_ ),
    .B1(\u_cpu.ALU.u_wallace._3260_ ),
    .C1(\u_cpu.ALU.u_wallace._3529_ ),
    .X(\u_cpu.ALU.u_wallace._3540_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9072_  (.A1(\u_cpu.ALU.u_wallace._3253_ ),
    .A2(\u_cpu.ALU.u_wallace._2402_ ),
    .B1(\u_cpu.ALU.u_wallace._3534_ ),
    .B2(\u_cpu.ALU.u_wallace._3535_ ),
    .X(\u_cpu.ALU.u_wallace._3541_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9073_  (.A1(\u_cpu.ALU.u_wallace._3532_ ),
    .A2(\u_cpu.ALU.u_wallace._3540_ ),
    .B1(\u_cpu.ALU.u_wallace._3538_ ),
    .C1(\u_cpu.ALU.u_wallace._3541_ ),
    .Y(\u_cpu.ALU.u_wallace._3542_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._9074_  (.A1_N(\u_cpu.ALU.u_wallace._3539_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3542_ ),
    .B1(\u_cpu.ALU.u_wallace._4813_ ),
    .B2(\u_cpu.ALU.u_wallace._2131_ ),
    .Y(\u_cpu.ALU.u_wallace._3543_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9075_  (.A(\u_cpu.ALU.u_wallace._4813_ ),
    .B(\u_cpu.ALU.u_wallace._2131_ ),
    .Y(\u_cpu.ALU.u_wallace._3544_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9076_  (.A(\u_cpu.ALU.u_wallace._3177_ ),
    .B(\u_cpu.ALU.u_wallace._3178_ ),
    .C(\u_cpu.ALU.u_wallace._2343_ ),
    .D(\u_cpu.ALU.u_wallace._1615_ ),
    .X(\u_cpu.ALU.u_wallace._3545_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9077_  (.A1(\u_cpu.ALU.u_wallace._3172_ ),
    .A2(\u_cpu.ALU.u_wallace._3176_ ),
    .B1(\u_cpu.ALU.u_wallace._3182_ ),
    .Y(\u_cpu.ALU.u_wallace._3546_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9078_  (.A1(\u_cpu.ALU.u_wallace._3545_ ),
    .A2(\u_cpu.ALU.u_wallace._3546_ ),
    .B1(\u_cpu.ALU.u_wallace._3190_ ),
    .B2(\u_cpu.ALU.u_wallace._3186_ ),
    .Y(\u_cpu.ALU.u_wallace._3548_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._9079_  (.A(\u_cpu.ALU.SrcB[28] ),
    .Y(\u_cpu.ALU.u_wallace._3549_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9080_  (.A(\u_cpu.ALU.u_wallace._0198_ ),
    .B(\u_cpu.ALU.u_wallace._1136_ ),
    .C(\u_cpu.ALU.SrcB[21] ),
    .D(\u_cpu.ALU.SrcB[22] ),
    .Y(\u_cpu.ALU.u_wallace._3550_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.ALU.u_wallace._9081_  (.A(\u_cpu.ALU.u_wallace._0032_ ),
    .B(\u_cpu.ALU.u_wallace._3549_ ),
    .C(\u_cpu.ALU.u_wallace._3550_ ),
    .X(\u_cpu.ALU.u_wallace._3551_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._9082_  (.A(\u_cpu.ALU.u_wallace._3551_ ),
    .X(\u_cpu.ALU.u_wallace._3552_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9083_  (.A1(\u_cpu.ALU.u_wallace._0043_ ),
    .A2(\u_cpu.ALU.u_wallace._3549_ ),
    .B1(\u_cpu.ALU.u_wallace._3550_ ),
    .Y(\u_cpu.ALU.u_wallace._3553_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9084_  (.A(\u_cpu.ALU.u_wallace._3548_ ),
    .B(\u_cpu.ALU.u_wallace._3552_ ),
    .C(\u_cpu.ALU.u_wallace._3553_ ),
    .Y(\u_cpu.ALU.u_wallace._3554_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9085_  (.A1(\u_cpu.ALU.u_wallace._3172_ ),
    .A2(\u_cpu.ALU.u_wallace._3176_ ),
    .B1(\u_cpu.ALU.u_wallace._3179_ ),
    .C1(\u_cpu.ALU.u_wallace._3182_ ),
    .Y(\u_cpu.ALU.u_wallace._3555_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9086_  (.A(\u_cpu.ALU.u_wallace._3552_ ),
    .B(\u_cpu.ALU.u_wallace._3553_ ),
    .Y(\u_cpu.ALU.u_wallace._3556_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9087_  (.A1(\u_cpu.ALU.u_wallace._3190_ ),
    .A2(\u_cpu.ALU.u_wallace._3186_ ),
    .B1(\u_cpu.ALU.u_wallace._3555_ ),
    .C1(\u_cpu.ALU.u_wallace._3556_ ),
    .Y(\u_cpu.ALU.u_wallace._3557_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9088_  (.A1(\u_cpu.ALU.u_wallace._3554_ ),
    .A2(\u_cpu.ALU.u_wallace._3557_ ),
    .B1(\u_cpu.ALU.u_wallace._3279_ ),
    .Y(\u_cpu.ALU.u_wallace._3559_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9089_  (.A(\u_cpu.ALU.u_wallace._3554_ ),
    .B(\u_cpu.ALU.u_wallace._3557_ ),
    .C(\u_cpu.ALU.u_wallace._3279_ ),
    .X(\u_cpu.ALU.u_wallace._3560_ ));
 sky130_fd_sc_hd__a311oi_2 \u_cpu.ALU.u_wallace._9090_  (.A1(\u_cpu.ALU.u_wallace._3539_ ),
    .A2(\u_cpu.ALU.u_wallace._3544_ ),
    .A3(\u_cpu.ALU.u_wallace._3542_ ),
    .B1(\u_cpu.ALU.u_wallace._3559_ ),
    .C1(\u_cpu.ALU.u_wallace._3560_ ),
    .Y(\u_cpu.ALU.u_wallace._3561_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9091_  (.A(\u_cpu.ALU.u_wallace._2787_ ),
    .B(\u_cpu.ALU.u_wallace._2789_ ),
    .C(\u_cpu.ALU.u_wallace._2791_ ),
    .X(\u_cpu.ALU.u_wallace._3562_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9092_  (.A1(\u_cpu.ALU.u_wallace._3562_ ),
    .A2(\u_cpu.ALU.u_wallace._2794_ ),
    .B1(\u_cpu.ALU.u_wallace._3554_ ),
    .B2(\u_cpu.ALU.u_wallace._3557_ ),
    .X(\u_cpu.ALU.u_wallace._3563_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9093_  (.A(\u_cpu.ALU.u_wallace._3554_ ),
    .B(\u_cpu.ALU.u_wallace._3557_ ),
    .C(\u_cpu.ALU.u_wallace._3562_ ),
    .D(\u_cpu.ALU.u_wallace._2794_ ),
    .Y(\u_cpu.ALU.u_wallace._3564_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9094_  (.A1(\u_cpu.ALU.u_wallace._3532_ ),
    .A2(\u_cpu.ALU.u_wallace._3540_ ),
    .B1(\u_cpu.ALU.u_wallace._3538_ ),
    .Y(\u_cpu.ALU.u_wallace._3565_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._9095_  (.A1(\u_cpu.ALU.u_wallace._3537_ ),
    .A2(\u_cpu.ALU.u_wallace._3565_ ),
    .B1(\u_cpu.ALU.u_wallace._1333_ ),
    .C1(\u_cpu.ALU.u_wallace._2134_ ),
    .D1(\u_cpu.ALU.u_wallace._3539_ ),
    .Y(\u_cpu.ALU.u_wallace._3566_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9096_  (.A1(\u_cpu.ALU.u_wallace._3563_ ),
    .A2(\u_cpu.ALU.u_wallace._3564_ ),
    .B1(\u_cpu.ALU.u_wallace._3543_ ),
    .B2(\u_cpu.ALU.u_wallace._3566_ ),
    .Y(\u_cpu.ALU.u_wallace._3567_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9097_  (.A1(\u_cpu.ALU.u_wallace._3543_ ),
    .A2(\u_cpu.ALU.u_wallace._3561_ ),
    .B1(\u_cpu.ALU.u_wallace._3567_ ),
    .Y(\u_cpu.ALU.u_wallace._3568_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9098_  (.A1(\u_cpu.ALU.u_wallace._3224_ ),
    .A2(\u_cpu.ALU.u_wallace._3248_ ),
    .B1(\u_cpu.ALU.u_wallace._3568_ ),
    .Y(\u_cpu.ALU.u_wallace._3570_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._9099_  (.A1(\u_cpu.ALU.u_wallace._2943_ ),
    .A2(\u_cpu.ALU.u_wallace._2836_ ),
    .A3(\u_cpu.ALU.u_wallace._2844_ ),
    .B1(\u_cpu.ALU.u_wallace._3046_ ),
    .X(\u_cpu.ALU.u_wallace._3571_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9100_  (.A1(\u_cpu.ALU.u_wallace._3571_ ),
    .A2(\u_cpu.ALU.u_wallace._2853_ ),
    .B1(\u_cpu.ALU.u_wallace._3226_ ),
    .X(\u_cpu.ALU.u_wallace._3572_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9101_  (.A1(\u_cpu.ALU.u_wallace._3539_ ),
    .A2(\u_cpu.ALU.u_wallace._3542_ ),
    .B1(\u_cpu.ALU.u_wallace._3544_ ),
    .Y(\u_cpu.ALU.u_wallace._3573_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9102_  (.A(\u_cpu.ALU.u_wallace._3563_ ),
    .B(\u_cpu.ALU.u_wallace._3564_ ),
    .C(\u_cpu.ALU.u_wallace._3566_ ),
    .Y(\u_cpu.ALU.u_wallace._3574_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9103_  (.A1(\u_cpu.ALU.u_wallace._3537_ ),
    .A2(\u_cpu.ALU.u_wallace._3565_ ),
    .B1(\u_cpu.ALU.u_wallace._3544_ ),
    .C1(\u_cpu.ALU.u_wallace._3539_ ),
    .X(\u_cpu.ALU.u_wallace._3575_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9104_  (.A1(\u_cpu.ALU.u_wallace._3559_ ),
    .A2(\u_cpu.ALU.u_wallace._3560_ ),
    .B1(\u_cpu.ALU.u_wallace._3573_ ),
    .B2(\u_cpu.ALU.u_wallace._3575_ ),
    .Y(\u_cpu.ALU.u_wallace._3576_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9105_  (.A1(\u_cpu.ALU.u_wallace._3573_ ),
    .A2(\u_cpu.ALU.u_wallace._3574_ ),
    .B1(\u_cpu.ALU.u_wallace._3576_ ),
    .Y(\u_cpu.ALU.u_wallace._3577_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9106_  (.A1(\u_cpu.ALU.u_wallace._3232_ ),
    .A2(\u_cpu.ALU.u_wallace._3231_ ),
    .B1(\u_cpu.ALU.u_wallace._3572_ ),
    .C1(\u_cpu.ALU.u_wallace._3577_ ),
    .Y(\u_cpu.ALU.u_wallace._3578_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._9107_  (.A1(\u_cpu.ALU.u_wallace._2556_ ),
    .A2(\u_cpu.ALU.u_wallace._2514_ ),
    .A3(\u_cpu.ALU.u_wallace._3280_ ),
    .B1(\u_cpu.ALU.u_wallace._3288_ ),
    .B2(\u_cpu.ALU.u_wallace._3277_ ),
    .X(\u_cpu.ALU.u_wallace._3579_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9108_  (.A1(\u_cpu.ALU.u_wallace._3570_ ),
    .A2(\u_cpu.ALU.u_wallace._3578_ ),
    .B1(\u_cpu.ALU.u_wallace._3579_ ),
    .Y(\u_cpu.ALU.u_wallace._3581_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU.u_wallace._9109_  (.A1(\u_cpu.ALU.u_wallace._3224_ ),
    .A2(\u_cpu.ALU.u_wallace._3248_ ),
    .A3(\u_cpu.ALU.u_wallace._3568_ ),
    .B1(\u_cpu.ALU.u_wallace._3570_ ),
    .C1(\u_cpu.ALU.u_wallace._3579_ ),
    .X(\u_cpu.ALU.u_wallace._3582_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9110_  (.A(\u_cpu.ALU.u_wallace._3581_ ),
    .B(\u_cpu.ALU.u_wallace._3582_ ),
    .Y(\u_cpu.ALU.u_wallace._3583_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9111_  (.A(\u_cpu.ALU.u_wallace._3515_ ),
    .B(\u_cpu.ALU.u_wallace._3521_ ),
    .C(\u_cpu.ALU.u_wallace._3583_ ),
    .Y(\u_cpu.ALU.u_wallace._3584_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.ALU.u_wallace._9112_  (.A1_N(\u_cpu.ALU.u_wallace._3581_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3582_ ),
    .B1(\u_cpu.ALU.u_wallace._3515_ ),
    .B2(\u_cpu.ALU.u_wallace._3521_ ),
    .X(\u_cpu.ALU.u_wallace._3585_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9113_  (.A1(\u_cpu.ALU.u_wallace._3301_ ),
    .A2(\u_cpu.ALU.u_wallace._3341_ ),
    .B1(\u_cpu.ALU.u_wallace._3584_ ),
    .C1(\u_cpu.ALU.u_wallace._3585_ ),
    .X(\u_cpu.ALU.u_wallace._3586_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._9114_  (.A(\u_cpu.ALU.u_wallace._3291_ ),
    .Y(\u_cpu.ALU.u_wallace._3587_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._9115_  (.A1(\u_cpu.ALU.u_wallace._2958_ ),
    .A2(\u_cpu.ALU.u_wallace._2808_ ),
    .A3(\u_cpu.ALU.u_wallace._3286_ ),
    .B1(\u_cpu.ALU.u_wallace._3292_ ),
    .Y(\u_cpu.ALU.u_wallace._3588_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._9116_  (.A1(\u_cpu.ALU.u_wallace._3340_ ),
    .A2(\u_cpu.ALU.u_wallace._3300_ ),
    .B1(\u_cpu.ALU.u_wallace._3252_ ),
    .X(\u_cpu.ALU.u_wallace._3589_ ));
 sky130_fd_sc_hd__a21bo_2 \u_cpu.ALU.u_wallace._9117_  (.A1(\u_cpu.ALU.u_wallace._3515_ ),
    .A2(\u_cpu.ALU.u_wallace._3521_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3583_ ),
    .X(\u_cpu.ALU.u_wallace._3590_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9118_  (.A1(\u_cpu.ALU.u_wallace._3581_ ),
    .A2(\u_cpu.ALU.u_wallace._3582_ ),
    .B1(\u_cpu.ALU.u_wallace._3515_ ),
    .C1(\u_cpu.ALU.u_wallace._3521_ ),
    .Y(\u_cpu.ALU.u_wallace._3592_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9119_  (.A(\u_cpu.ALU.u_wallace._3589_ ),
    .B(\u_cpu.ALU.u_wallace._3590_ ),
    .C(\u_cpu.ALU.u_wallace._3592_ ),
    .Y(\u_cpu.ALU.u_wallace._3593_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9120_  (.A1(\u_cpu.ALU.u_wallace._3587_ ),
    .A2(\u_cpu.ALU.u_wallace._3588_ ),
    .B1(\u_cpu.ALU.u_wallace._3593_ ),
    .Y(\u_cpu.ALU.u_wallace._3594_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9121_  (.A1(\u_cpu.ALU.u_wallace._3301_ ),
    .A2(\u_cpu.ALU.u_wallace._3341_ ),
    .B1(\u_cpu.ALU.u_wallace._3584_ ),
    .C1(\u_cpu.ALU.u_wallace._3585_ ),
    .Y(\u_cpu.ALU.u_wallace._3595_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU.u_wallace._9122_  (.A(\u_cpu.ALU.u_wallace._3587_ ),
    .B(\u_cpu.ALU.u_wallace._3588_ ),
    .X(\u_cpu.ALU.u_wallace._3596_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9123_  (.A1(\u_cpu.ALU.u_wallace._3595_ ),
    .A2(\u_cpu.ALU.u_wallace._3593_ ),
    .B1(\u_cpu.ALU.u_wallace._3596_ ),
    .X(\u_cpu.ALU.u_wallace._3597_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._9124_  (.A1(\u_cpu.ALU.u_wallace._3586_ ),
    .A2(\u_cpu.ALU.u_wallace._3594_ ),
    .B1(\u_cpu.ALU.u_wallace._3307_ ),
    .B2(\u_cpu.ALU.u_wallace._3318_ ),
    .C1(\u_cpu.ALU.u_wallace._3597_ ),
    .Y(\u_cpu.ALU.u_wallace._3598_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9125_  (.A1(\u_cpu.ALU.u_wallace._3595_ ),
    .A2(\u_cpu.ALU.u_wallace._3593_ ),
    .B1(\u_cpu.ALU.u_wallace._3596_ ),
    .Y(\u_cpu.ALU.u_wallace._3599_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9126_  (.A1(\u_cpu.ALU.u_wallace._3587_ ),
    .A2(\u_cpu.ALU.u_wallace._3588_ ),
    .B1(\u_cpu.ALU.u_wallace._3595_ ),
    .C1(\u_cpu.ALU.u_wallace._3593_ ),
    .X(\u_cpu.ALU.u_wallace._3600_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._9127_  (.A1(\u_cpu.ALU.u_wallace._3308_ ),
    .A2(\u_cpu.ALU.u_wallace._3304_ ),
    .B1(\u_cpu.ALU.u_wallace._3312_ ),
    .X(\u_cpu.ALU.u_wallace._3601_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9128_  (.A1(\u_cpu.ALU.u_wallace._3599_ ),
    .A2(\u_cpu.ALU.u_wallace._3600_ ),
    .B1(\u_cpu.ALU.u_wallace._3601_ ),
    .Y(\u_cpu.ALU.u_wallace._3603_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9129_  (.A(\u_cpu.ALU.u_wallace._3598_ ),
    .B(\u_cpu.ALU.u_wallace._3603_ ),
    .Y(\u_cpu.ALU.u_wallace._3604_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._9130_  (.A1(\u_cpu.ALU.u_wallace._3586_ ),
    .A2(\u_cpu.ALU.u_wallace._3594_ ),
    .B1(\u_cpu.ALU.u_wallace._3307_ ),
    .B2(\u_cpu.ALU.u_wallace._3318_ ),
    .C1(\u_cpu.ALU.u_wallace._3597_ ),
    .X(\u_cpu.ALU.u_wallace._3605_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9131_  (.A(\u_cpu.ALU.u_wallace._3337_ ),
    .B(\u_cpu.ALU.u_wallace._3603_ ),
    .Y(\u_cpu.ALU.u_wallace._3606_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._9132_  (.A1_N(\u_cpu.ALU.u_wallace._3339_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3604_ ),
    .B1(\u_cpu.ALU.u_wallace._3605_ ),
    .B2(\u_cpu.ALU.u_wallace._3606_ ),
    .Y(\u_cpu.ALU.u_wallace._3607_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._9133_  (.A(\u_cpu.ALU.u_wallace._3335_ ),
    .B(\u_cpu.ALU.u_wallace._3607_ ),
    .X(\u_cpu.ALU.u_wallace._3608_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9134_  (.A(\u_cpu.ALU.u_wallace._3037_ ),
    .B(\u_cpu.ALU.u_wallace._3040_ ),
    .C(\u_cpu.ALU.u_wallace._3332_ ),
    .D(\u_cpu.ALU.u_wallace._2468_ ),
    .Y(\u_cpu.ALU.u_wallace._3609_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9135_  (.A1(\u_cpu.ALU.u_wallace._3320_ ),
    .A2(\u_cpu.ALU.u_wallace._3330_ ),
    .B1(\u_cpu.ALU.u_wallace._3323_ ),
    .C1(\u_cpu.ALU.u_wallace._3327_ ),
    .Y(\u_cpu.ALU.u_wallace._3610_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9136_  (.A(\u_cpu.ALU.u_wallace._3031_ ),
    .B(\u_cpu.ALU.u_wallace._3039_ ),
    .C(\u_cpu.ALU.u_wallace._3036_ ),
    .D(\u_cpu.ALU.u_wallace._2751_ ),
    .Y(\u_cpu.ALU.u_wallace._3611_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._9137_  (.A1(\u_cpu.ALU.u_wallace._3036_ ),
    .A2(\u_cpu.ALU.u_wallace._3610_ ),
    .A3(\u_cpu.ALU.u_wallace._3611_ ),
    .B1(\u_cpu.ALU.u_wallace._3329_ ),
    .X(\u_cpu.ALU.u_wallace._3612_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9138_  (.A(\u_cpu.ALU.u_wallace._3609_ ),
    .B(\u_cpu.ALU.u_wallace._3612_ ),
    .Y(\u_cpu.ALU.u_wallace._3614_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._9139_  (.A(\u_cpu.ALU.u_wallace._3608_ ),
    .B(\u_cpu.ALU.u_wallace._3614_ ),
    .X(\u_cpu.ALU.Product_Wallace[28] ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9140_  (.A(\u_cpu.ALU.u_wallace._3614_ ),
    .B(\u_cpu.ALU.u_wallace._3608_ ),
    .Y(\u_cpu.ALU.u_wallace._3615_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9141_  (.A1(\u_cpu.ALU.u_wallace._3384_ ),
    .A2(\u_cpu.ALU.u_wallace._3387_ ),
    .B1(\u_cpu.ALU.u_wallace._3391_ ),
    .C1(\u_cpu.ALU.u_wallace._3510_ ),
    .Y(\u_cpu.ALU.u_wallace._3616_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9142_  (.A(\u_cpu.ALU.u_wallace._3505_ ),
    .B(\u_cpu.ALU.u_wallace._3616_ ),
    .Y(\u_cpu.ALU.u_wallace._3617_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9143_  (.A(\u_cpu.ALU.u_wallace._4798_ ),
    .B(\u_cpu.ALU.u_wallace._0958_ ),
    .Y(\u_cpu.ALU.u_wallace._3618_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9144_  (.A(\u_cpu.ALU.u_wallace._3618_ ),
    .B(\u_cpu.ALU.u_wallace._1176_ ),
    .C(\u_cpu.ALU.u_wallace._0847_ ),
    .Y(\u_cpu.ALU.u_wallace._3619_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9145_  (.A(\u_cpu.ALU.u_wallace._0847_ ),
    .B(\u_cpu.ALU.u_wallace._1208_ ),
    .Y(\u_cpu.ALU.u_wallace._3620_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9146_  (.A(\u_cpu.ALU.u_wallace._3620_ ),
    .B(\u_cpu.ALU.u_wallace._0958_ ),
    .C(\u_cpu.ALU.u_wallace._1129_ ),
    .Y(\u_cpu.ALU.u_wallace._3621_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9147_  (.A1(\u_cpu.ALU.u_wallace._4573_ ),
    .A2(\u_cpu.ALU.u_wallace._2053_ ),
    .B1(\u_cpu.ALU.u_wallace._3619_ ),
    .C1(\u_cpu.ALU.u_wallace._3621_ ),
    .Y(\u_cpu.ALU.u_wallace._3622_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9148_  (.A1(\u_cpu.ALU.u_wallace._4798_ ),
    .A2(\u_cpu.ALU.u_wallace._0958_ ),
    .B1(\u_cpu.ALU.u_wallace._1176_ ),
    .B2(\u_cpu.ALU.u_wallace._4643_ ),
    .X(\u_cpu.ALU.u_wallace._3624_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9149_  (.A(\u_cpu.ALU.u_wallace._0847_ ),
    .B(\u_cpu.ALU.u_wallace._1129_ ),
    .C(\u_cpu.ALU.u_wallace._0958_ ),
    .D(\u_cpu.ALU.u_wallace._1176_ ),
    .Y(\u_cpu.ALU.u_wallace._3625_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9150_  (.A(\u_cpu.ALU.u_wallace._3624_ ),
    .B(\u_cpu.ALU.u_wallace._1615_ ),
    .C(\u_cpu.ALU.u_wallace._0607_ ),
    .D(\u_cpu.ALU.u_wallace._3625_ ),
    .Y(\u_cpu.ALU.u_wallace._3626_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9151_  (.A(\u_cpu.ALU.u_wallace._4661_ ),
    .B(\u_cpu.ALU.u_wallace._1615_ ),
    .Y(\u_cpu.ALU.u_wallace._3627_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9152_  (.A1(\u_cpu.ALU.u_wallace._3627_ ),
    .A2(\u_cpu.ALU.u_wallace._3364_ ),
    .B1(\u_cpu.ALU.u_wallace._3365_ ),
    .Y(\u_cpu.ALU.u_wallace._3628_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9153_  (.A1(\u_cpu.ALU.u_wallace._3622_ ),
    .A2(\u_cpu.ALU.u_wallace._3626_ ),
    .B1(\u_cpu.ALU.u_wallace._3628_ ),
    .Y(\u_cpu.ALU.u_wallace._3629_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9154_  (.A(\u_cpu.ALU.u_wallace._3628_ ),
    .B(\u_cpu.ALU.u_wallace._3622_ ),
    .C(\u_cpu.ALU.u_wallace._3626_ ),
    .X(\u_cpu.ALU.u_wallace._3630_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9155_  (.A(\u_cpu.ALU.u_wallace._4661_ ),
    .B(\u_cpu.ALU.u_wallace._2343_ ),
    .C(\u_cpu.ALU.u_wallace._1610_ ),
    .D(\u_cpu.ALU.u_wallace._1824_ ),
    .X(\u_cpu.ALU.u_wallace._3631_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9156_  (.A1(\u_cpu.ALU.u_wallace._4661_ ),
    .A2(\u_cpu.ALU.u_wallace._1611_ ),
    .B1(\u_cpu.ALU.u_wallace._1855_ ),
    .B2(\u_cpu.ALU.u_wallace._2343_ ),
    .Y(\u_cpu.ALU.u_wallace._3632_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9157_  (.A(\u_cpu.ALU.u_wallace._3631_ ),
    .B(\u_cpu.ALU.u_wallace._3632_ ),
    .Y(\u_cpu.ALU.u_wallace._3633_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._9158_  (.A1(\u_cpu.ALU.u_wallace._3629_ ),
    .A2(\u_cpu.ALU.u_wallace._3630_ ),
    .B1(\u_cpu.ALU.u_wallace._3633_ ),
    .X(\u_cpu.ALU.u_wallace._3635_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._9159_  (.A(\u_cpu.ALU.u_wallace._3629_ ),
    .B(\u_cpu.ALU.u_wallace._3630_ ),
    .C(\u_cpu.ALU.u_wallace._3633_ ),
    .Y(\u_cpu.ALU.u_wallace._3636_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9160_  (.A(\u_cpu.ALU.u_wallace._4894_ ),
    .B(\u_cpu.ALU.u_wallace._1075_ ),
    .Y(\u_cpu.ALU.u_wallace._3637_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9161_  (.A(\u_cpu.ALU.u_wallace._4732_ ),
    .B(\u_cpu.ALU.u_wallace._1286_ ),
    .Y(\u_cpu.ALU.u_wallace._3638_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9162_  (.A(\u_cpu.ALU.u_wallace._0034_ ),
    .B(\u_cpu.ALU.u_wallace._1974_ ),
    .Y(\u_cpu.ALU.u_wallace._3639_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9163_  (.A1(\u_cpu.ALU.u_wallace._3637_ ),
    .A2(\u_cpu.ALU.u_wallace._3638_ ),
    .B1(\u_cpu.ALU.u_wallace._3639_ ),
    .Y(\u_cpu.ALU.u_wallace._3640_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9164_  (.A1(\u_cpu.ALU.u_wallace._0121_ ),
    .A2(\u_cpu.ALU.u_wallace._0826_ ),
    .B1(\u_cpu.ALU.u_wallace._0279_ ),
    .B2(\u_cpu.ALU.u_wallace._0320_ ),
    .X(\u_cpu.ALU.u_wallace._3641_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9165_  (.A(\u_cpu.ALU.u_wallace._0652_ ),
    .B(\u_cpu.ALU.u_wallace._0121_ ),
    .C(\u_cpu.ALU.u_wallace._0826_ ),
    .D(\u_cpu.ALU.u_wallace._0279_ ),
    .Y(\u_cpu.ALU.u_wallace._3642_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9166_  (.A(\u_cpu.ALU.u_wallace._3641_ ),
    .B(\u_cpu.ALU.u_wallace._3642_ ),
    .C(\u_cpu.ALU.u_wallace._1578_ ),
    .D(\u_cpu.ALU.u_wallace._0551_ ),
    .Y(\u_cpu.ALU.u_wallace._3643_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9167_  (.A1(\u_cpu.ALU.u_wallace._0121_ ),
    .A2(\u_cpu.ALU.u_wallace._0826_ ),
    .B1(\u_cpu.ALU.u_wallace._0280_ ),
    .B2(\u_cpu.ALU.u_wallace._0652_ ),
    .Y(\u_cpu.ALU.u_wallace._3644_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9168_  (.A(\u_cpu.ALU.u_wallace._0320_ ),
    .B(\u_cpu.ALU.u_wallace._0121_ ),
    .C(\u_cpu.ALU.u_wallace._0826_ ),
    .D(\u_cpu.ALU.u_wallace._0279_ ),
    .X(\u_cpu.ALU.u_wallace._3646_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9169_  (.A1(\u_cpu.ALU.u_wallace._0458_ ),
    .A2(\u_cpu.ALU.u_wallace._0554_ ),
    .B1(\u_cpu.ALU.u_wallace._3644_ ),
    .B2(\u_cpu.ALU.u_wallace._3646_ ),
    .Y(\u_cpu.ALU.u_wallace._3647_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9170_  (.A1(\u_cpu.ALU.u_wallace._3472_ ),
    .A2(\u_cpu.ALU.u_wallace._3640_ ),
    .B1(\u_cpu.ALU.u_wallace._3643_ ),
    .C1(\u_cpu.ALU.u_wallace._3647_ ),
    .X(\u_cpu.ALU.u_wallace._3648_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9171_  (.A(\u_cpu.ALU.u_wallace._3472_ ),
    .B(\u_cpu.ALU.u_wallace._3640_ ),
    .Y(\u_cpu.ALU.u_wallace._3649_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9172_  (.A(\u_cpu.ALU.u_wallace._3643_ ),
    .B(\u_cpu.ALU.u_wallace._3647_ ),
    .Y(\u_cpu.ALU.u_wallace._3650_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9173_  (.A(\u_cpu.ALU.u_wallace._1578_ ),
    .B(\u_cpu.ALU.u_wallace._0652_ ),
    .C(\u_cpu.ALU.u_wallace._0121_ ),
    .D(\u_cpu.ALU.u_wallace._0280_ ),
    .X(\u_cpu.ALU.u_wallace._3651_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9174_  (.A(\u_cpu.ALU.u_wallace._3344_ ),
    .B(\u_cpu.ALU.u_wallace._3204_ ),
    .C(\u_cpu.ALU.u_wallace._2658_ ),
    .X(\u_cpu.ALU.u_wallace._3652_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._9175_  (.A1_N(\u_cpu.ALU.u_wallace._3649_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3650_ ),
    .B1(\u_cpu.ALU.u_wallace._3651_ ),
    .B2(\u_cpu.ALU.u_wallace._3652_ ),
    .Y(\u_cpu.ALU.u_wallace._3653_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._9176_  (.A1(\u_cpu.ALU.u_wallace._3639_ ),
    .A2(\u_cpu.ALU.u_wallace._3471_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3472_ ),
    .Y(\u_cpu.ALU.u_wallace._3654_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9177_  (.A1(\u_cpu.ALU.u_wallace._3643_ ),
    .A2(\u_cpu.ALU.u_wallace._3647_ ),
    .B1(\u_cpu.ALU.u_wallace._3654_ ),
    .Y(\u_cpu.ALU.u_wallace._3655_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._9178_  (.A1(\u_cpu.ALU.u_wallace._3344_ ),
    .A2(\u_cpu.ALU.u_wallace._3204_ ),
    .A3(\u_cpu.ALU.u_wallace._2658_ ),
    .B1(\u_cpu.ALU.u_wallace._3651_ ),
    .Y(\u_cpu.ALU.u_wallace._3657_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9179_  (.A1(\u_cpu.ALU.u_wallace._3648_ ),
    .A2(\u_cpu.ALU.u_wallace._3655_ ),
    .B1(\u_cpu.ALU.u_wallace._3657_ ),
    .Y(\u_cpu.ALU.u_wallace._3658_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._9180_  (.A1_N(\u_cpu.ALU.u_wallace._3351_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3355_ ),
    .B1(\u_cpu.ALU.u_wallace._3353_ ),
    .B2(\u_cpu.ALU.u_wallace._3354_ ),
    .Y(\u_cpu.ALU.u_wallace._3659_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9181_  (.A1(\u_cpu.ALU.u_wallace._3648_ ),
    .A2(\u_cpu.ALU.u_wallace._3653_ ),
    .B1(\u_cpu.ALU.u_wallace._3658_ ),
    .C1(\u_cpu.ALU.u_wallace._3659_ ),
    .X(\u_cpu.ALU.u_wallace._3660_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9182_  (.A1(\u_cpu.ALU.u_wallace._3650_ ),
    .A2(\u_cpu.ALU.u_wallace._3649_ ),
    .B1(\u_cpu.ALU.u_wallace._3657_ ),
    .Y(\u_cpu.ALU.u_wallace._3661_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9183_  (.A1(\u_cpu.ALU.u_wallace._3649_ ),
    .A2(\u_cpu.ALU.u_wallace._3650_ ),
    .B1(\u_cpu.ALU.u_wallace._3661_ ),
    .Y(\u_cpu.ALU.u_wallace._3662_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9184_  (.A1(\u_cpu.ALU.u_wallace._3662_ ),
    .A2(\u_cpu.ALU.u_wallace._3658_ ),
    .B1(\u_cpu.ALU.u_wallace._3659_ ),
    .Y(\u_cpu.ALU.u_wallace._3663_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9185_  (.A1(\u_cpu.ALU.u_wallace._3635_ ),
    .A2(\u_cpu.ALU.u_wallace._3636_ ),
    .B1(\u_cpu.ALU.u_wallace._3660_ ),
    .B2(\u_cpu.ALU.u_wallace._3663_ ),
    .Y(\u_cpu.ALU.u_wallace._3664_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9186_  (.A1(\u_cpu.ALU.u_wallace._3662_ ),
    .A2(\u_cpu.ALU.u_wallace._3658_ ),
    .B1(\u_cpu.ALU.u_wallace._3659_ ),
    .X(\u_cpu.ALU.u_wallace._3665_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9187_  (.A(\u_cpu.ALU.u_wallace._3635_ ),
    .B(\u_cpu.ALU.u_wallace._3636_ ),
    .Y(\u_cpu.ALU.u_wallace._3666_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9188_  (.A1(\u_cpu.ALU.u_wallace._3648_ ),
    .A2(\u_cpu.ALU.u_wallace._3653_ ),
    .B1(\u_cpu.ALU.u_wallace._3658_ ),
    .C1(\u_cpu.ALU.u_wallace._3659_ ),
    .Y(\u_cpu.ALU.u_wallace._3668_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9189_  (.A(\u_cpu.ALU.u_wallace._3665_ ),
    .B(\u_cpu.ALU.u_wallace._3666_ ),
    .C(\u_cpu.ALU.u_wallace._3668_ ),
    .Y(\u_cpu.ALU.u_wallace._3669_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9190_  (.A(\u_cpu.ALU.u_wallace._3487_ ),
    .B(\u_cpu.ALU.u_wallace._3501_ ),
    .C(\u_cpu.ALU.u_wallace._3664_ ),
    .D(\u_cpu.ALU.u_wallace._3669_ ),
    .Y(\u_cpu.ALU.u_wallace._3670_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9191_  (.A1(\u_cpu.ALU.u_wallace._3483_ ),
    .A2(\u_cpu.ALU.u_wallace._3484_ ),
    .B1(\u_cpu.ALU.u_wallace._3482_ ),
    .Y(\u_cpu.ALU.u_wallace._3671_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9192_  (.A1(\u_cpu.ALU.u_wallace._3485_ ),
    .A2(\u_cpu.ALU.u_wallace._3671_ ),
    .B1(\u_cpu.ALU.u_wallace._3487_ ),
    .Y(\u_cpu.ALU.u_wallace._3672_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9193_  (.A1(\u_cpu.ALU.u_wallace._3635_ ),
    .A2(\u_cpu.ALU.u_wallace._3636_ ),
    .B1(\u_cpu.ALU.u_wallace._3668_ ),
    .C1(\u_cpu.ALU.u_wallace._3665_ ),
    .Y(\u_cpu.ALU.u_wallace._3673_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9194_  (.A1(\u_cpu.ALU.u_wallace._3660_ ),
    .A2(\u_cpu.ALU.u_wallace._3663_ ),
    .B1(\u_cpu.ALU.u_wallace._3666_ ),
    .Y(\u_cpu.ALU.u_wallace._3674_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9195_  (.A(\u_cpu.ALU.u_wallace._3672_ ),
    .B(\u_cpu.ALU.u_wallace._3673_ ),
    .C(\u_cpu.ALU.u_wallace._3674_ ),
    .Y(\u_cpu.ALU.u_wallace._3675_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._9196_  (.A1(\u_cpu.ALU.u_wallace._3358_ ),
    .A2(\u_cpu.ALU.u_wallace._3352_ ),
    .A3(\u_cpu.ALU.u_wallace._3356_ ),
    .B1(\u_cpu.ALU.u_wallace._3376_ ),
    .B2(\u_cpu.ALU.u_wallace._3379_ ),
    .X(\u_cpu.ALU.u_wallace._3676_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9197_  (.A1(\u_cpu.ALU.u_wallace._3670_ ),
    .A2(\u_cpu.ALU.u_wallace._3675_ ),
    .B1(\u_cpu.ALU.u_wallace._3676_ ),
    .X(\u_cpu.ALU.u_wallace._3677_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9198_  (.A(\u_cpu.ALU.u_wallace._3676_ ),
    .B(\u_cpu.ALU.u_wallace._3670_ ),
    .C(\u_cpu.ALU.u_wallace._3675_ ),
    .Y(\u_cpu.ALU.u_wallace._3679_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9199_  (.A1(\u_cpu.ALU.u_wallace._3490_ ),
    .A2(\u_cpu.ALU.u_wallace._3497_ ),
    .B1(\u_cpu.ALU.u_wallace._3458_ ),
    .X(\u_cpu.ALU.u_wallace._3680_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._9200_  (.A1(\u_cpu.ALU.u_wallace._3468_ ),
    .A2(\u_cpu.ALU.u_wallace._3465_ ),
    .A3(\u_cpu.ALU.u_wallace._3466_ ),
    .B1(\u_cpu.ALU.u_wallace._3478_ ),
    .B2(\u_cpu.ALU.u_wallace._3475_ ),
    .X(\u_cpu.ALU.u_wallace._3681_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9201_  (.A(\u_cpu.ALU.u_wallace._4605_ ),
    .B(\u_cpu.ALU.u_wallace._2916_ ),
    .Y(\u_cpu.ALU.u_wallace._3682_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9202_  (.A1(\u_cpu.ALU.u_wallace._4313_ ),
    .A2(\u_cpu.ALU.u_wallace._2907_ ),
    .B1(\u_cpu.ALU.u_wallace._3088_ ),
    .B2(\u_cpu.ALU.u_wallace._4029_ ),
    .Y(\u_cpu.ALU.u_wallace._3683_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9203_  (.A1(\u_cpu.ALU.u_wallace._3682_ ),
    .A2(\u_cpu.ALU.u_wallace._3683_ ),
    .B1(\u_cpu.ALU.u_wallace._3464_ ),
    .Y(\u_cpu.ALU.u_wallace._3684_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9204_  (.A(\u_cpu.ALU.u_wallace._4717_ ),
    .B(\u_cpu.ALU.u_wallace._4599_ ),
    .C(\u_cpu.ALU.u_wallace._1531_ ),
    .Y(\u_cpu.ALU.u_wallace._3685_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9205_  (.A1(\u_cpu.ALU.u_wallace._4599_ ),
    .A2(\u_cpu.ALU.u_wallace._1275_ ),
    .B1(\u_cpu.ALU.u_wallace._1531_ ),
    .B2(\u_cpu.ALU.u_wallace._4717_ ),
    .X(\u_cpu.ALU.u_wallace._3686_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._9206_  (.A1(\u_cpu.ALU.u_wallace._1271_ ),
    .A2(\u_cpu.ALU.u_wallace._3685_ ),
    .B1(\u_cpu.ALU.u_wallace._4605_ ),
    .C1(\u_cpu.ALU.u_wallace._2907_ ),
    .D1(\u_cpu.ALU.u_wallace._3686_ ),
    .Y(\u_cpu.ALU.u_wallace._3687_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9207_  (.A(\u_cpu.ALU.u_wallace._4029_ ),
    .B(\u_cpu.ALU.u_wallace._4313_ ),
    .C(\u_cpu.ALU.u_wallace._3088_ ),
    .D(\u_cpu.ALU.u_wallace._2618_ ),
    .Y(\u_cpu.ALU.u_wallace._3688_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9208_  (.A1(\u_cpu.ALU.u_wallace._4605_ ),
    .A2(\u_cpu.ALU.u_wallace._2907_ ),
    .B1(\u_cpu.ALU.u_wallace._3686_ ),
    .B2(\u_cpu.ALU.u_wallace._3688_ ),
    .X(\u_cpu.ALU.u_wallace._3690_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9209_  (.A(\u_cpu.ALU.u_wallace._3684_ ),
    .B(\u_cpu.ALU.u_wallace._3687_ ),
    .C(\u_cpu.ALU.u_wallace._3690_ ),
    .Y(\u_cpu.ALU.u_wallace._3691_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._9210_  (.A(\u_cpu.ALU.u_wallace._4604_ ),
    .B(\u_cpu.ALU.u_wallace._1101_ ),
    .X(\u_cpu.ALU.u_wallace._3692_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9211_  (.A1(\u_cpu.ALU.u_wallace._1271_ ),
    .A2(\u_cpu.ALU.u_wallace._3685_ ),
    .B1(\u_cpu.ALU.u_wallace._3692_ ),
    .C1(\u_cpu.ALU.u_wallace._3686_ ),
    .X(\u_cpu.ALU.u_wallace._3693_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9212_  (.A1(\u_cpu.ALU.u_wallace._3686_ ),
    .A2(\u_cpu.ALU.u_wallace._3688_ ),
    .B1(\u_cpu.ALU.u_wallace._3692_ ),
    .Y(\u_cpu.ALU.u_wallace._3694_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._9213_  (.A1(\u_cpu.ALU.u_wallace._3693_ ),
    .A2(\u_cpu.ALU.u_wallace._3694_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3684_ ),
    .Y(\u_cpu.ALU.u_wallace._3695_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9214_  (.A1(\u_cpu.ALU.u_wallace._4894_ ),
    .A2(\u_cpu.ALU.u_wallace._1286_ ),
    .B1(\u_cpu.ALU.u_wallace._2916_ ),
    .B2(\u_cpu.ALU.u_wallace._4732_ ),
    .X(\u_cpu.ALU.u_wallace._3696_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9215_  (.A(\u_cpu.ALU.u_wallace._4732_ ),
    .B(\u_cpu.ALU.u_wallace._4894_ ),
    .C(\u_cpu.ALU.u_wallace._2621_ ),
    .D(\u_cpu.ALU.u_wallace._2916_ ),
    .Y(\u_cpu.ALU.u_wallace._3697_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._9216_  (.A(\u_cpu.ALU.u_wallace._0034_ ),
    .B(\u_cpu.ALU.u_wallace._2248_ ),
    .X(\u_cpu.ALU.u_wallace._3698_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9217_  (.A(\u_cpu.ALU.u_wallace._3696_ ),
    .B(\u_cpu.ALU.u_wallace._3697_ ),
    .C(\u_cpu.ALU.u_wallace._3698_ ),
    .X(\u_cpu.ALU.u_wallace._3699_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9218_  (.A1(\u_cpu.ALU.u_wallace._4894_ ),
    .A2(\u_cpu.ALU.u_wallace._2621_ ),
    .B1(\u_cpu.ALU.u_wallace._2916_ ),
    .B2(\u_cpu.ALU.u_wallace._4732_ ),
    .Y(\u_cpu.ALU.u_wallace._3701_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9219_  (.A(\u_cpu.ALU.u_wallace._4732_ ),
    .B(\u_cpu.ALU.u_wallace._4894_ ),
    .C(\u_cpu.ALU.u_wallace._1286_ ),
    .D(\u_cpu.ALU.u_wallace._0815_ ),
    .X(\u_cpu.ALU.u_wallace._3702_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._9220_  (.A1(\u_cpu.ALU.u_wallace._0124_ ),
    .A2(\u_cpu.ALU.u_wallace._0442_ ),
    .B1(\u_cpu.ALU.u_wallace._3701_ ),
    .B2(\u_cpu.ALU.u_wallace._3702_ ),
    .X(\u_cpu.ALU.u_wallace._3703_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._9221_  (.A1_N(\u_cpu.ALU.u_wallace._3691_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3695_ ),
    .B1(\u_cpu.ALU.u_wallace._3699_ ),
    .B2(\u_cpu.ALU.u_wallace._3703_ ),
    .Y(\u_cpu.ALU.u_wallace._3704_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9222_  (.A(\u_cpu.ALU.u_wallace._0117_ ),
    .B(\u_cpu.ALU.u_wallace._2248_ ),
    .Y(\u_cpu.ALU.u_wallace._3705_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9223_  (.A(\u_cpu.ALU.u_wallace._3705_ ),
    .B(\u_cpu.ALU.u_wallace._3696_ ),
    .C(\u_cpu.ALU.u_wallace._3697_ ),
    .X(\u_cpu.ALU.u_wallace._3706_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9224_  (.A1(\u_cpu.ALU.u_wallace._3701_ ),
    .A2(\u_cpu.ALU.u_wallace._3702_ ),
    .B1(\u_cpu.ALU.u_wallace._0117_ ),
    .C1(\u_cpu.ALU.u_wallace._2248_ ),
    .X(\u_cpu.ALU.u_wallace._3707_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9225_  (.A1(\u_cpu.ALU.u_wallace._3706_ ),
    .A2(\u_cpu.ALU.u_wallace._3707_ ),
    .B1(\u_cpu.ALU.u_wallace._3691_ ),
    .C1(\u_cpu.ALU.u_wallace._3695_ ),
    .Y(\u_cpu.ALU.u_wallace._3708_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9226_  (.A(\u_cpu.ALU.u_wallace._3434_ ),
    .B(\u_cpu.ALU.u_wallace._3436_ ),
    .Y(\u_cpu.ALU.u_wallace._3709_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._9227_  (.A1_N(\u_cpu.ALU.u_wallace._3440_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3435_ ),
    .B1(\u_cpu.ALU.u_wallace._3709_ ),
    .B2(\u_cpu.ALU.u_wallace._3431_ ),
    .Y(\u_cpu.ALU.u_wallace._3710_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9228_  (.A1(\u_cpu.ALU.u_wallace._3704_ ),
    .A2(\u_cpu.ALU.u_wallace._3708_ ),
    .B1(\u_cpu.ALU.u_wallace._3710_ ),
    .X(\u_cpu.ALU.u_wallace._3712_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9229_  (.A(\u_cpu.ALU.u_wallace._3681_ ),
    .B(\u_cpu.ALU.u_wallace._3712_ ),
    .Y(\u_cpu.ALU.u_wallace._3713_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9230_  (.A(\u_cpu.ALU.u_wallace._3710_ ),
    .B(\u_cpu.ALU.u_wallace._3704_ ),
    .C(\u_cpu.ALU.u_wallace._3708_ ),
    .X(\u_cpu.ALU.u_wallace._3714_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9231_  (.A1(\u_cpu.ALU.u_wallace._3704_ ),
    .A2(\u_cpu.ALU.u_wallace._3708_ ),
    .B1(\u_cpu.ALU.u_wallace._3710_ ),
    .Y(\u_cpu.ALU.u_wallace._3715_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9232_  (.A1(\u_cpu.ALU.u_wallace._3475_ ),
    .A2(\u_cpu.ALU.u_wallace._3478_ ),
    .B1(\u_cpu.ALU.u_wallace._3467_ ),
    .Y(\u_cpu.ALU.u_wallace._3716_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9233_  (.A1(\u_cpu.ALU.u_wallace._3715_ ),
    .A2(\u_cpu.ALU.u_wallace._3714_ ),
    .B1(\u_cpu.ALU.u_wallace._3716_ ),
    .Y(\u_cpu.ALU.u_wallace._3717_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._9234_  (.A(\u_cpu.ALU.u_wallace._1102_ ),
    .X(\u_cpu.ALU.u_wallace._3718_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._9235_  (.A(\u_cpu.ALU.u_wallace._4431_ ),
    .X(\u_cpu.ALU.u_wallace._3719_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9236_  (.A1(\u_cpu.ALU.u_wallace._0475_ ),
    .A2(\u_cpu.ALU.u_wallace._3718_ ),
    .B1(\u_cpu.ALU.u_wallace._2882_ ),
    .B2(\u_cpu.ALU.u_wallace._3719_ ),
    .Y(\u_cpu.ALU.u_wallace._3720_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9237_  (.A(\u_cpu.ALU.u_wallace._0086_ ),
    .B(\u_cpu.ALU.SrcA[29] ),
    .Y(\u_cpu.ALU.u_wallace._3721_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9238_  (.A(\u_cpu.ALU.u_wallace._3719_ ),
    .B(\u_cpu.ALU.u_wallace._0475_ ),
    .C(\u_cpu.ALU.u_wallace._3718_ ),
    .D(\u_cpu.ALU.u_wallace._2002_ ),
    .X(\u_cpu.ALU.u_wallace._3723_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._9239_  (.A(\u_cpu.ALU.u_wallace._3720_ ),
    .B(\u_cpu.ALU.u_wallace._3721_ ),
    .C(\u_cpu.ALU.u_wallace._3723_ ),
    .Y(\u_cpu.ALU.u_wallace._3724_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9240_  (.A(\u_cpu.ALU.u_wallace._2779_ ),
    .B(\u_cpu.ALU.u_wallace._4917_ ),
    .C(\u_cpu.ALU.u_wallace._0629_ ),
    .D(\u_cpu.ALU.u_wallace._2002_ ),
    .Y(\u_cpu.ALU.u_wallace._3725_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9241_  (.A1(\u_cpu.ALU.u_wallace._4917_ ),
    .A2(\u_cpu.ALU.u_wallace._0629_ ),
    .B1(\u_cpu.ALU.u_wallace._2002_ ),
    .B2(\u_cpu.ALU.u_wallace._2779_ ),
    .X(\u_cpu.ALU.u_wallace._3726_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9242_  (.A1(\u_cpu.ALU.u_wallace._0884_ ),
    .A2(\u_cpu.ALU.SrcA[29] ),
    .B1(\u_cpu.ALU.u_wallace._3725_ ),
    .B2(\u_cpu.ALU.u_wallace._3726_ ),
    .Y(\u_cpu.ALU.u_wallace._3727_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9243_  (.A(\u_cpu.ALU.u_wallace._0086_ ),
    .B(\u_cpu.ALU.u_wallace._3399_ ),
    .Y(\u_cpu.ALU.u_wallace._3728_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9244_  (.A(\u_cpu.ALU.u_wallace._3719_ ),
    .B(\u_cpu.ALU.u_wallace._4798_ ),
    .C(\u_cpu.ALU.u_wallace._3718_ ),
    .D(\u_cpu.ALU.u_wallace._2598_ ),
    .Y(\u_cpu.ALU.u_wallace._3729_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9245_  (.A1(\u_cpu.ALU.u_wallace._3728_ ),
    .A2(\u_cpu.ALU.u_wallace._3401_ ),
    .B1(\u_cpu.ALU.u_wallace._3729_ ),
    .Y(\u_cpu.ALU.u_wallace._3730_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._9246_  (.A1(\u_cpu.ALU.u_wallace._3724_ ),
    .A2(\u_cpu.ALU.u_wallace._3727_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3730_ ),
    .Y(\u_cpu.ALU.u_wallace._3731_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9247_  (.A1(\u_cpu.ALU.u_wallace._0304_ ),
    .A2(\u_cpu.ALU.SrcA[27] ),
    .B1(\u_cpu.ALU.u_wallace._3399_ ),
    .B2(\u_cpu.ALU.u_wallace._1158_ ),
    .X(\u_cpu.ALU.u_wallace._3732_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9248_  (.A(\u_cpu.ALU.u_wallace._0217_ ),
    .B(\u_cpu.ALU.u_wallace._4796_ ),
    .C(\u_cpu.ALU.u_wallace._3058_ ),
    .D(\u_cpu.ALU.u_wallace._3399_ ),
    .Y(\u_cpu.ALU.u_wallace._3734_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9249_  (.A1(\u_cpu.ALU.u_wallace._4663_ ),
    .A2(\u_cpu.ALU.u_wallace._2869_ ),
    .B1(\u_cpu.ALU.u_wallace._3732_ ),
    .B2(\u_cpu.ALU.u_wallace._3734_ ),
    .Y(\u_cpu.ALU.u_wallace._3735_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9250_  (.A(\u_cpu.ALU.u_wallace._3732_ ),
    .B(\u_cpu.ALU.u_wallace._3734_ ),
    .C(\u_cpu.ALU.u_wallace._0983_ ),
    .D(\u_cpu.ALU.u_wallace._2869_ ),
    .X(\u_cpu.ALU.u_wallace._3736_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9251_  (.A(\u_cpu.ALU.u_wallace._3735_ ),
    .B(\u_cpu.ALU.u_wallace._3736_ ),
    .Y(\u_cpu.ALU.u_wallace._3737_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9252_  (.A(\u_cpu.ALU.u_wallace._4798_ ),
    .B(\u_cpu.ALU.u_wallace._3718_ ),
    .Y(\u_cpu.ALU.u_wallace._3738_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9253_  (.A(\u_cpu.ALU.u_wallace._3719_ ),
    .B(\u_cpu.ALU.u_wallace._1742_ ),
    .Y(\u_cpu.ALU.u_wallace._3739_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9254_  (.A1(\u_cpu.ALU.u_wallace._3738_ ),
    .A2(\u_cpu.ALU.u_wallace._3739_ ),
    .B1(\u_cpu.ALU.u_wallace._3728_ ),
    .Y(\u_cpu.ALU.u_wallace._3740_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9255_  (.A(\u_cpu.ALU.u_wallace._3726_ ),
    .B(\u_cpu.ALU.SrcA[29] ),
    .C(\u_cpu.ALU.u_wallace._0884_ ),
    .D(\u_cpu.ALU.u_wallace._3725_ ),
    .Y(\u_cpu.ALU.u_wallace._3741_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._9256_  (.A(\u_cpu.ALU.SrcA[29] ),
    .Y(\u_cpu.ALU.u_wallace._3742_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._9257_  (.A1_N(\u_cpu.ALU.u_wallace._3725_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3726_ ),
    .B1(\u_cpu.ALU.u_wallace._4934_ ),
    .B2(\u_cpu.ALU.u_wallace._3742_ ),
    .Y(\u_cpu.ALU.u_wallace._3743_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9258_  (.A1(\u_cpu.ALU.u_wallace._3402_ ),
    .A2(\u_cpu.ALU.u_wallace._3740_ ),
    .B1(\u_cpu.ALU.u_wallace._3741_ ),
    .C1(\u_cpu.ALU.u_wallace._3743_ ),
    .Y(\u_cpu.ALU.u_wallace._3745_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9259_  (.A(\u_cpu.ALU.u_wallace._3731_ ),
    .B(\u_cpu.ALU.u_wallace._3737_ ),
    .C(\u_cpu.ALU.u_wallace._3745_ ),
    .Y(\u_cpu.ALU.u_wallace._3746_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9260_  (.A1(\u_cpu.ALU.u_wallace._3402_ ),
    .A2(\u_cpu.ALU.u_wallace._3740_ ),
    .B1(\u_cpu.ALU.u_wallace._3741_ ),
    .C1(\u_cpu.ALU.u_wallace._3743_ ),
    .X(\u_cpu.ALU.u_wallace._3747_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9261_  (.A1(\u_cpu.ALU.u_wallace._3741_ ),
    .A2(\u_cpu.ALU.u_wallace._3743_ ),
    .B1(\u_cpu.ALU.u_wallace._3730_ ),
    .Y(\u_cpu.ALU.u_wallace._3748_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9262_  (.A1(\u_cpu.ALU.u_wallace._3735_ ),
    .A2(\u_cpu.ALU.u_wallace._3736_ ),
    .B1(\u_cpu.ALU.u_wallace._3747_ ),
    .B2(\u_cpu.ALU.u_wallace._3748_ ),
    .Y(\u_cpu.ALU.u_wallace._3749_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9263_  (.A1(\u_cpu.ALU.u_wallace._3417_ ),
    .A2(\u_cpu.ALU.u_wallace._3411_ ),
    .B1(\u_cpu.ALU.u_wallace._3746_ ),
    .C1(\u_cpu.ALU.u_wallace._3749_ ),
    .X(\u_cpu.ALU.u_wallace._3750_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9264_  (.A1(\u_cpu.ALU.u_wallace._3747_ ),
    .A2(\u_cpu.ALU.u_wallace._3748_ ),
    .B1(\u_cpu.ALU.u_wallace._3737_ ),
    .Y(\u_cpu.ALU.u_wallace._3751_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9265_  (.A1(\u_cpu.ALU.u_wallace._3735_ ),
    .A2(\u_cpu.ALU.u_wallace._3736_ ),
    .B1(\u_cpu.ALU.u_wallace._3745_ ),
    .C1(\u_cpu.ALU.u_wallace._3731_ ),
    .Y(\u_cpu.ALU.u_wallace._3752_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9266_  (.A1(\u_cpu.ALU.u_wallace._3413_ ),
    .A2(\u_cpu.ALU.u_wallace._3414_ ),
    .B1(\u_cpu.ALU.u_wallace._3079_ ),
    .X(\u_cpu.ALU.u_wallace._3753_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9267_  (.A1(\u_cpu.ALU.u_wallace._0097_ ),
    .A2(\u_cpu.ALU.u_wallace._3399_ ),
    .B1(\u_cpu.ALU.u_wallace._3397_ ),
    .B2(\u_cpu.ALU.u_wallace._3729_ ),
    .Y(\u_cpu.ALU.u_wallace._3754_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9268_  (.A1(\u_cpu.ALU.u_wallace._3057_ ),
    .A2(\u_cpu.ALU.u_wallace._3753_ ),
    .B1(\u_cpu.ALU.u_wallace._3754_ ),
    .Y(\u_cpu.ALU.u_wallace._3756_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9269_  (.A1(\u_cpu.ALU.u_wallace._1737_ ),
    .A2(\u_cpu.ALU.u_wallace._3395_ ),
    .B1(\u_cpu.ALU.u_wallace._3396_ ),
    .C1(\u_cpu.ALU.u_wallace._3397_ ),
    .X(\u_cpu.ALU.u_wallace._3757_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9270_  (.A1(\u_cpu.ALU.u_wallace._3757_ ),
    .A2(\u_cpu.ALU.u_wallace._3754_ ),
    .B1(\u_cpu.ALU.u_wallace._3394_ ),
    .Y(\u_cpu.ALU.u_wallace._3758_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9271_  (.A1(\u_cpu.ALU.u_wallace._3398_ ),
    .A2(\u_cpu.ALU.u_wallace._3756_ ),
    .B1(\u_cpu.ALU.u_wallace._3758_ ),
    .B2(\u_cpu.ALU.u_wallace._3420_ ),
    .Y(\u_cpu.ALU.u_wallace._3759_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9272_  (.A(\u_cpu.ALU.u_wallace._3751_ ),
    .B(\u_cpu.ALU.u_wallace._3752_ ),
    .C(\u_cpu.ALU.u_wallace._3759_ ),
    .Y(\u_cpu.ALU.u_wallace._3760_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9273_  (.A(\u_cpu.ALU.u_wallace._3408_ ),
    .B(\u_cpu.ALU.u_wallace._3447_ ),
    .Y(\u_cpu.ALU.u_wallace._3761_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9274_  (.A1(\u_cpu.ALU.u_wallace._1508_ ),
    .A2(\u_cpu.ALU.u_wallace._2569_ ),
    .B1(\u_cpu.ALU.u_wallace._3449_ ),
    .B2(\u_cpu.ALU.u_wallace._2166_ ),
    .Y(\u_cpu.ALU.u_wallace._3762_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9275_  (.A(\u_cpu.ALU.u_wallace._1476_ ),
    .B(\u_cpu.ALU.u_wallace._1508_ ),
    .C(\u_cpu.ALU.u_wallace._2222_ ),
    .D(\u_cpu.ALU.u_wallace._3449_ ),
    .X(\u_cpu.ALU.u_wallace._3763_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9276_  (.A1(\u_cpu.ALU.u_wallace._2284_ ),
    .A2(\u_cpu.ALU.u_wallace._1737_ ),
    .B1(\u_cpu.ALU.u_wallace._3762_ ),
    .B2(\u_cpu.ALU.u_wallace._3763_ ),
    .Y(\u_cpu.ALU.u_wallace._3764_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9277_  (.A1(\u_cpu.ALU.u_wallace._1508_ ),
    .A2(\u_cpu.ALU.u_wallace._2569_ ),
    .B1(\u_cpu.ALU.u_wallace._3449_ ),
    .B2(\u_cpu.ALU.u_wallace._1476_ ),
    .X(\u_cpu.ALU.u_wallace._3765_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9278_  (.A(\u_cpu.ALU.u_wallace._2166_ ),
    .B(\u_cpu.ALU.u_wallace._1508_ ),
    .C(\u_cpu.ALU.u_wallace._2569_ ),
    .D(\u_cpu.ALU.u_wallace._3449_ ),
    .Y(\u_cpu.ALU.u_wallace._3767_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9279_  (.A(\u_cpu.ALU.u_wallace._3765_ ),
    .B(\u_cpu.ALU.u_wallace._3767_ ),
    .C(\u_cpu.ALU.u_wallace._0015_ ),
    .D(\u_cpu.ALU.u_wallace._2598_ ),
    .Y(\u_cpu.ALU.u_wallace._3768_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9280_  (.A1(\u_cpu.ALU.u_wallace._3446_ ),
    .A2(\u_cpu.ALU.u_wallace._3761_ ),
    .B1(\u_cpu.ALU.u_wallace._3764_ ),
    .C1(\u_cpu.ALU.u_wallace._3768_ ),
    .Y(\u_cpu.ALU.u_wallace._3769_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._9281_  (.A1(\u_cpu.ALU.u_wallace._2284_ ),
    .A2(\u_cpu.ALU.u_wallace._1522_ ),
    .A3(\u_cpu.ALU.u_wallace._3428_ ),
    .B1(\u_cpu.ALU.u_wallace._3425_ ),
    .X(\u_cpu.ALU.u_wallace._3770_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9282_  (.A1(\u_cpu.ALU.u_wallace._3408_ ),
    .A2(\u_cpu.ALU.u_wallace._3447_ ),
    .B1(\u_cpu.ALU.u_wallace._3406_ ),
    .Y(\u_cpu.ALU.u_wallace._3771_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9283_  (.A1(\u_cpu.ALU.u_wallace._3764_ ),
    .A2(\u_cpu.ALU.u_wallace._3768_ ),
    .B1(\u_cpu.ALU.u_wallace._3771_ ),
    .Y(\u_cpu.ALU.u_wallace._3772_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9284_  (.A(\u_cpu.ALU.u_wallace._3770_ ),
    .B(\u_cpu.ALU.u_wallace._3772_ ),
    .Y(\u_cpu.ALU.u_wallace._3773_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9285_  (.A1(\u_cpu.ALU.u_wallace._2917_ ),
    .A2(\u_cpu.ALU.u_wallace._2598_ ),
    .B1(\u_cpu.ALU.u_wallace._3765_ ),
    .B2(\u_cpu.ALU.u_wallace._3767_ ),
    .Y(\u_cpu.ALU.u_wallace._3774_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9286_  (.A(\u_cpu.ALU.u_wallace._0015_ ),
    .B(\u_cpu.ALU.u_wallace._2598_ ),
    .Y(\u_cpu.ALU.u_wallace._3775_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._9287_  (.A(\u_cpu.ALU.u_wallace._3775_ ),
    .B(\u_cpu.ALU.u_wallace._3762_ ),
    .C(\u_cpu.ALU.u_wallace._3763_ ),
    .Y(\u_cpu.ALU.u_wallace._3776_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._9288_  (.A1(\u_cpu.ALU.u_wallace._3774_ ),
    .A2(\u_cpu.ALU.u_wallace._3776_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3771_ ),
    .Y(\u_cpu.ALU.u_wallace._3778_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._9289_  (.A1(\u_cpu.ALU.u_wallace._3424_ ),
    .A2(\u_cpu.ALU.u_wallace._2618_ ),
    .A3(\u_cpu.ALU.u_wallace._2917_ ),
    .B1(\u_cpu.ALU.u_wallace._3430_ ),
    .X(\u_cpu.ALU.u_wallace._3779_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9290_  (.A1(\u_cpu.ALU.u_wallace._3778_ ),
    .A2(\u_cpu.ALU.u_wallace._3769_ ),
    .B1(\u_cpu.ALU.u_wallace._3779_ ),
    .Y(\u_cpu.ALU.u_wallace._3780_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9291_  (.A1(\u_cpu.ALU.u_wallace._3769_ ),
    .A2(\u_cpu.ALU.u_wallace._3773_ ),
    .B1(\u_cpu.ALU.u_wallace._3780_ ),
    .Y(\u_cpu.ALU.u_wallace._3781_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9292_  (.A(\u_cpu.ALU.u_wallace._3760_ ),
    .B(\u_cpu.ALU.u_wallace._3781_ ),
    .Y(\u_cpu.ALU.u_wallace._3782_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9293_  (.A1(\u_cpu.ALU.u_wallace._3417_ ),
    .A2(\u_cpu.ALU.u_wallace._3452_ ),
    .B1(\u_cpu.ALU.u_wallace._3421_ ),
    .Y(\u_cpu.ALU.u_wallace._3783_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.ALU.u_wallace._9294_  (.A1(\u_cpu.ALU.u_wallace._3078_ ),
    .A2(\u_cpu.ALU.u_wallace._3080_ ),
    .A3(\u_cpu.ALU.u_wallace._3081_ ),
    .B1(\u_cpu.ALU.u_wallace._3072_ ),
    .B2(\u_cpu.ALU.u_wallace._3067_ ),
    .X(\u_cpu.ALU.u_wallace._3784_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9295_  (.A1(\u_cpu.ALU.u_wallace._3435_ ),
    .A2(\u_cpu.ALU.u_wallace._3439_ ),
    .B1(\u_cpu.ALU.u_wallace._3440_ ),
    .X(\u_cpu.ALU.u_wallace._3785_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9296_  (.A1(\u_cpu.ALU.u_wallace._3431_ ),
    .A2(\u_cpu.ALU.u_wallace._3709_ ),
    .B1(\u_cpu.ALU.u_wallace._3435_ ),
    .C1(\u_cpu.ALU.u_wallace._3440_ ),
    .Y(\u_cpu.ALU.u_wallace._3786_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9297_  (.A(\u_cpu.ALU.u_wallace._3785_ ),
    .B(\u_cpu.ALU.u_wallace._3786_ ),
    .Y(\u_cpu.ALU.u_wallace._3787_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9298_  (.A1(\u_cpu.ALU.u_wallace._3783_ ),
    .A2(\u_cpu.ALU.u_wallace._3784_ ),
    .B1(\u_cpu.ALU.u_wallace._3787_ ),
    .Y(\u_cpu.ALU.u_wallace._3789_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9299_  (.A(\u_cpu.ALU.u_wallace._3779_ ),
    .B(\u_cpu.ALU.u_wallace._3778_ ),
    .C(\u_cpu.ALU.u_wallace._3769_ ),
    .X(\u_cpu.ALU.u_wallace._3790_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._9300_  (.A1(\u_cpu.ALU.u_wallace._3746_ ),
    .A2(\u_cpu.ALU.u_wallace._3749_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3759_ ),
    .Y(\u_cpu.ALU.u_wallace._3791_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9301_  (.A1(\u_cpu.ALU.u_wallace._3780_ ),
    .A2(\u_cpu.ALU.u_wallace._3790_ ),
    .B1(\u_cpu.ALU.u_wallace._3750_ ),
    .B2(\u_cpu.ALU.u_wallace._3791_ ),
    .Y(\u_cpu.ALU.u_wallace._3792_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._9302_  (.A1(\u_cpu.ALU.u_wallace._3750_ ),
    .A2(\u_cpu.ALU.u_wallace._3782_ ),
    .B1(\u_cpu.ALU.u_wallace._3455_ ),
    .B2(\u_cpu.ALU.u_wallace._3789_ ),
    .C1(\u_cpu.ALU.u_wallace._3792_ ),
    .Y(\u_cpu.ALU.u_wallace._3793_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9303_  (.A1(\u_cpu.ALU.u_wallace._3417_ ),
    .A2(\u_cpu.ALU.u_wallace._3411_ ),
    .B1(\u_cpu.ALU.u_wallace._3749_ ),
    .Y(\u_cpu.ALU.u_wallace._3794_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._9304_  (.A(\u_cpu.ALU.u_wallace._3746_ ),
    .Y(\u_cpu.ALU.u_wallace._3795_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9305_  (.A1(\u_cpu.ALU.u_wallace._3794_ ),
    .A2(\u_cpu.ALU.u_wallace._3795_ ),
    .B1(\u_cpu.ALU.u_wallace._3781_ ),
    .C1(\u_cpu.ALU.u_wallace._3760_ ),
    .Y(\u_cpu.ALU.u_wallace._3796_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9306_  (.A1(\u_cpu.ALU.u_wallace._3787_ ),
    .A2(\u_cpu.ALU.u_wallace._3456_ ),
    .B1(\u_cpu.ALU.u_wallace._3453_ ),
    .Y(\u_cpu.ALU.u_wallace._3797_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9307_  (.A1(\u_cpu.ALU.u_wallace._3796_ ),
    .A2(\u_cpu.ALU.u_wallace._3792_ ),
    .B1(\u_cpu.ALU.u_wallace._3797_ ),
    .X(\u_cpu.ALU.u_wallace._3798_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._9308_  (.A1(\u_cpu.ALU.u_wallace._3713_ ),
    .A2(\u_cpu.ALU.u_wallace._3714_ ),
    .B1(\u_cpu.ALU.u_wallace._3717_ ),
    .C1(\u_cpu.ALU.u_wallace._3793_ ),
    .D1(\u_cpu.ALU.u_wallace._3798_ ),
    .Y(\u_cpu.ALU.u_wallace._3800_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9309_  (.A(\u_cpu.ALU.u_wallace._3710_ ),
    .B(\u_cpu.ALU.u_wallace._3704_ ),
    .C(\u_cpu.ALU.u_wallace._3708_ ),
    .Y(\u_cpu.ALU.u_wallace._3801_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9310_  (.A1(\u_cpu.ALU.u_wallace._3712_ ),
    .A2(\u_cpu.ALU.u_wallace._3801_ ),
    .B1(\u_cpu.ALU.u_wallace._3681_ ),
    .Y(\u_cpu.ALU.u_wallace._3802_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9311_  (.A(\u_cpu.ALU.u_wallace._3681_ ),
    .B(\u_cpu.ALU.u_wallace._3712_ ),
    .C(\u_cpu.ALU.u_wallace._3801_ ),
    .X(\u_cpu.ALU.u_wallace._3803_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._9312_  (.A1(\u_cpu.ALU.u_wallace._3750_ ),
    .A2(\u_cpu.ALU.u_wallace._3782_ ),
    .B1(\u_cpu.ALU.u_wallace._3455_ ),
    .B2(\u_cpu.ALU.u_wallace._3789_ ),
    .C1(\u_cpu.ALU.u_wallace._3792_ ),
    .X(\u_cpu.ALU.u_wallace._3804_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9313_  (.A1(\u_cpu.ALU.u_wallace._3796_ ),
    .A2(\u_cpu.ALU.u_wallace._3792_ ),
    .B1(\u_cpu.ALU.u_wallace._3797_ ),
    .Y(\u_cpu.ALU.u_wallace._3805_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9314_  (.A1(\u_cpu.ALU.u_wallace._3802_ ),
    .A2(\u_cpu.ALU.u_wallace._3803_ ),
    .B1(\u_cpu.ALU.u_wallace._3804_ ),
    .B2(\u_cpu.ALU.u_wallace._3805_ ),
    .Y(\u_cpu.ALU.u_wallace._3806_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9315_  (.A(\u_cpu.ALU.u_wallace._3680_ ),
    .B(\u_cpu.ALU.u_wallace._3800_ ),
    .C(\u_cpu.ALU.u_wallace._3806_ ),
    .Y(\u_cpu.ALU.u_wallace._3807_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9316_  (.A1(\u_cpu.ALU.u_wallace._3714_ ),
    .A2(\u_cpu.ALU.u_wallace._3713_ ),
    .B1(\u_cpu.ALU.u_wallace._3717_ ),
    .Y(\u_cpu.ALU.u_wallace._3808_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._9317_  (.A1(\u_cpu.ALU.u_wallace._3804_ ),
    .A2(\u_cpu.ALU.u_wallace._3805_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3808_ ),
    .Y(\u_cpu.ALU.u_wallace._3809_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9318_  (.A1(\u_cpu.ALU.u_wallace._3802_ ),
    .A2(\u_cpu.ALU.u_wallace._3803_ ),
    .B1(\u_cpu.ALU.u_wallace._3793_ ),
    .C1(\u_cpu.ALU.u_wallace._3798_ ),
    .Y(\u_cpu.ALU.u_wallace._3811_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9319_  (.A1(\u_cpu.ALU.u_wallace._3490_ ),
    .A2(\u_cpu.ALU.u_wallace._3497_ ),
    .B1(\u_cpu.ALU.u_wallace._3458_ ),
    .Y(\u_cpu.ALU.u_wallace._3812_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9320_  (.A(\u_cpu.ALU.u_wallace._3809_ ),
    .B(\u_cpu.ALU.u_wallace._3811_ ),
    .C(\u_cpu.ALU.u_wallace._3812_ ),
    .Y(\u_cpu.ALU.u_wallace._3813_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9321_  (.A(\u_cpu.ALU.u_wallace._3677_ ),
    .B(\u_cpu.ALU.u_wallace._3679_ ),
    .C(\u_cpu.ALU.u_wallace._3807_ ),
    .D(\u_cpu.ALU.u_wallace._3813_ ),
    .Y(\u_cpu.ALU.u_wallace._3814_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9322_  (.A1(\u_cpu.ALU.u_wallace._3677_ ),
    .A2(\u_cpu.ALU.u_wallace._3679_ ),
    .B1(\u_cpu.ALU.u_wallace._3807_ ),
    .B2(\u_cpu.ALU.u_wallace._3813_ ),
    .X(\u_cpu.ALU.u_wallace._3815_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9323_  (.A(\u_cpu.ALU.u_wallace._3617_ ),
    .B(\u_cpu.ALU.u_wallace._3814_ ),
    .C(\u_cpu.ALU.u_wallace._3815_ ),
    .Y(\u_cpu.ALU.u_wallace._3816_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9324_  (.A(\u_cpu.ALU.u_wallace._3677_ ),
    .B(\u_cpu.ALU.u_wallace._3679_ ),
    .Y(\u_cpu.ALU.u_wallace._3817_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9325_  (.A1(\u_cpu.ALU.u_wallace._3807_ ),
    .A2(\u_cpu.ALU.u_wallace._3813_ ),
    .B1(\u_cpu.ALU.u_wallace._3817_ ),
    .X(\u_cpu.ALU.u_wallace._3818_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9326_  (.A1(\u_cpu.ALU.u_wallace._3670_ ),
    .A2(\u_cpu.ALU.u_wallace._3675_ ),
    .B1(\u_cpu.ALU.u_wallace._3676_ ),
    .Y(\u_cpu.ALU.u_wallace._3819_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9327_  (.A(\u_cpu.ALU.u_wallace._3676_ ),
    .B(\u_cpu.ALU.u_wallace._3670_ ),
    .C(\u_cpu.ALU.u_wallace._3675_ ),
    .X(\u_cpu.ALU.u_wallace._3820_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9328_  (.A1(\u_cpu.ALU.u_wallace._3819_ ),
    .A2(\u_cpu.ALU.u_wallace._3820_ ),
    .B1(\u_cpu.ALU.u_wallace._3807_ ),
    .C1(\u_cpu.ALU.u_wallace._3813_ ),
    .Y(\u_cpu.ALU.u_wallace._3822_ ));
 sky130_fd_sc_hd__a32oi_2 \u_cpu.ALU.u_wallace._9329_  (.A1(\u_cpu.ALU.u_wallace._3377_ ),
    .A2(\u_cpu.ALU.u_wallace._3380_ ),
    .A3(\u_cpu.ALU.u_wallace._3383_ ),
    .B1(\u_cpu.ALU.u_wallace._3223_ ),
    .B2(\u_cpu.ALU.u_wallace._3220_ ),
    .Y(\u_cpu.ALU.u_wallace._3823_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9330_  (.A1(\u_cpu.ALU.u_wallace._3388_ ),
    .A2(\u_cpu.ALU.u_wallace._3389_ ),
    .B1(\u_cpu.ALU.u_wallace._3390_ ),
    .Y(\u_cpu.ALU.u_wallace._3824_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9331_  (.A1(\u_cpu.ALU.u_wallace._3389_ ),
    .A2(\u_cpu.ALU.u_wallace._3823_ ),
    .B1(\u_cpu.ALU.u_wallace._3824_ ),
    .Y(\u_cpu.ALU.u_wallace._3825_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._9332_  (.A1(\u_cpu.ALU.u_wallace._3825_ ),
    .A2(\u_cpu.ALU.u_wallace._3510_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3505_ ),
    .Y(\u_cpu.ALU.u_wallace._3826_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9333_  (.A(\u_cpu.ALU.u_wallace._3818_ ),
    .B(\u_cpu.ALU.u_wallace._3822_ ),
    .C(\u_cpu.ALU.u_wallace._3826_ ),
    .Y(\u_cpu.ALU.u_wallace._3827_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9334_  (.A1(\u_cpu.ALU.u_wallace._3381_ ),
    .A2(\u_cpu.ALU.u_wallace._3159_ ),
    .B1(\u_cpu.ALU.u_wallace._3386_ ),
    .Y(\u_cpu.ALU.u_wallace._3828_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9335_  (.A(\u_cpu.ALU.u_wallace._3376_ ),
    .B(\u_cpu.ALU.u_wallace._3378_ ),
    .C(\u_cpu.ALU.u_wallace._3379_ ),
    .X(\u_cpu.ALU.u_wallace._3829_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._9336_  (.A1_N(\u_cpu.ALU.u_wallace._3390_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3388_ ),
    .B1(\u_cpu.ALU.u_wallace._3828_ ),
    .B2(\u_cpu.ALU.u_wallace._3829_ ),
    .Y(\u_cpu.ALU.u_wallace._3830_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._9337_  (.A(\u_cpu.ALU.u_wallace._3534_ ),
    .Y(\u_cpu.ALU.u_wallace._3831_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9338_  (.A1(\u_cpu.ALU.u_wallace._3529_ ),
    .A2(\u_cpu.ALU.u_wallace._3522_ ),
    .B1(\u_cpu.ALU.u_wallace._3531_ ),
    .Y(\u_cpu.ALU.u_wallace._3833_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9339_  (.A1(\u_cpu.ALU.u_wallace._4527_ ),
    .A2(\u_cpu.ALU.SrcB[26] ),
    .B1(\u_cpu.ALU.SrcB[27] ),
    .B2(\u_cpu.ALU.u_wallace._0359_ ),
    .Y(\u_cpu.ALU.u_wallace._3834_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9340_  (.A(\u_cpu.ALU.u_wallace._4545_ ),
    .B(\u_cpu.ALU.u_wallace._4527_ ),
    .C(\u_cpu.ALU.u_wallace._3258_ ),
    .D(\u_cpu.ALU.u_wallace._3254_ ),
    .Y(\u_cpu.ALU.u_wallace._3835_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._9341_  (.A_N(\u_cpu.ALU.u_wallace._3834_ ),
    .B(\u_cpu.ALU.u_wallace._3835_ ),
    .C(\u_cpu.ALU.u_wallace._0917_ ),
    .D(\u_cpu.ALU.u_wallace._2480_ ),
    .Y(\u_cpu.ALU.u_wallace._3836_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9342_  (.A(\u_cpu.ALU.u_wallace._0359_ ),
    .B(\u_cpu.ALU.u_wallace._4527_ ),
    .C(\u_cpu.ALU.SrcB[26] ),
    .D(\u_cpu.ALU.SrcB[27] ),
    .X(\u_cpu.ALU.u_wallace._3837_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9343_  (.A1(\u_cpu.ALU.u_wallace._0939_ ),
    .A2(\u_cpu.ALU.u_wallace._2481_ ),
    .B1(\u_cpu.ALU.u_wallace._3834_ ),
    .B2(\u_cpu.ALU.u_wallace._3837_ ),
    .Y(\u_cpu.ALU.u_wallace._3838_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.ALU.u_wallace._9344_  (.A1(\u_cpu.ALU.u_wallace._0621_ ),
    .A2(\u_cpu.ALU.u_wallace._2481_ ),
    .A3(\u_cpu.ALU.u_wallace._3523_ ),
    .B1(\u_cpu.ALU.u_wallace._3527_ ),
    .Y(\u_cpu.ALU.u_wallace._3839_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9345_  (.A1(\u_cpu.ALU.u_wallace._3836_ ),
    .A2(\u_cpu.ALU.u_wallace._3838_ ),
    .B1(\u_cpu.ALU.u_wallace._3839_ ),
    .Y(\u_cpu.ALU.u_wallace._3840_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9346_  (.A(\u_cpu.ALU.u_wallace._3839_ ),
    .B(\u_cpu.ALU.u_wallace._3836_ ),
    .C(\u_cpu.ALU.u_wallace._3838_ ),
    .X(\u_cpu.ALU.u_wallace._3841_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._9347_  (.A1_N(\u_cpu.ALU.u_wallace._1333_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2402_ ),
    .B1(\u_cpu.ALU.u_wallace._3840_ ),
    .B2(\u_cpu.ALU.u_wallace._3841_ ),
    .Y(\u_cpu.ALU.u_wallace._3842_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9348_  (.A1(\u_cpu.ALU.u_wallace._3836_ ),
    .A2(\u_cpu.ALU.u_wallace._3838_ ),
    .B1(\u_cpu.ALU.u_wallace._3839_ ),
    .X(\u_cpu.ALU.u_wallace._3844_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9349_  (.A(\u_cpu.ALU.u_wallace._3839_ ),
    .B(\u_cpu.ALU.u_wallace._3836_ ),
    .C(\u_cpu.ALU.u_wallace._3838_ ),
    .Y(\u_cpu.ALU.u_wallace._3845_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9350_  (.A(\u_cpu.ALU.u_wallace._3844_ ),
    .B(\u_cpu.ALU.u_wallace._3845_ ),
    .C(\u_cpu.ALU.u_wallace._1333_ ),
    .D(\u_cpu.ALU.u_wallace._2402_ ),
    .Y(\u_cpu.ALU.u_wallace._3846_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9351_  (.A1(\u_cpu.ALU.u_wallace._3831_ ),
    .A2(\u_cpu.ALU.u_wallace._3833_ ),
    .B1(\u_cpu.ALU.u_wallace._3842_ ),
    .C1(\u_cpu.ALU.u_wallace._3846_ ),
    .X(\u_cpu.ALU.u_wallace._3847_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9352_  (.A1(\u_cpu.ALU.u_wallace._3531_ ),
    .A2(\u_cpu.ALU.u_wallace._3540_ ),
    .B1(\u_cpu.ALU.u_wallace._3534_ ),
    .Y(\u_cpu.ALU.u_wallace._3848_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9353_  (.A1(\u_cpu.ALU.u_wallace._3842_ ),
    .A2(\u_cpu.ALU.u_wallace._3846_ ),
    .B1(\u_cpu.ALU.u_wallace._3848_ ),
    .X(\u_cpu.ALU.u_wallace._3849_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9354_  (.A(\u_cpu.ALU.u_wallace._4454_ ),
    .B(\u_cpu.ALU.u_wallace._2131_ ),
    .Y(\u_cpu.ALU.u_wallace._3850_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._9355_  (.A_N(\u_cpu.ALU.u_wallace._3847_ ),
    .B(\u_cpu.ALU.u_wallace._3849_ ),
    .C(\u_cpu.ALU.u_wallace._3850_ ),
    .Y(\u_cpu.ALU.u_wallace._3851_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9356_  (.A1(\u_cpu.ALU.u_wallace._3842_ ),
    .A2(\u_cpu.ALU.u_wallace._3846_ ),
    .B1(\u_cpu.ALU.u_wallace._3848_ ),
    .Y(\u_cpu.ALU.u_wallace._3852_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9357_  (.A1(\u_cpu.ALU.u_wallace._4454_ ),
    .A2(\u_cpu.ALU.u_wallace._2131_ ),
    .B1(\u_cpu.ALU.u_wallace._3847_ ),
    .B2(\u_cpu.ALU.u_wallace._3852_ ),
    .Y(\u_cpu.ALU.u_wallace._3853_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9358_  (.A1(\u_cpu.ALU.u_wallace._0173_ ),
    .A2(\u_cpu.ALU.SrcB[28] ),
    .B1(\u_cpu.ALU.SrcB[29] ),
    .B2(\u_cpu.ALU.u_wallace._0118_ ),
    .Y(\u_cpu.ALU.u_wallace._3855_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9359_  (.A(\u_cpu.ALU.u_wallace._1070_ ),
    .B(\u_cpu.ALU.u_wallace._0272_ ),
    .C(\u_cpu.ALU.SrcB[28] ),
    .D(\u_cpu.ALU.SrcB[29] ),
    .X(\u_cpu.ALU.u_wallace._3856_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.ALU.u_wallace._9360_  (.A1(\u_cpu.ALU.u_wallace._3855_ ),
    .A2(\u_cpu.ALU.u_wallace._3856_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3362_ ),
    .X(\u_cpu.ALU.u_wallace._3857_ ));
 sky130_fd_sc_hd__nor3b_2 \u_cpu.ALU.u_wallace._9361_  (.A(\u_cpu.ALU.u_wallace._3855_ ),
    .B(\u_cpu.ALU.u_wallace._3856_ ),
    .C_N(\u_cpu.ALU.u_wallace._3362_ ),
    .Y(\u_cpu.ALU.u_wallace._3858_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9362_  (.A1(\u_cpu.ALU.u_wallace._3366_ ),
    .A2(\u_cpu.ALU.u_wallace._3368_ ),
    .B1(\u_cpu.ALU.u_wallace._3369_ ),
    .Y(\u_cpu.ALU.u_wallace._3859_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._9363_  (.A1(\u_cpu.ALU.u_wallace._3857_ ),
    .A2(\u_cpu.ALU.u_wallace._3858_ ),
    .B1(\u_cpu.ALU.u_wallace._3363_ ),
    .B2(\u_cpu.ALU.u_wallace._3859_ ),
    .C1(\u_cpu.ALU.u_wallace._3372_ ),
    .Y(\u_cpu.ALU.u_wallace._3860_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9364_  (.A1(\u_cpu.ALU.u_wallace._3363_ ),
    .A2(\u_cpu.ALU.u_wallace._3859_ ),
    .B1(\u_cpu.ALU.u_wallace._3372_ ),
    .Y(\u_cpu.ALU.u_wallace._3861_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9365_  (.A(\u_cpu.ALU.u_wallace._3857_ ),
    .B(\u_cpu.ALU.u_wallace._3858_ ),
    .Y(\u_cpu.ALU.u_wallace._3862_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9366_  (.A(\u_cpu.ALU.u_wallace._3861_ ),
    .B(\u_cpu.ALU.u_wallace._3862_ ),
    .Y(\u_cpu.ALU.u_wallace._3863_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9367_  (.A1(\u_cpu.ALU.u_wallace._3552_ ),
    .A2(\u_cpu.ALU.u_wallace._3554_ ),
    .B1(\u_cpu.ALU.u_wallace._3860_ ),
    .B2(\u_cpu.ALU.u_wallace._3863_ ),
    .Y(\u_cpu.ALU.u_wallace._3864_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9368_  (.A(\u_cpu.ALU.u_wallace._3552_ ),
    .B(\u_cpu.ALU.u_wallace._3554_ ),
    .C(\u_cpu.ALU.u_wallace._3860_ ),
    .D(\u_cpu.ALU.u_wallace._3863_ ),
    .X(\u_cpu.ALU.u_wallace._3866_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._9369_  (.A1(\u_cpu.ALU.u_wallace._3851_ ),
    .A2(\u_cpu.ALU.u_wallace._3853_ ),
    .B1(\u_cpu.ALU.u_wallace._3864_ ),
    .C1(\u_cpu.ALU.u_wallace._3866_ ),
    .X(\u_cpu.ALU.u_wallace._3867_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9370_  (.A1(\u_cpu.ALU.u_wallace._3864_ ),
    .A2(\u_cpu.ALU.u_wallace._3866_ ),
    .B1(\u_cpu.ALU.u_wallace._3851_ ),
    .C1(\u_cpu.ALU.u_wallace._3853_ ),
    .Y(\u_cpu.ALU.u_wallace._3868_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9371_  (.A(\u_cpu.ALU.u_wallace._3830_ ),
    .B(\u_cpu.ALU.u_wallace._3867_ ),
    .C(\u_cpu.ALU.u_wallace._3868_ ),
    .Y(\u_cpu.ALU.u_wallace._3869_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9372_  (.A1(\u_cpu.ALU.u_wallace._3552_ ),
    .A2(\u_cpu.ALU.u_wallace._3554_ ),
    .B1(\u_cpu.ALU.u_wallace._3860_ ),
    .B2(\u_cpu.ALU.u_wallace._3863_ ),
    .X(\u_cpu.ALU.u_wallace._3870_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9373_  (.A(\u_cpu.ALU.u_wallace._3552_ ),
    .B(\u_cpu.ALU.u_wallace._3554_ ),
    .C(\u_cpu.ALU.u_wallace._3860_ ),
    .D(\u_cpu.ALU.u_wallace._3863_ ),
    .Y(\u_cpu.ALU.u_wallace._3871_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9374_  (.A(\u_cpu.ALU.u_wallace._3870_ ),
    .B(\u_cpu.ALU.u_wallace._3871_ ),
    .Y(\u_cpu.ALU.u_wallace._3872_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9375_  (.A1(\u_cpu.ALU.u_wallace._3851_ ),
    .A2(\u_cpu.ALU.u_wallace._3853_ ),
    .B1(\u_cpu.ALU.u_wallace._3872_ ),
    .Y(\u_cpu.ALU.u_wallace._3873_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9376_  (.A1(\u_cpu.ALU.u_wallace._3864_ ),
    .A2(\u_cpu.ALU.u_wallace._3866_ ),
    .B1(\u_cpu.ALU.u_wallace._3851_ ),
    .C1(\u_cpu.ALU.u_wallace._3853_ ),
    .X(\u_cpu.ALU.u_wallace._3874_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9377_  (.A1(\u_cpu.ALU.u_wallace._3873_ ),
    .A2(\u_cpu.ALU.u_wallace._3874_ ),
    .B1(\u_cpu.ALU.u_wallace._3389_ ),
    .C1(\u_cpu.ALU.u_wallace._3512_ ),
    .Y(\u_cpu.ALU.u_wallace._3875_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._9378_  (.A1(\u_cpu.ALU.u_wallace._3563_ ),
    .A2(\u_cpu.ALU.u_wallace._3543_ ),
    .A3(\u_cpu.ALU.u_wallace._3566_ ),
    .B1(\u_cpu.ALU.u_wallace._3560_ ),
    .X(\u_cpu.ALU.u_wallace._3877_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9379_  (.A1(\u_cpu.ALU.u_wallace._3869_ ),
    .A2(\u_cpu.ALU.u_wallace._3875_ ),
    .B1(\u_cpu.ALU.u_wallace._3877_ ),
    .Y(\u_cpu.ALU.u_wallace._3878_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9380_  (.A(\u_cpu.ALU.u_wallace._3877_ ),
    .B(\u_cpu.ALU.u_wallace._3869_ ),
    .C(\u_cpu.ALU.u_wallace._3875_ ),
    .X(\u_cpu.ALU.u_wallace._3879_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9381_  (.A(\u_cpu.ALU.u_wallace._3878_ ),
    .B(\u_cpu.ALU.u_wallace._3879_ ),
    .Y(\u_cpu.ALU.u_wallace._3880_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9382_  (.A1(\u_cpu.ALU.u_wallace._3816_ ),
    .A2(\u_cpu.ALU.u_wallace._3827_ ),
    .B1(\u_cpu.ALU.u_wallace._3880_ ),
    .Y(\u_cpu.ALU.u_wallace._3881_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9383_  (.A(\u_cpu.ALU.u_wallace._3880_ ),
    .B(\u_cpu.ALU.u_wallace._3816_ ),
    .C(\u_cpu.ALU.u_wallace._3827_ ),
    .X(\u_cpu.ALU.u_wallace._3882_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._9384_  (.A1(\u_cpu.ALU.u_wallace._3517_ ),
    .A2(\u_cpu.ALU.u_wallace._3511_ ),
    .A3(\u_cpu.ALU.u_wallace._3513_ ),
    .B1(\u_cpu.ALU.u_wallace._3521_ ),
    .B2(\u_cpu.ALU.u_wallace._3583_ ),
    .X(\u_cpu.ALU.u_wallace._3883_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._9385_  (.A1(\u_cpu.ALU.u_wallace._3881_ ),
    .A2(\u_cpu.ALU.u_wallace._3882_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3883_ ),
    .Y(\u_cpu.ALU.u_wallace._3884_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9386_  (.A1(\u_cpu.ALU.u_wallace._3505_ ),
    .A2(\u_cpu.ALU.u_wallace._3616_ ),
    .B1(\u_cpu.ALU.u_wallace._3818_ ),
    .B2(\u_cpu.ALU.u_wallace._3822_ ),
    .Y(\u_cpu.ALU.u_wallace._3885_ ));
 sky130_fd_sc_hd__a311o_2 \u_cpu.ALU.u_wallace._9387_  (.A1(\u_cpu.ALU.u_wallace._3818_ ),
    .A2(\u_cpu.ALU.u_wallace._3822_ ),
    .A3(\u_cpu.ALU.u_wallace._3826_ ),
    .B1(\u_cpu.ALU.u_wallace._3878_ ),
    .C1(\u_cpu.ALU.u_wallace._3879_ ),
    .X(\u_cpu.ALU.u_wallace._3886_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.ALU.u_wallace._9388_  (.A1_N(\u_cpu.ALU.u_wallace._3878_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3879_ ),
    .B1(\u_cpu.ALU.u_wallace._3816_ ),
    .B2(\u_cpu.ALU.u_wallace._3827_ ),
    .X(\u_cpu.ALU.u_wallace._3888_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9389_  (.A1(\u_cpu.ALU.u_wallace._3885_ ),
    .A2(\u_cpu.ALU.u_wallace._3886_ ),
    .B1(\u_cpu.ALU.u_wallace._3888_ ),
    .C1(\u_cpu.ALU.u_wallace._3883_ ),
    .Y(\u_cpu.ALU.u_wallace._3889_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._9390_  (.A(\u_cpu.ALU.u_wallace._3570_ ),
    .Y(\u_cpu.ALU.u_wallace._3890_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._9391_  (.A1(\u_cpu.ALU.u_wallace._3884_ ),
    .A2(\u_cpu.ALU.u_wallace._3889_ ),
    .B1(\u_cpu.ALU.u_wallace._3890_ ),
    .C1(\u_cpu.ALU.u_wallace._3582_ ),
    .X(\u_cpu.ALU.u_wallace._3891_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9392_  (.A1(\u_cpu.ALU.u_wallace._3890_ ),
    .A2(\u_cpu.ALU.u_wallace._3582_ ),
    .B1(\u_cpu.ALU.u_wallace._3884_ ),
    .C1(\u_cpu.ALU.u_wallace._3889_ ),
    .Y(\u_cpu.ALU.u_wallace._3892_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9393_  (.A1(\u_cpu.ALU.u_wallace._3596_ ),
    .A2(\u_cpu.ALU.u_wallace._3593_ ),
    .B1(\u_cpu.ALU.u_wallace._3586_ ),
    .X(\u_cpu.ALU.u_wallace._3893_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9394_  (.A1(\u_cpu.ALU.u_wallace._3891_ ),
    .A2(\u_cpu.ALU.u_wallace._3892_ ),
    .B1(\u_cpu.ALU.u_wallace._3893_ ),
    .X(\u_cpu.ALU.u_wallace._3894_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9395_  (.A(\u_cpu.ALU.u_wallace._3893_ ),
    .B(\u_cpu.ALU.u_wallace._3891_ ),
    .C(\u_cpu.ALU.u_wallace._3892_ ),
    .Y(\u_cpu.ALU.u_wallace._3895_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.ALU.u_wallace._9396_  (.A1_N(\u_cpu.ALU.u_wallace._3537_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3565_ ),
    .B1(\u_cpu.ALU.u_wallace._3544_ ),
    .B2(\u_cpu.ALU.u_wallace._3539_ ),
    .X(\u_cpu.ALU.u_wallace._3896_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9397_  (.A1(\u_cpu.ALU.u_wallace._3894_ ),
    .A2(\u_cpu.ALU.u_wallace._3895_ ),
    .B1(\u_cpu.ALU.u_wallace._3896_ ),
    .Y(\u_cpu.ALU.u_wallace._3897_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9398_  (.A(\u_cpu.ALU.u_wallace._3896_ ),
    .B(\u_cpu.ALU.u_wallace._3894_ ),
    .C(\u_cpu.ALU.u_wallace._3895_ ),
    .X(\u_cpu.ALU.u_wallace._3899_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9399_  (.A1(\u_cpu.ALU.u_wallace._3897_ ),
    .A2(\u_cpu.ALU.u_wallace._3899_ ),
    .B1(\u_cpu.ALU.u_wallace._3598_ ),
    .C1(\u_cpu.ALU.u_wallace._3606_ ),
    .Y(\u_cpu.ALU.u_wallace._3900_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._9400_  (.A1(\u_cpu.ALU.u_wallace._3598_ ),
    .A2(\u_cpu.ALU.u_wallace._3606_ ),
    .B1(\u_cpu.ALU.u_wallace._3897_ ),
    .C1(\u_cpu.ALU.u_wallace._3899_ ),
    .X(\u_cpu.ALU.u_wallace._3901_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._9401_  (.A1(\u_cpu.ALU.u_wallace._3335_ ),
    .A2(\u_cpu.ALU.u_wallace._3607_ ),
    .B1(\u_cpu.ALU.u_wallace._3615_ ),
    .C1(\u_cpu.ALU.u_wallace._3900_ ),
    .D1(\u_cpu.ALU.u_wallace._3901_ ),
    .Y(\u_cpu.ALU.u_wallace._3902_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9402_  (.A1(\u_cpu.ALU.u_wallace._3325_ ),
    .A2(\u_cpu.ALU.u_wallace._3326_ ),
    .B1(\u_cpu.ALU.u_wallace._3607_ ),
    .X(\u_cpu.ALU.u_wallace._3903_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9403_  (.A1(\u_cpu.ALU.u_wallace._3903_ ),
    .A2(\u_cpu.ALU.u_wallace._3615_ ),
    .B1(\u_cpu.ALU.u_wallace._3900_ ),
    .B2(\u_cpu.ALU.u_wallace._3901_ ),
    .X(\u_cpu.ALU.u_wallace._3904_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9404_  (.A(\u_cpu.ALU.u_wallace._3902_ ),
    .B(\u_cpu.ALU.u_wallace._3904_ ),
    .Y(\u_cpu.ALU.Product_Wallace[29] ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._9405_  (.A1(\u_cpu.ALU.u_wallace._3903_ ),
    .A2(\u_cpu.ALU.u_wallace._3901_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3900_ ),
    .Y(\u_cpu.ALU.u_wallace._3905_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9406_  (.A(\u_cpu.ALU.u_wallace._3608_ ),
    .B(\u_cpu.ALU.u_wallace._3900_ ),
    .C(\u_cpu.ALU.u_wallace._3901_ ),
    .Y(\u_cpu.ALU.u_wallace._3906_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9407_  (.A1(\u_cpu.ALU.u_wallace._3609_ ),
    .A2(\u_cpu.ALU.u_wallace._3612_ ),
    .B1(\u_cpu.ALU.u_wallace._3906_ ),
    .Y(\u_cpu.ALU.u_wallace._3907_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._9408_  (.A1(\u_cpu.ALU.u_wallace._3896_ ),
    .A2(\u_cpu.ALU.u_wallace._3894_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3895_ ),
    .Y(\u_cpu.ALU.u_wallace._3909_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9409_  (.A1(\u_cpu.ALU.u_wallace._3849_ ),
    .A2(\u_cpu.ALU.u_wallace._3850_ ),
    .B1(\u_cpu.ALU.u_wallace._3847_ ),
    .Y(\u_cpu.ALU.u_wallace._3910_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9410_  (.A(\u_cpu.ALU.u_wallace._3675_ ),
    .B(\u_cpu.ALU.u_wallace._3679_ ),
    .Y(\u_cpu.ALU.u_wallace._3911_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9411_  (.A1(\u_cpu.ALU.u_wallace._3253_ ),
    .A2(\u_cpu.ALU.u_wallace._3258_ ),
    .B1(\u_cpu.ALU.u_wallace._3254_ ),
    .B2(\u_cpu.ALU.u_wallace._2986_ ),
    .X(\u_cpu.ALU.u_wallace._3912_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9412_  (.A(\u_cpu.ALU.u_wallace._3253_ ),
    .B(\u_cpu.ALU.u_wallace._2986_ ),
    .C(\u_cpu.ALU.u_wallace._3258_ ),
    .D(\u_cpu.ALU.u_wallace._3254_ ),
    .Y(\u_cpu.ALU.u_wallace._3913_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9413_  (.A(\u_cpu.ALU.u_wallace._3912_ ),
    .B(\u_cpu.ALU.u_wallace._3913_ ),
    .C(\u_cpu.ALU.u_wallace._1333_ ),
    .D(\u_cpu.ALU.u_wallace._2480_ ),
    .Y(\u_cpu.ALU.u_wallace._3914_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9414_  (.A1(\u_cpu.ALU.u_wallace._3253_ ),
    .A2(\u_cpu.ALU.u_wallace._3258_ ),
    .B1(\u_cpu.ALU.u_wallace._3254_ ),
    .B2(\u_cpu.ALU.u_wallace._2986_ ),
    .Y(\u_cpu.ALU.u_wallace._3915_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9415_  (.A(\u_cpu.ALU.u_wallace._0917_ ),
    .B(\u_cpu.ALU.u_wallace._4541_ ),
    .C(\u_cpu.ALU.u_wallace._3258_ ),
    .D(\u_cpu.ALU.u_wallace._3254_ ),
    .X(\u_cpu.ALU.u_wallace._3916_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9416_  (.A1(\u_cpu.ALU.u_wallace._4813_ ),
    .A2(\u_cpu.ALU.u_wallace._2482_ ),
    .B1(\u_cpu.ALU.u_wallace._3915_ ),
    .B2(\u_cpu.ALU.u_wallace._3916_ ),
    .Y(\u_cpu.ALU.u_wallace._3917_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.ALU.u_wallace._9417_  (.A1(\u_cpu.ALU.u_wallace._0939_ ),
    .A2(\u_cpu.ALU.u_wallace._2482_ ),
    .A3(\u_cpu.ALU.u_wallace._3834_ ),
    .B1(\u_cpu.ALU.u_wallace._3835_ ),
    .Y(\u_cpu.ALU.u_wallace._3918_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9418_  (.A1(\u_cpu.ALU.u_wallace._3914_ ),
    .A2(\u_cpu.ALU.u_wallace._3917_ ),
    .B1(\u_cpu.ALU.u_wallace._3918_ ),
    .Y(\u_cpu.ALU.u_wallace._3920_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9419_  (.A(\u_cpu.ALU.u_wallace._3918_ ),
    .B(\u_cpu.ALU.u_wallace._3914_ ),
    .C(\u_cpu.ALU.u_wallace._3917_ ),
    .X(\u_cpu.ALU.u_wallace._3921_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._9420_  (.A1_N(\u_cpu.ALU.u_wallace._0198_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2402_ ),
    .B1(\u_cpu.ALU.u_wallace._3920_ ),
    .B2(\u_cpu.ALU.u_wallace._3921_ ),
    .Y(\u_cpu.ALU.u_wallace._3922_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9421_  (.A(\u_cpu.ALU.u_wallace._3918_ ),
    .B(\u_cpu.ALU.u_wallace._3914_ ),
    .C(\u_cpu.ALU.u_wallace._3917_ ),
    .Y(\u_cpu.ALU.u_wallace._3923_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.ALU.u_wallace._9422_  (.A_N(\u_cpu.ALU.u_wallace._3920_ ),
    .B(\u_cpu.ALU.u_wallace._3923_ ),
    .C(\u_cpu.ALU.u_wallace._0198_ ),
    .D(\u_cpu.ALU.u_wallace._2402_ ),
    .Y(\u_cpu.ALU.u_wallace._3924_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._9423_  (.A1(\u_cpu.ALU.u_wallace._3844_ ),
    .A2(\u_cpu.ALU.u_wallace._2402_ ),
    .A3(\u_cpu.ALU.u_wallace._1333_ ),
    .B1(\u_cpu.ALU.u_wallace._3841_ ),
    .X(\u_cpu.ALU.u_wallace._3925_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9424_  (.A1(\u_cpu.ALU.u_wallace._3922_ ),
    .A2(\u_cpu.ALU.u_wallace._3924_ ),
    .B1(\u_cpu.ALU.u_wallace._3925_ ),
    .X(\u_cpu.ALU.u_wallace._3926_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9425_  (.A(\u_cpu.ALU.u_wallace._3925_ ),
    .B(\u_cpu.ALU.u_wallace._3922_ ),
    .C(\u_cpu.ALU.u_wallace._3924_ ),
    .Y(\u_cpu.ALU.u_wallace._3927_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9426_  (.A(\u_cpu.ALU.u_wallace._2343_ ),
    .B(\u_cpu.ALU.u_wallace._2134_ ),
    .Y(\u_cpu.ALU.u_wallace._3928_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9427_  (.A1(\u_cpu.ALU.u_wallace._3926_ ),
    .A2(\u_cpu.ALU.u_wallace._3927_ ),
    .B1(\u_cpu.ALU.u_wallace._3928_ ),
    .Y(\u_cpu.ALU.u_wallace._3929_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9428_  (.A1(\u_cpu.ALU.u_wallace._0203_ ),
    .A2(\u_cpu.ALU.u_wallace._2131_ ),
    .B1(\u_cpu.ALU.u_wallace._3926_ ),
    .C1(\u_cpu.ALU.u_wallace._3927_ ),
    .X(\u_cpu.ALU.u_wallace._3931_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9429_  (.A1(\u_cpu.ALU.u_wallace._0272_ ),
    .A2(\u_cpu.ALU.SrcB[29] ),
    .B1(\u_cpu.ALU.SrcB[30] ),
    .B2(\u_cpu.ALU.u_wallace._1070_ ),
    .X(\u_cpu.ALU.u_wallace._3932_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9430_  (.A(\u_cpu.ALU.u_wallace._0118_ ),
    .B(\u_cpu.ALU.u_wallace._0272_ ),
    .C(\u_cpu.ALU.SrcB[29] ),
    .D(\u_cpu.ALU.SrcB[30] ),
    .Y(\u_cpu.ALU.u_wallace._3933_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9431_  (.A(\u_cpu.ALU.u_wallace._3932_ ),
    .B(\u_cpu.ALU.u_wallace._3933_ ),
    .C(\u_cpu.ALU.u_wallace._0370_ ),
    .D(\u_cpu.ALU.SrcB[28] ),
    .Y(\u_cpu.ALU.u_wallace._3934_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9432_  (.A1(\u_cpu.ALU.u_wallace._0173_ ),
    .A2(\u_cpu.ALU.SrcB[29] ),
    .B1(\u_cpu.ALU.SrcB[30] ),
    .B2(\u_cpu.ALU.u_wallace._0118_ ),
    .Y(\u_cpu.ALU.u_wallace._3935_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9433_  (.A(\u_cpu.ALU.u_wallace._1070_ ),
    .B(\u_cpu.ALU.u_wallace._0272_ ),
    .C(\u_cpu.ALU.SrcB[29] ),
    .D(\u_cpu.ALU.SrcB[30] ),
    .X(\u_cpu.ALU.u_wallace._3936_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9434_  (.A1(\u_cpu.ALU.u_wallace._0414_ ),
    .A2(\u_cpu.ALU.u_wallace._3549_ ),
    .B1(\u_cpu.ALU.u_wallace._3935_ ),
    .B2(\u_cpu.ALU.u_wallace._3936_ ),
    .Y(\u_cpu.ALU.u_wallace._3937_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9435_  (.A(\u_cpu.ALU.u_wallace._2343_ ),
    .B(\u_cpu.ALU.u_wallace._1855_ ),
    .Y(\u_cpu.ALU.u_wallace._3938_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9436_  (.A(\u_cpu.ALU.u_wallace._4661_ ),
    .B(\u_cpu.ALU.u_wallace._1611_ ),
    .Y(\u_cpu.ALU.u_wallace._3939_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._9437_  (.A1_N(\u_cpu.ALU.u_wallace._3934_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3937_ ),
    .B1(\u_cpu.ALU.u_wallace._3938_ ),
    .B2(\u_cpu.ALU.u_wallace._3939_ ),
    .Y(\u_cpu.ALU.u_wallace._3940_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9438_  (.A(\u_cpu.ALU.u_wallace._3937_ ),
    .B(\u_cpu.ALU.u_wallace._3631_ ),
    .C(\u_cpu.ALU.u_wallace._3934_ ),
    .Y(\u_cpu.ALU.u_wallace._3942_ ));
 sky130_fd_sc_hd__a21bo_2 \u_cpu.ALU.u_wallace._9439_  (.A1(\u_cpu.ALU.u_wallace._3940_ ),
    .A2(\u_cpu.ALU.u_wallace._3942_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3856_ ),
    .X(\u_cpu.ALU.u_wallace._3943_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9440_  (.A(\u_cpu.ALU.u_wallace._0129_ ),
    .B(\u_cpu.ALU.u_wallace._0184_ ),
    .C(\u_cpu.ALU.SrcB[29] ),
    .Y(\u_cpu.ALU.u_wallace._3944_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9441_  (.A1(\u_cpu.ALU.u_wallace._3549_ ),
    .A2(\u_cpu.ALU.u_wallace._3944_ ),
    .B1(\u_cpu.ALU.u_wallace._3940_ ),
    .C1(\u_cpu.ALU.u_wallace._3942_ ),
    .Y(\u_cpu.ALU.u_wallace._3945_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9442_  (.A(\u_cpu.ALU.u_wallace._3624_ ),
    .B(\u_cpu.ALU.u_wallace._1615_ ),
    .C(\u_cpu.ALU.u_wallace._0607_ ),
    .D(\u_cpu.ALU.u_wallace._3625_ ),
    .X(\u_cpu.ALU.u_wallace._3946_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9443_  (.A(\u_cpu.ALU.u_wallace._3628_ ),
    .B(\u_cpu.ALU.u_wallace._3622_ ),
    .Y(\u_cpu.ALU.u_wallace._3947_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU.u_wallace._9444_  (.A(\u_cpu.ALU.u_wallace._3631_ ),
    .B(\u_cpu.ALU.u_wallace._3632_ ),
    .X(\u_cpu.ALU.u_wallace._3948_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._9445_  (.A1(\u_cpu.ALU.u_wallace._3946_ ),
    .A2(\u_cpu.ALU.u_wallace._3947_ ),
    .B1(\u_cpu.ALU.u_wallace._3948_ ),
    .B2(\u_cpu.ALU.u_wallace._3629_ ),
    .X(\u_cpu.ALU.u_wallace._3949_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9446_  (.A(\u_cpu.ALU.u_wallace._3943_ ),
    .B(\u_cpu.ALU.u_wallace._3945_ ),
    .C(\u_cpu.ALU.u_wallace._3949_ ),
    .Y(\u_cpu.ALU.u_wallace._3950_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9447_  (.A(\u_cpu.ALU.u_wallace._3622_ ),
    .B(\u_cpu.ALU.u_wallace._3626_ ),
    .Y(\u_cpu.ALU.u_wallace._3951_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._9448_  (.A1(\u_cpu.ALU.u_wallace._4677_ ),
    .A2(\u_cpu.ALU.u_wallace._2053_ ),
    .A3(\u_cpu.ALU.u_wallace._3364_ ),
    .B1(\u_cpu.ALU.u_wallace._3365_ ),
    .X(\u_cpu.ALU.u_wallace._3953_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9449_  (.A1(\u_cpu.ALU.u_wallace._3951_ ),
    .A2(\u_cpu.ALU.u_wallace._3953_ ),
    .B1(\u_cpu.ALU.u_wallace._3948_ ),
    .Y(\u_cpu.ALU.u_wallace._3954_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9450_  (.A(\u_cpu.ALU.u_wallace._3940_ ),
    .B(\u_cpu.ALU.u_wallace._3942_ ),
    .C(\u_cpu.ALU.u_wallace._3856_ ),
    .Y(\u_cpu.ALU.u_wallace._3955_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._9451_  (.A1_N(\u_cpu.ALU.u_wallace._3940_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3942_ ),
    .B1(\u_cpu.ALU.u_wallace._3549_ ),
    .B2(\u_cpu.ALU.u_wallace._3944_ ),
    .Y(\u_cpu.ALU.u_wallace._3956_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9452_  (.A1(\u_cpu.ALU.u_wallace._3630_ ),
    .A2(\u_cpu.ALU.u_wallace._3954_ ),
    .B1(\u_cpu.ALU.u_wallace._3955_ ),
    .C1(\u_cpu.ALU.u_wallace._3956_ ),
    .Y(\u_cpu.ALU.u_wallace._3957_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9453_  (.A1(\u_cpu.ALU.u_wallace._3950_ ),
    .A2(\u_cpu.ALU.u_wallace._3957_ ),
    .B1(\u_cpu.ALU.u_wallace._3858_ ),
    .Y(\u_cpu.ALU.u_wallace._3958_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._9454_  (.A1(\u_cpu.ALU.u_wallace._3857_ ),
    .A2(\u_cpu.ALU.u_wallace._3858_ ),
    .B1(\u_cpu.ALU.u_wallace._3363_ ),
    .B2(\u_cpu.ALU.u_wallace._3859_ ),
    .C1(\u_cpu.ALU.u_wallace._3372_ ),
    .X(\u_cpu.ALU.u_wallace._3959_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9455_  (.A1(\u_cpu.ALU.u_wallace._3552_ ),
    .A2(\u_cpu.ALU.u_wallace._3863_ ),
    .B1(\u_cpu.ALU.u_wallace._3959_ ),
    .Y(\u_cpu.ALU.u_wallace._3960_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9456_  (.A(\u_cpu.ALU.u_wallace._3950_ ),
    .B(\u_cpu.ALU.u_wallace._3957_ ),
    .C(\u_cpu.ALU.u_wallace._3858_ ),
    .Y(\u_cpu.ALU.u_wallace._3961_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._9457_  (.A_N(\u_cpu.ALU.u_wallace._3958_ ),
    .B(\u_cpu.ALU.u_wallace._3960_ ),
    .C(\u_cpu.ALU.u_wallace._3961_ ),
    .Y(\u_cpu.ALU.u_wallace._3962_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._9458_  (.A1(\u_cpu.ALU.u_wallace._0043_ ),
    .A2(\u_cpu.ALU.u_wallace._3549_ ),
    .A3(\u_cpu.ALU.u_wallace._3550_ ),
    .B1(\u_cpu.ALU.u_wallace._3863_ ),
    .X(\u_cpu.ALU.u_wallace._3964_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9459_  (.A(\u_cpu.ALU.u_wallace._3950_ ),
    .B(\u_cpu.ALU.u_wallace._3957_ ),
    .C(\u_cpu.ALU.u_wallace._3858_ ),
    .X(\u_cpu.ALU.u_wallace._3965_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9460_  (.A1(\u_cpu.ALU.u_wallace._3959_ ),
    .A2(\u_cpu.ALU.u_wallace._3964_ ),
    .B1(\u_cpu.ALU.u_wallace._3965_ ),
    .B2(\u_cpu.ALU.u_wallace._3958_ ),
    .Y(\u_cpu.ALU.u_wallace._3966_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9461_  (.A1(\u_cpu.ALU.u_wallace._3929_ ),
    .A2(\u_cpu.ALU.u_wallace._3931_ ),
    .B1(\u_cpu.ALU.u_wallace._3962_ ),
    .C1(\u_cpu.ALU.u_wallace._3966_ ),
    .Y(\u_cpu.ALU.u_wallace._3967_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9462_  (.A1(\u_cpu.ALU.u_wallace._3926_ ),
    .A2(\u_cpu.ALU.u_wallace._3927_ ),
    .B1(\u_cpu.ALU.u_wallace._3928_ ),
    .X(\u_cpu.ALU.u_wallace._3968_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9463_  (.A1(\u_cpu.ALU.u_wallace._0203_ ),
    .A2(\u_cpu.ALU.u_wallace._2131_ ),
    .B1(\u_cpu.ALU.u_wallace._3926_ ),
    .C1(\u_cpu.ALU.u_wallace._3927_ ),
    .Y(\u_cpu.ALU.u_wallace._3969_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9464_  (.A(\u_cpu.ALU.u_wallace._3968_ ),
    .B(\u_cpu.ALU.u_wallace._3969_ ),
    .Y(\u_cpu.ALU.u_wallace._3970_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9465_  (.A1(\u_cpu.ALU.u_wallace._3962_ ),
    .A2(\u_cpu.ALU.u_wallace._3966_ ),
    .B1(\u_cpu.ALU.u_wallace._3970_ ),
    .X(\u_cpu.ALU.u_wallace._3971_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9466_  (.A(\u_cpu.ALU.u_wallace._3911_ ),
    .B(\u_cpu.ALU.u_wallace._3967_ ),
    .C(\u_cpu.ALU.u_wallace._3971_ ),
    .Y(\u_cpu.ALU.u_wallace._3972_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9467_  (.A1(\u_cpu.ALU.u_wallace._3929_ ),
    .A2(\u_cpu.ALU.u_wallace._3931_ ),
    .B1(\u_cpu.ALU.u_wallace._3962_ ),
    .C1(\u_cpu.ALU.u_wallace._3966_ ),
    .X(\u_cpu.ALU.u_wallace._3973_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9468_  (.A1(\u_cpu.ALU.u_wallace._3962_ ),
    .A2(\u_cpu.ALU.u_wallace._3966_ ),
    .B1(\u_cpu.ALU.u_wallace._3970_ ),
    .Y(\u_cpu.ALU.u_wallace._3975_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._9469_  (.A1(\u_cpu.ALU.u_wallace._3676_ ),
    .A2(\u_cpu.ALU.u_wallace._3670_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3675_ ),
    .Y(\u_cpu.ALU.u_wallace._3976_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9470_  (.A1(\u_cpu.ALU.u_wallace._3973_ ),
    .A2(\u_cpu.ALU.u_wallace._3975_ ),
    .B1(\u_cpu.ALU.u_wallace._3976_ ),
    .Y(\u_cpu.ALU.u_wallace._3977_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.ALU.u_wallace._9471_  (.A_N(\u_cpu.ALU.u_wallace._3556_ ),
    .B(\u_cpu.ALU.u_wallace._3860_ ),
    .C(\u_cpu.ALU.u_wallace._3863_ ),
    .D(\u_cpu.ALU.u_wallace._3548_ ),
    .X(\u_cpu.ALU.u_wallace._3978_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._9472_  (.A1(\u_cpu.ALU.u_wallace._3872_ ),
    .A2(\u_cpu.ALU.u_wallace._3851_ ),
    .A3(\u_cpu.ALU.u_wallace._3853_ ),
    .B1(\u_cpu.ALU.u_wallace._3978_ ),
    .X(\u_cpu.ALU.u_wallace._3979_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9473_  (.A1(\u_cpu.ALU.u_wallace._3972_ ),
    .A2(\u_cpu.ALU.u_wallace._3977_ ),
    .B1(\u_cpu.ALU.u_wallace._3979_ ),
    .Y(\u_cpu.ALU.u_wallace._3980_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9474_  (.A(\u_cpu.ALU.u_wallace._3979_ ),
    .B(\u_cpu.ALU.u_wallace._3972_ ),
    .C(\u_cpu.ALU.u_wallace._3977_ ),
    .X(\u_cpu.ALU.u_wallace._3981_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9475_  (.A1(\u_cpu.ALU.u_wallace._0607_ ),
    .A2(\u_cpu.ALU.u_wallace._1611_ ),
    .B1(\u_cpu.ALU.u_wallace._1855_ ),
    .B2(\u_cpu.ALU.u_wallace._4661_ ),
    .Y(\u_cpu.ALU.u_wallace._3982_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9476_  (.A(\u_cpu.ALU.u_wallace._4661_ ),
    .B(\u_cpu.ALU.u_wallace._0607_ ),
    .C(\u_cpu.ALU.u_wallace._1611_ ),
    .D(\u_cpu.ALU.u_wallace._1855_ ),
    .X(\u_cpu.ALU.u_wallace._3983_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9477_  (.A1(\u_cpu.ALU.u_wallace._2658_ ),
    .A2(\u_cpu.ALU.u_wallace._0959_ ),
    .B1(\u_cpu.ALU.u_wallace._1176_ ),
    .B2(\u_cpu.ALU.u_wallace._1129_ ),
    .X(\u_cpu.ALU.u_wallace._3984_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9478_  (.A(\u_cpu.ALU.u_wallace._1129_ ),
    .B(\u_cpu.ALU.u_wallace._2658_ ),
    .C(\u_cpu.ALU.u_wallace._0959_ ),
    .D(\u_cpu.ALU.u_wallace._1176_ ),
    .Y(\u_cpu.ALU.u_wallace._3986_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9479_  (.A(\u_cpu.ALU.u_wallace._3984_ ),
    .B(\u_cpu.ALU.u_wallace._3986_ ),
    .C(\u_cpu.ALU.u_wallace._0847_ ),
    .D(\u_cpu.ALU.u_wallace._1615_ ),
    .Y(\u_cpu.ALU.u_wallace._3987_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._9480_  (.A1_N(\u_cpu.ALU.u_wallace._3984_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3986_ ),
    .B1(\u_cpu.ALU.u_wallace._4904_ ),
    .B2(\u_cpu.ALU.u_wallace._2053_ ),
    .Y(\u_cpu.ALU.u_wallace._3988_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9481_  (.A(\u_cpu.ALU.u_wallace._0847_ ),
    .B(\u_cpu.ALU.u_wallace._1129_ ),
    .C(\u_cpu.ALU.u_wallace._0959_ ),
    .D(\u_cpu.ALU.u_wallace._1176_ ),
    .X(\u_cpu.ALU.u_wallace._3989_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._9482_  (.A1(\u_cpu.ALU.u_wallace._3624_ ),
    .A2(\u_cpu.ALU.u_wallace._1615_ ),
    .A3(\u_cpu.ALU.u_wallace._0607_ ),
    .B1(\u_cpu.ALU.u_wallace._3989_ ),
    .X(\u_cpu.ALU.u_wallace._3990_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9483_  (.A1(\u_cpu.ALU.u_wallace._3987_ ),
    .A2(\u_cpu.ALU.u_wallace._3988_ ),
    .B1(\u_cpu.ALU.u_wallace._3990_ ),
    .Y(\u_cpu.ALU.u_wallace._3991_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9484_  (.A(\u_cpu.ALU.u_wallace._3990_ ),
    .B(\u_cpu.ALU.u_wallace._3987_ ),
    .C(\u_cpu.ALU.u_wallace._3988_ ),
    .X(\u_cpu.ALU.u_wallace._3992_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9485_  (.A1(\u_cpu.ALU.u_wallace._3982_ ),
    .A2(\u_cpu.ALU.u_wallace._3983_ ),
    .B1(\u_cpu.ALU.u_wallace._3991_ ),
    .B2(\u_cpu.ALU.u_wallace._3992_ ),
    .Y(\u_cpu.ALU.u_wallace._3993_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9486_  (.A1(\u_cpu.ALU.u_wallace._3989_ ),
    .A2(\u_cpu.ALU.u_wallace._3946_ ),
    .B1(\u_cpu.ALU.u_wallace._3987_ ),
    .C1(\u_cpu.ALU.u_wallace._3988_ ),
    .Y(\u_cpu.ALU.u_wallace._3994_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9487_  (.A(\u_cpu.ALU.u_wallace._3982_ ),
    .B(\u_cpu.ALU.u_wallace._3983_ ),
    .Y(\u_cpu.ALU.u_wallace._3995_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._9488_  (.A_N(\u_cpu.ALU.u_wallace._3991_ ),
    .B(\u_cpu.ALU.u_wallace._3994_ ),
    .C(\u_cpu.ALU.u_wallace._3995_ ),
    .Y(\u_cpu.ALU.u_wallace._3997_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9489_  (.A(\u_cpu.ALU.u_wallace._0122_ ),
    .B(\u_cpu.ALU.u_wallace._1974_ ),
    .Y(\u_cpu.ALU.u_wallace._3998_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9490_  (.A(\u_cpu.ALU.u_wallace._0280_ ),
    .B(\u_cpu.ALU.u_wallace._2248_ ),
    .Y(\u_cpu.ALU.u_wallace._3999_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._9491_  (.A(\u_cpu.ALU.u_wallace._0652_ ),
    .B(\u_cpu.ALU.u_wallace._3204_ ),
    .X(\u_cpu.ALU.u_wallace._4000_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9492_  (.A1(\u_cpu.ALU.u_wallace._1974_ ),
    .A2(\u_cpu.ALU.u_wallace._0280_ ),
    .B1(\u_cpu.ALU.u_wallace._2248_ ),
    .B2(\u_cpu.ALU.u_wallace._0122_ ),
    .X(\u_cpu.ALU.u_wallace._4001_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9493_  (.A1(\u_cpu.ALU.u_wallace._3998_ ),
    .A2(\u_cpu.ALU.u_wallace._3999_ ),
    .B1(\u_cpu.ALU.u_wallace._4000_ ),
    .C1(\u_cpu.ALU.u_wallace._4001_ ),
    .X(\u_cpu.ALU.u_wallace._4002_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9494_  (.A1(\u_cpu.ALU.u_wallace._1974_ ),
    .A2(\u_cpu.ALU.u_wallace._0280_ ),
    .B1(\u_cpu.ALU.u_wallace._2248_ ),
    .B2(\u_cpu.ALU.u_wallace._0122_ ),
    .Y(\u_cpu.ALU.u_wallace._4003_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9495_  (.A(\u_cpu.ALU.u_wallace._0122_ ),
    .B(\u_cpu.ALU.u_wallace._1974_ ),
    .C(\u_cpu.ALU.u_wallace._0280_ ),
    .D(\u_cpu.ALU.u_wallace._2248_ ),
    .X(\u_cpu.ALU.u_wallace._4004_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._9496_  (.A1(\u_cpu.ALU.u_wallace._1323_ ),
    .A2(\u_cpu.ALU.u_wallace._0554_ ),
    .B1(\u_cpu.ALU.u_wallace._4003_ ),
    .B2(\u_cpu.ALU.u_wallace._4004_ ),
    .X(\u_cpu.ALU.u_wallace._4005_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9497_  (.A1(\u_cpu.ALU.u_wallace._3705_ ),
    .A2(\u_cpu.ALU.u_wallace._3701_ ),
    .B1(\u_cpu.ALU.u_wallace._3697_ ),
    .Y(\u_cpu.ALU.u_wallace._4006_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._9498_  (.A1(\u_cpu.ALU.u_wallace._4002_ ),
    .A2(\u_cpu.ALU.u_wallace._4005_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4006_ ),
    .Y(\u_cpu.ALU.u_wallace._4008_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._9499_  (.A1(\u_cpu.ALU.u_wallace._3998_ ),
    .A2(\u_cpu.ALU.u_wallace._3999_ ),
    .B1(\u_cpu.ALU.u_wallace._0652_ ),
    .C1(\u_cpu.ALU.u_wallace._3204_ ),
    .D1(\u_cpu.ALU.u_wallace._4001_ ),
    .Y(\u_cpu.ALU.u_wallace._4009_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9500_  (.A1(\u_cpu.ALU.u_wallace._1323_ ),
    .A2(\u_cpu.ALU.u_wallace._0554_ ),
    .B1(\u_cpu.ALU.u_wallace._4003_ ),
    .B2(\u_cpu.ALU.u_wallace._4004_ ),
    .Y(\u_cpu.ALU.u_wallace._4010_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9501_  (.A(\u_cpu.ALU.u_wallace._4006_ ),
    .B(\u_cpu.ALU.u_wallace._4009_ ),
    .C(\u_cpu.ALU.u_wallace._4010_ ),
    .Y(\u_cpu.ALU.u_wallace._4011_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._9502_  (.A1(\u_cpu.ALU.u_wallace._3641_ ),
    .A2(\u_cpu.ALU.u_wallace._3204_ ),
    .A3(\u_cpu.ALU.u_wallace._1578_ ),
    .B1(\u_cpu.ALU.u_wallace._3646_ ),
    .X(\u_cpu.ALU.u_wallace._4012_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9503_  (.A1(\u_cpu.ALU.u_wallace._4008_ ),
    .A2(\u_cpu.ALU.u_wallace._4011_ ),
    .B1(\u_cpu.ALU.u_wallace._4012_ ),
    .Y(\u_cpu.ALU.u_wallace._4013_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9504_  (.A(\u_cpu.ALU.u_wallace._3641_ ),
    .B(\u_cpu.ALU.u_wallace._3642_ ),
    .C(\u_cpu.ALU.u_wallace._1578_ ),
    .D(\u_cpu.ALU.u_wallace._3204_ ),
    .X(\u_cpu.ALU.u_wallace._4014_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9505_  (.A1(\u_cpu.ALU.u_wallace._3646_ ),
    .A2(\u_cpu.ALU.u_wallace._4014_ ),
    .B1(\u_cpu.ALU.u_wallace._4008_ ),
    .C1(\u_cpu.ALU.u_wallace._4011_ ),
    .X(\u_cpu.ALU.u_wallace._4015_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._9506_  (.A1(\u_cpu.ALU.u_wallace._3657_ ),
    .A2(\u_cpu.ALU.u_wallace._3655_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3648_ ),
    .Y(\u_cpu.ALU.u_wallace._4016_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._9507_  (.A1(\u_cpu.ALU.u_wallace._4013_ ),
    .A2(\u_cpu.ALU.u_wallace._4015_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4016_ ),
    .Y(\u_cpu.ALU.u_wallace._4017_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9508_  (.A1(\u_cpu.ALU.u_wallace._4009_ ),
    .A2(\u_cpu.ALU.u_wallace._4010_ ),
    .B1(\u_cpu.ALU.u_wallace._4006_ ),
    .Y(\u_cpu.ALU.u_wallace._4019_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9509_  (.A1(\u_cpu.ALU.u_wallace._3696_ ),
    .A2(\u_cpu.ALU.u_wallace._3698_ ),
    .B1(\u_cpu.ALU.u_wallace._3702_ ),
    .Y(\u_cpu.ALU.u_wallace._4020_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._9510_  (.A(\u_cpu.ALU.u_wallace._4020_ ),
    .B(\u_cpu.ALU.u_wallace._4002_ ),
    .C(\u_cpu.ALU.u_wallace._4005_ ),
    .Y(\u_cpu.ALU.u_wallace._4021_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._9511_  (.A1(\u_cpu.ALU.u_wallace._4019_ ),
    .A2(\u_cpu.ALU.u_wallace._4021_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4012_ ),
    .Y(\u_cpu.ALU.u_wallace._4022_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9512_  (.A1(\u_cpu.ALU.u_wallace._3646_ ),
    .A2(\u_cpu.ALU.u_wallace._4014_ ),
    .B1(\u_cpu.ALU.u_wallace._4008_ ),
    .C1(\u_cpu.ALU.u_wallace._4011_ ),
    .Y(\u_cpu.ALU.u_wallace._4023_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9513_  (.A1(\u_cpu.ALU.u_wallace._3648_ ),
    .A2(\u_cpu.ALU.u_wallace._3661_ ),
    .B1(\u_cpu.ALU.u_wallace._4022_ ),
    .C1(\u_cpu.ALU.u_wallace._4023_ ),
    .Y(\u_cpu.ALU.u_wallace._4024_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9514_  (.A1(\u_cpu.ALU.u_wallace._3993_ ),
    .A2(\u_cpu.ALU.u_wallace._3997_ ),
    .B1(\u_cpu.ALU.u_wallace._4017_ ),
    .B2(\u_cpu.ALU.u_wallace._4024_ ),
    .Y(\u_cpu.ALU.u_wallace._4025_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._9515_  (.A1(\u_cpu.ALU.u_wallace._3648_ ),
    .A2(\u_cpu.ALU.u_wallace._3661_ ),
    .B1(\u_cpu.ALU.u_wallace._4023_ ),
    .X(\u_cpu.ALU.u_wallace._4026_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9516_  (.A(\u_cpu.ALU.u_wallace._3993_ ),
    .B(\u_cpu.ALU.u_wallace._3997_ ),
    .Y(\u_cpu.ALU.u_wallace._4027_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9517_  (.A1(\u_cpu.ALU.u_wallace._4022_ ),
    .A2(\u_cpu.ALU.u_wallace._4023_ ),
    .B1(\u_cpu.ALU.u_wallace._4016_ ),
    .Y(\u_cpu.ALU.u_wallace._4028_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU.u_wallace._9518_  (.A1(\u_cpu.ALU.u_wallace._4026_ ),
    .A2(\u_cpu.ALU.u_wallace._4022_ ),
    .B1(\u_cpu.ALU.u_wallace._4027_ ),
    .C1(\u_cpu.ALU.u_wallace._4028_ ),
    .Y(\u_cpu.ALU.u_wallace._4030_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9519_  (.A1(\u_cpu.ALU.u_wallace._3716_ ),
    .A2(\u_cpu.ALU.u_wallace._3715_ ),
    .B1(\u_cpu.ALU.u_wallace._3801_ ),
    .Y(\u_cpu.ALU.u_wallace._4031_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._9520_  (.A1(\u_cpu.ALU.u_wallace._4025_ ),
    .A2(\u_cpu.ALU.u_wallace._4030_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4031_ ),
    .Y(\u_cpu.ALU.u_wallace._4032_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9521_  (.A1(\u_cpu.ALU.u_wallace._3648_ ),
    .A2(\u_cpu.ALU.u_wallace._3661_ ),
    .B1(\u_cpu.ALU.u_wallace._4022_ ),
    .C1(\u_cpu.ALU.u_wallace._4023_ ),
    .X(\u_cpu.ALU.u_wallace._4033_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._9522_  (.A1_N(\u_cpu.ALU.u_wallace._3993_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3997_ ),
    .B1(\u_cpu.ALU.u_wallace._4028_ ),
    .B2(\u_cpu.ALU.u_wallace._4033_ ),
    .Y(\u_cpu.ALU.u_wallace._4034_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9523_  (.A(\u_cpu.ALU.u_wallace._3993_ ),
    .B(\u_cpu.ALU.u_wallace._3997_ ),
    .C(\u_cpu.ALU.u_wallace._4017_ ),
    .D(\u_cpu.ALU.u_wallace._4024_ ),
    .Y(\u_cpu.ALU.u_wallace._4035_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9524_  (.A(\u_cpu.ALU.u_wallace._4031_ ),
    .B(\u_cpu.ALU.u_wallace._4034_ ),
    .C(\u_cpu.ALU.u_wallace._4035_ ),
    .Y(\u_cpu.ALU.u_wallace._4036_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._9525_  (.A1(\u_cpu.ALU.u_wallace._3666_ ),
    .A2(\u_cpu.ALU.u_wallace._3663_ ),
    .B1(\u_cpu.ALU.u_wallace._3668_ ),
    .X(\u_cpu.ALU.u_wallace._4037_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._9526_  (.A1(\u_cpu.ALU.u_wallace._4032_ ),
    .A2(\u_cpu.ALU.u_wallace._4036_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4037_ ),
    .Y(\u_cpu.ALU.u_wallace._4038_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._9527_  (.A1(\u_cpu.ALU.u_wallace._3635_ ),
    .A2(\u_cpu.ALU.u_wallace._3636_ ),
    .B1(\u_cpu.ALU.u_wallace._3665_ ),
    .X(\u_cpu.ALU.u_wallace._4039_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9528_  (.A1(\u_cpu.ALU.u_wallace._3660_ ),
    .A2(\u_cpu.ALU.u_wallace._4039_ ),
    .B1(\u_cpu.ALU.u_wallace._4032_ ),
    .C1(\u_cpu.ALU.u_wallace._4036_ ),
    .X(\u_cpu.ALU.u_wallace._4041_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9529_  (.A1(\u_cpu.ALU.u_wallace._3446_ ),
    .A2(\u_cpu.ALU.u_wallace._3761_ ),
    .B1(\u_cpu.ALU.u_wallace._3764_ ),
    .C1(\u_cpu.ALU.u_wallace._3768_ ),
    .X(\u_cpu.ALU.u_wallace._4042_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._9530_  (.A(\u_cpu.ALU.u_wallace._4605_ ),
    .B(\u_cpu.ALU.u_wallace._3088_ ),
    .X(\u_cpu.ALU.u_wallace._4043_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9531_  (.A1(\u_cpu.ALU.u_wallace._4313_ ),
    .A2(\u_cpu.ALU.u_wallace._2618_ ),
    .B1(\u_cpu.ALU.u_wallace._2598_ ),
    .B2(\u_cpu.ALU.u_wallace._4029_ ),
    .X(\u_cpu.ALU.u_wallace._4044_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9532_  (.A1(\u_cpu.ALU.u_wallace._1737_ ),
    .A2(\u_cpu.ALU.u_wallace._3685_ ),
    .B1(\u_cpu.ALU.u_wallace._4043_ ),
    .C1(\u_cpu.ALU.u_wallace._4044_ ),
    .X(\u_cpu.ALU.u_wallace._4045_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9533_  (.A(\u_cpu.ALU.u_wallace._4029_ ),
    .B(\u_cpu.ALU.u_wallace._4313_ ),
    .C(\u_cpu.ALU.u_wallace._2618_ ),
    .D(\u_cpu.ALU.u_wallace._2598_ ),
    .Y(\u_cpu.ALU.u_wallace._4046_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9534_  (.A1(\u_cpu.ALU.u_wallace._4044_ ),
    .A2(\u_cpu.ALU.u_wallace._4046_ ),
    .B1(\u_cpu.ALU.u_wallace._4043_ ),
    .Y(\u_cpu.ALU.u_wallace._4047_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU.u_wallace._9535_  (.A1_N(\u_cpu.ALU.u_wallace._3692_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3686_ ),
    .B1(\u_cpu.ALU.u_wallace._1271_ ),
    .B2(\u_cpu.ALU.u_wallace._3685_ ),
    .X(\u_cpu.ALU.u_wallace._4048_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9536_  (.A1(\u_cpu.ALU.u_wallace._4045_ ),
    .A2(\u_cpu.ALU.u_wallace._4047_ ),
    .B1(\u_cpu.ALU.u_wallace._4048_ ),
    .Y(\u_cpu.ALU.u_wallace._4049_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.ALU.u_wallace._9537_  (.A1_N(\u_cpu.ALU.u_wallace._1271_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3685_ ),
    .B1(\u_cpu.ALU.u_wallace._3692_ ),
    .B2(\u_cpu.ALU.u_wallace._3686_ ),
    .X(\u_cpu.ALU.u_wallace._4050_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._9538_  (.A1(\u_cpu.ALU.u_wallace._1737_ ),
    .A2(\u_cpu.ALU.u_wallace._3685_ ),
    .B1(\u_cpu.ALU.u_wallace._4605_ ),
    .C1(\u_cpu.ALU.u_wallace._3088_ ),
    .D1(\u_cpu.ALU.u_wallace._4044_ ),
    .Y(\u_cpu.ALU.u_wallace._4052_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9539_  (.A1(\u_cpu.ALU.u_wallace._4605_ ),
    .A2(\u_cpu.ALU.u_wallace._3088_ ),
    .B1(\u_cpu.ALU.u_wallace._4044_ ),
    .B2(\u_cpu.ALU.u_wallace._4046_ ),
    .X(\u_cpu.ALU.u_wallace._4053_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9540_  (.A(\u_cpu.ALU.u_wallace._4050_ ),
    .B(\u_cpu.ALU.u_wallace._4052_ ),
    .C(\u_cpu.ALU.u_wallace._4053_ ),
    .Y(\u_cpu.ALU.u_wallace._4054_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9541_  (.A1(\u_cpu.ALU.u_wallace._4894_ ),
    .A2(\u_cpu.ALU.u_wallace._2916_ ),
    .B1(\u_cpu.ALU.u_wallace._2907_ ),
    .B2(\u_cpu.ALU.u_wallace._4733_ ),
    .Y(\u_cpu.ALU.u_wallace._4055_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9542_  (.A(\u_cpu.ALU.u_wallace._4732_ ),
    .B(\u_cpu.ALU.u_wallace._4894_ ),
    .C(\u_cpu.ALU.u_wallace._2916_ ),
    .D(\u_cpu.ALU.u_wallace._2907_ ),
    .X(\u_cpu.ALU.u_wallace._4056_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9543_  (.A1(\u_cpu.ALU.u_wallace._4055_ ),
    .A2(\u_cpu.ALU.u_wallace._4056_ ),
    .B1(\u_cpu.ALU.u_wallace._0117_ ),
    .C1(\u_cpu.ALU.u_wallace._2621_ ),
    .Y(\u_cpu.ALU.u_wallace._4057_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._9544_  (.A1(\u_cpu.ALU.u_wallace._0117_ ),
    .A2(\u_cpu.ALU.u_wallace._2621_ ),
    .B1(\u_cpu.ALU.u_wallace._4055_ ),
    .C1(\u_cpu.ALU.u_wallace._4056_ ),
    .X(\u_cpu.ALU.u_wallace._4058_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9545_  (.A(\u_cpu.ALU.u_wallace._4057_ ),
    .B(\u_cpu.ALU.u_wallace._4058_ ),
    .Y(\u_cpu.ALU.u_wallace._4059_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9546_  (.A1(\u_cpu.ALU.u_wallace._4049_ ),
    .A2(\u_cpu.ALU.u_wallace._4054_ ),
    .B1(\u_cpu.ALU.u_wallace._4059_ ),
    .X(\u_cpu.ALU.u_wallace._4060_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9547_  (.A(\u_cpu.ALU.u_wallace._4049_ ),
    .B(\u_cpu.ALU.u_wallace._4059_ ),
    .C(\u_cpu.ALU.u_wallace._4054_ ),
    .Y(\u_cpu.ALU.u_wallace._4061_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9548_  (.A1(\u_cpu.ALU.u_wallace._4042_ ),
    .A2(\u_cpu.ALU.u_wallace._3773_ ),
    .B1(\u_cpu.ALU.u_wallace._4060_ ),
    .C1(\u_cpu.ALU.u_wallace._4061_ ),
    .Y(\u_cpu.ALU.u_wallace._4063_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._9549_  (.A(\u_cpu.ALU.u_wallace._4063_ ),
    .Y(\u_cpu.ALU.u_wallace._4064_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9550_  (.A(\u_cpu.ALU.u_wallace._3691_ ),
    .B(\u_cpu.ALU.u_wallace._3708_ ),
    .Y(\u_cpu.ALU.u_wallace._4065_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9551_  (.A1(\u_cpu.ALU.u_wallace._4049_ ),
    .A2(\u_cpu.ALU.u_wallace._4054_ ),
    .B1(\u_cpu.ALU.u_wallace._4059_ ),
    .Y(\u_cpu.ALU.u_wallace._4066_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9552_  (.A(\u_cpu.ALU.u_wallace._4049_ ),
    .B(\u_cpu.ALU.u_wallace._4059_ ),
    .C(\u_cpu.ALU.u_wallace._4054_ ),
    .X(\u_cpu.ALU.u_wallace._4067_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9553_  (.A1(\u_cpu.ALU.u_wallace._3770_ ),
    .A2(\u_cpu.ALU.u_wallace._3772_ ),
    .B1(\u_cpu.ALU.u_wallace._3769_ ),
    .Y(\u_cpu.ALU.u_wallace._4068_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._9554_  (.A1(\u_cpu.ALU.u_wallace._4066_ ),
    .A2(\u_cpu.ALU.u_wallace._4067_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4068_ ),
    .Y(\u_cpu.ALU.u_wallace._4069_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9555_  (.A(\u_cpu.ALU.u_wallace._4065_ ),
    .B(\u_cpu.ALU.u_wallace._4069_ ),
    .Y(\u_cpu.ALU.u_wallace._4070_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9556_  (.A1(\u_cpu.ALU.u_wallace._4063_ ),
    .A2(\u_cpu.ALU.u_wallace._4069_ ),
    .B1(\u_cpu.ALU.u_wallace._4065_ ),
    .X(\u_cpu.ALU.u_wallace._4071_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9557_  (.A1(\u_cpu.ALU.u_wallace._3731_ ),
    .A2(\u_cpu.ALU.u_wallace._3737_ ),
    .B1(\u_cpu.ALU.u_wallace._3747_ ),
    .Y(\u_cpu.ALU.u_wallace._4072_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9558_  (.A(\u_cpu.ALU.u_wallace._0475_ ),
    .B(\u_cpu.ALU.u_wallace._3718_ ),
    .Y(\u_cpu.ALU.u_wallace._4074_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9559_  (.A(\u_cpu.ALU.u_wallace._3719_ ),
    .B(\u_cpu.ALU.u_wallace._2882_ ),
    .Y(\u_cpu.ALU.u_wallace._4075_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9560_  (.A1(\u_cpu.ALU.u_wallace._4074_ ),
    .A2(\u_cpu.ALU.u_wallace._4075_ ),
    .B1(\u_cpu.ALU.u_wallace._3721_ ),
    .Y(\u_cpu.ALU.u_wallace._4076_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9561_  (.A1(\u_cpu.ALU.u_wallace._1578_ ),
    .A2(\u_cpu.ALU.u_wallace._3718_ ),
    .B1(\u_cpu.ALU.u_wallace._2569_ ),
    .B2(\u_cpu.ALU.u_wallace._3719_ ),
    .X(\u_cpu.ALU.u_wallace._4077_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9562_  (.A(\u_cpu.ALU.u_wallace._3719_ ),
    .B(\u_cpu.ALU.u_wallace._1578_ ),
    .C(\u_cpu.ALU.u_wallace._3718_ ),
    .D(\u_cpu.ALU.u_wallace._2569_ ),
    .Y(\u_cpu.ALU.u_wallace._4078_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9563_  (.A(\u_cpu.ALU.u_wallace._4077_ ),
    .B(\u_cpu.ALU.u_wallace._4078_ ),
    .C(\u_cpu.ALU.u_wallace._0097_ ),
    .D(\u_cpu.ALU.SrcA[30] ),
    .Y(\u_cpu.ALU.u_wallace._4079_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._9564_  (.A(\u_cpu.ALU.SrcA[30] ),
    .Y(\u_cpu.ALU.u_wallace._4080_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9565_  (.A1(\u_cpu.ALU.u_wallace._0319_ ),
    .A2(\u_cpu.ALU.u_wallace._3718_ ),
    .B1(\u_cpu.ALU.u_wallace._2222_ ),
    .B2(\u_cpu.ALU.u_wallace._3719_ ),
    .Y(\u_cpu.ALU.u_wallace._4081_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9566_  (.A(\u_cpu.ALU.u_wallace._2779_ ),
    .B(\u_cpu.ALU.u_wallace._0319_ ),
    .C(\u_cpu.ALU.u_wallace._0629_ ),
    .D(\u_cpu.ALU.u_wallace._2222_ ),
    .X(\u_cpu.ALU.u_wallace._4082_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9567_  (.A1(\u_cpu.ALU.u_wallace._4934_ ),
    .A2(\u_cpu.ALU.u_wallace._4080_ ),
    .B1(\u_cpu.ALU.u_wallace._4081_ ),
    .B2(\u_cpu.ALU.u_wallace._4082_ ),
    .Y(\u_cpu.ALU.u_wallace._4083_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9568_  (.A1(\u_cpu.ALU.u_wallace._3723_ ),
    .A2(\u_cpu.ALU.u_wallace._4076_ ),
    .B1(\u_cpu.ALU.u_wallace._4079_ ),
    .C1(\u_cpu.ALU.u_wallace._4083_ ),
    .X(\u_cpu.ALU.u_wallace._4085_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9569_  (.A1(\u_cpu.ALU.u_wallace._3721_ ),
    .A2(\u_cpu.ALU.u_wallace._3720_ ),
    .B1(\u_cpu.ALU.u_wallace._3725_ ),
    .Y(\u_cpu.ALU.u_wallace._4086_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9570_  (.A1(\u_cpu.ALU.u_wallace._4079_ ),
    .A2(\u_cpu.ALU.u_wallace._4083_ ),
    .B1(\u_cpu.ALU.u_wallace._4086_ ),
    .Y(\u_cpu.ALU.u_wallace._4087_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9571_  (.A1(\u_cpu.ALU.u_wallace._0315_ ),
    .A2(\u_cpu.ALU.u_wallace._3399_ ),
    .B1(\u_cpu.ALU.SrcA[29] ),
    .B2(\u_cpu.ALU.u_wallace._0217_ ),
    .X(\u_cpu.ALU.u_wallace._4088_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9572_  (.A(\u_cpu.ALU.u_wallace._0228_ ),
    .B(\u_cpu.ALU.u_wallace._0315_ ),
    .C(\u_cpu.ALU.u_wallace._3399_ ),
    .D(\u_cpu.ALU.SrcA[29] ),
    .Y(\u_cpu.ALU.u_wallace._4089_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9573_  (.A(\u_cpu.ALU.u_wallace._4088_ ),
    .B(\u_cpu.ALU.u_wallace._3058_ ),
    .C(\u_cpu.ALU.u_wallace._4663_ ),
    .D(\u_cpu.ALU.u_wallace._4089_ ),
    .Y(\u_cpu.ALU.u_wallace._4090_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._9574_  (.A1_N(\u_cpu.ALU.u_wallace._4089_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4088_ ),
    .B1(\u_cpu.ALU.u_wallace._4678_ ),
    .B2(\u_cpu.ALU.u_wallace._3060_ ),
    .Y(\u_cpu.ALU.u_wallace._4091_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9575_  (.A(\u_cpu.ALU.u_wallace._4090_ ),
    .B(\u_cpu.ALU.u_wallace._4091_ ),
    .Y(\u_cpu.ALU.u_wallace._4092_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._9576_  (.A1(\u_cpu.ALU.u_wallace._4085_ ),
    .A2(\u_cpu.ALU.u_wallace._4087_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4092_ ),
    .Y(\u_cpu.ALU.u_wallace._4093_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9577_  (.A1(\u_cpu.ALU.u_wallace._3723_ ),
    .A2(\u_cpu.ALU.u_wallace._4076_ ),
    .B1(\u_cpu.ALU.u_wallace._4083_ ),
    .Y(\u_cpu.ALU.u_wallace._4094_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9578_  (.A(\u_cpu.ALU.u_wallace._4077_ ),
    .B(\u_cpu.ALU.u_wallace._4078_ ),
    .C(\u_cpu.ALU.u_wallace._0097_ ),
    .D(\u_cpu.ALU.SrcA[30] ),
    .X(\u_cpu.ALU.u_wallace._4096_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9579_  (.A1(\u_cpu.ALU.u_wallace._4079_ ),
    .A2(\u_cpu.ALU.u_wallace._4083_ ),
    .B1(\u_cpu.ALU.u_wallace._4086_ ),
    .X(\u_cpu.ALU.u_wallace._4097_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9580_  (.A1(\u_cpu.ALU.u_wallace._4094_ ),
    .A2(\u_cpu.ALU.u_wallace._4096_ ),
    .B1(\u_cpu.ALU.u_wallace._4092_ ),
    .C1(\u_cpu.ALU.u_wallace._4097_ ),
    .Y(\u_cpu.ALU.u_wallace._4098_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9581_  (.A(\u_cpu.ALU.u_wallace._4072_ ),
    .B(\u_cpu.ALU.u_wallace._4093_ ),
    .C(\u_cpu.ALU.u_wallace._4098_ ),
    .Y(\u_cpu.ALU.u_wallace._4099_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._9582_  (.A(\u_cpu.ALU.u_wallace._2869_ ),
    .X(\u_cpu.ALU.u_wallace._4100_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9583_  (.A1(\u_cpu.ALU.u_wallace._4663_ ),
    .A2(\u_cpu.ALU.u_wallace._4100_ ),
    .B1(\u_cpu.ALU.u_wallace._3732_ ),
    .B2(\u_cpu.ALU.u_wallace._3734_ ),
    .X(\u_cpu.ALU.u_wallace._4101_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9584_  (.A(\u_cpu.ALU.u_wallace._3732_ ),
    .B(\u_cpu.ALU.u_wallace._3734_ ),
    .C(\u_cpu.ALU.u_wallace._4663_ ),
    .D(\u_cpu.ALU.u_wallace._4100_ ),
    .Y(\u_cpu.ALU.u_wallace._4102_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9585_  (.A(\u_cpu.ALU.u_wallace._4101_ ),
    .B(\u_cpu.ALU.u_wallace._4102_ ),
    .Y(\u_cpu.ALU.u_wallace._4103_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9586_  (.A1(\u_cpu.ALU.u_wallace._4103_ ),
    .A2(\u_cpu.ALU.u_wallace._3748_ ),
    .B1(\u_cpu.ALU.u_wallace._3745_ ),
    .Y(\u_cpu.ALU.u_wallace._4104_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._9587_  (.A1(\u_cpu.ALU.u_wallace._4094_ ),
    .A2(\u_cpu.ALU.u_wallace._4096_ ),
    .B1(\u_cpu.ALU.u_wallace._4091_ ),
    .C1(\u_cpu.ALU.u_wallace._4090_ ),
    .D1(\u_cpu.ALU.u_wallace._4097_ ),
    .Y(\u_cpu.ALU.u_wallace._4105_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._9588_  (.A1_N(\u_cpu.ALU.u_wallace._4090_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4091_ ),
    .B1(\u_cpu.ALU.u_wallace._4085_ ),
    .B2(\u_cpu.ALU.u_wallace._4087_ ),
    .Y(\u_cpu.ALU.u_wallace._4107_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9589_  (.A(\u_cpu.ALU.u_wallace._4104_ ),
    .B(\u_cpu.ALU.u_wallace._4105_ ),
    .C(\u_cpu.ALU.u_wallace._4107_ ),
    .Y(\u_cpu.ALU.u_wallace._4108_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9590_  (.A(\u_cpu.ALU.u_wallace._0228_ ),
    .B(\u_cpu.ALU.u_wallace._0315_ ),
    .C(\u_cpu.ALU.u_wallace._3058_ ),
    .D(\u_cpu.ALU.u_wallace._3399_ ),
    .X(\u_cpu.ALU.u_wallace._4109_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._9591_  (.A1(\u_cpu.ALU.u_wallace._3732_ ),
    .A2(\u_cpu.ALU.u_wallace._4100_ ),
    .A3(\u_cpu.ALU.u_wallace._4663_ ),
    .B1(\u_cpu.ALU.u_wallace._4109_ ),
    .X(\u_cpu.ALU.u_wallace._4110_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9592_  (.A1(\u_cpu.ALU.u_wallace._2198_ ),
    .A2(\u_cpu.ALU.u_wallace._3449_ ),
    .B1(\u_cpu.ALU.u_wallace._4100_ ),
    .B2(\u_cpu.ALU.u_wallace._2166_ ),
    .X(\u_cpu.ALU.u_wallace._4111_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9593_  (.A(\u_cpu.ALU.u_wallace._2166_ ),
    .B(\u_cpu.ALU.u_wallace._2198_ ),
    .C(\u_cpu.ALU.u_wallace._3449_ ),
    .D(\u_cpu.ALU.u_wallace._4100_ ),
    .Y(\u_cpu.ALU.u_wallace._4112_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9594_  (.A(\u_cpu.ALU.u_wallace._4111_ ),
    .B(\u_cpu.ALU.u_wallace._2882_ ),
    .C(\u_cpu.ALU.u_wallace._2917_ ),
    .D(\u_cpu.ALU.u_wallace._4112_ ),
    .Y(\u_cpu.ALU.u_wallace._4113_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9595_  (.A(\u_cpu.ALU.u_wallace._2166_ ),
    .B(\u_cpu.ALU.u_wallace._2198_ ),
    .C(\u_cpu.ALU.u_wallace._3449_ ),
    .D(\u_cpu.ALU.u_wallace._2869_ ),
    .X(\u_cpu.ALU.u_wallace._4114_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9596_  (.A1(\u_cpu.ALU.u_wallace._2198_ ),
    .A2(\u_cpu.ALU.u_wallace._3449_ ),
    .B1(\u_cpu.ALU.u_wallace._4100_ ),
    .B2(\u_cpu.ALU.u_wallace._2166_ ),
    .Y(\u_cpu.ALU.u_wallace._4115_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9597_  (.A1(\u_cpu.ALU.u_wallace._2284_ ),
    .A2(\u_cpu.ALU.u_wallace._1987_ ),
    .B1(\u_cpu.ALU.u_wallace._4114_ ),
    .B2(\u_cpu.ALU.u_wallace._4115_ ),
    .Y(\u_cpu.ALU.u_wallace._4116_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9598_  (.A(\u_cpu.ALU.u_wallace._4110_ ),
    .B(\u_cpu.ALU.u_wallace._4113_ ),
    .C(\u_cpu.ALU.u_wallace._4116_ ),
    .Y(\u_cpu.ALU.u_wallace._4118_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9599_  (.A(\u_cpu.ALU.u_wallace._4113_ ),
    .B(\u_cpu.ALU.u_wallace._4116_ ),
    .Y(\u_cpu.ALU.u_wallace._4119_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._9600_  (.A1(\u_cpu.ALU.u_wallace._3732_ ),
    .A2(\u_cpu.ALU.u_wallace._4100_ ),
    .A3(\u_cpu.ALU.u_wallace._4663_ ),
    .B1(\u_cpu.ALU.u_wallace._4109_ ),
    .Y(\u_cpu.ALU.u_wallace._4120_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._9601_  (.A1(\u_cpu.ALU.u_wallace._3765_ ),
    .A2(\u_cpu.ALU.u_wallace._2598_ ),
    .A3(\u_cpu.ALU.u_wallace._2917_ ),
    .B1(\u_cpu.ALU.u_wallace._3763_ ),
    .X(\u_cpu.ALU.u_wallace._4121_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._9602_  (.A1(\u_cpu.ALU.u_wallace._4119_ ),
    .A2(\u_cpu.ALU.u_wallace._4120_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4121_ ),
    .Y(\u_cpu.ALU.u_wallace._4122_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9603_  (.A(\u_cpu.ALU.u_wallace._2917_ ),
    .B(\u_cpu.ALU.u_wallace._2882_ ),
    .Y(\u_cpu.ALU.u_wallace._4123_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._9604_  (.A(\u_cpu.ALU.u_wallace._4115_ ),
    .B(\u_cpu.ALU.u_wallace._4123_ ),
    .C(\u_cpu.ALU.u_wallace._4114_ ),
    .Y(\u_cpu.ALU.u_wallace._4124_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._9605_  (.A1(\u_cpu.ALU.u_wallace._2284_ ),
    .A2(\u_cpu.ALU.u_wallace._1987_ ),
    .B1(\u_cpu.ALU.u_wallace._4114_ ),
    .B2(\u_cpu.ALU.u_wallace._4115_ ),
    .X(\u_cpu.ALU.u_wallace._4125_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9606_  (.A1(\u_cpu.ALU.u_wallace._4124_ ),
    .A2(\u_cpu.ALU.u_wallace._4125_ ),
    .B1(\u_cpu.ALU.u_wallace._4120_ ),
    .Y(\u_cpu.ALU.u_wallace._4126_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9607_  (.A(\u_cpu.ALU.u_wallace._4118_ ),
    .B(\u_cpu.ALU.u_wallace._4126_ ),
    .Y(\u_cpu.ALU.u_wallace._4127_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._9608_  (.A(\u_cpu.ALU.u_wallace._4121_ ),
    .Y(\u_cpu.ALU.u_wallace._4129_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9609_  (.A1(\u_cpu.ALU.u_wallace._4118_ ),
    .A2(\u_cpu.ALU.u_wallace._4122_ ),
    .B1(\u_cpu.ALU.u_wallace._4127_ ),
    .B2(\u_cpu.ALU.u_wallace._4129_ ),
    .Y(\u_cpu.ALU.u_wallace._4130_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9610_  (.A1(\u_cpu.ALU.u_wallace._4099_ ),
    .A2(\u_cpu.ALU.u_wallace._4108_ ),
    .B1(\u_cpu.ALU.u_wallace._4130_ ),
    .Y(\u_cpu.ALU.u_wallace._4131_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._9611_  (.A(\u_cpu.ALU.u_wallace._4118_ ),
    .B(\u_cpu.ALU.u_wallace._4126_ ),
    .X(\u_cpu.ALU.u_wallace._4132_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9612_  (.A1(\u_cpu.ALU.u_wallace._4120_ ),
    .A2(\u_cpu.ALU.u_wallace._4119_ ),
    .B1(\u_cpu.ALU.u_wallace._4122_ ),
    .Y(\u_cpu.ALU.u_wallace._4133_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.ALU.u_wallace._9613_  (.A1(\u_cpu.ALU.u_wallace._4121_ ),
    .A2(\u_cpu.ALU.u_wallace._4132_ ),
    .B1(\u_cpu.ALU.u_wallace._4133_ ),
    .C1(\u_cpu.ALU.u_wallace._4099_ ),
    .D1(\u_cpu.ALU.u_wallace._4108_ ),
    .X(\u_cpu.ALU.u_wallace._4134_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._9614_  (.A1_N(\u_cpu.ALU.u_wallace._3781_ ),
    .A2_N(\u_cpu.ALU.u_wallace._3760_ ),
    .B1(\u_cpu.ALU.u_wallace._3794_ ),
    .B2(\u_cpu.ALU.u_wallace._3795_ ),
    .Y(\u_cpu.ALU.u_wallace._4135_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._9615_  (.A1(\u_cpu.ALU.u_wallace._4131_ ),
    .A2(\u_cpu.ALU.u_wallace._4134_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4135_ ),
    .Y(\u_cpu.ALU.u_wallace._4136_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9616_  (.A(\u_cpu.ALU.u_wallace._3779_ ),
    .B(\u_cpu.ALU.u_wallace._3778_ ),
    .Y(\u_cpu.ALU.u_wallace._4137_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9617_  (.A1(\u_cpu.ALU.u_wallace._3772_ ),
    .A2(\u_cpu.ALU.u_wallace._4042_ ),
    .B1(\u_cpu.ALU.u_wallace._3770_ ),
    .Y(\u_cpu.ALU.u_wallace._4138_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9618_  (.A1(\u_cpu.ALU.u_wallace._4042_ ),
    .A2(\u_cpu.ALU.u_wallace._4137_ ),
    .B1(\u_cpu.ALU.u_wallace._4138_ ),
    .Y(\u_cpu.ALU.u_wallace._4140_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._9619_  (.A1(\u_cpu.ALU.u_wallace._3759_ ),
    .A2(\u_cpu.ALU.u_wallace._3751_ ),
    .A3(\u_cpu.ALU.u_wallace._3752_ ),
    .B1(\u_cpu.ALU.u_wallace._4140_ ),
    .Y(\u_cpu.ALU.u_wallace._4141_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9620_  (.A(\u_cpu.ALU.u_wallace._4121_ ),
    .B(\u_cpu.ALU.u_wallace._4118_ ),
    .C(\u_cpu.ALU.u_wallace._4126_ ),
    .X(\u_cpu.ALU.u_wallace._4142_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU.u_wallace._9621_  (.A1(\u_cpu.ALU.u_wallace._2284_ ),
    .A2(\u_cpu.ALU.u_wallace._1737_ ),
    .A3(\u_cpu.ALU.u_wallace._3762_ ),
    .B1(\u_cpu.ALU.u_wallace._3767_ ),
    .C1(\u_cpu.ALU.u_wallace._4127_ ),
    .X(\u_cpu.ALU.u_wallace._4143_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._9622_  (.A1_N(\u_cpu.ALU.u_wallace._4099_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4108_ ),
    .B1(\u_cpu.ALU.u_wallace._4142_ ),
    .B2(\u_cpu.ALU.u_wallace._4143_ ),
    .Y(\u_cpu.ALU.u_wallace._4144_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9623_  (.A1(\u_cpu.ALU.u_wallace._4118_ ),
    .A2(\u_cpu.ALU.u_wallace._4126_ ),
    .B1(\u_cpu.ALU.u_wallace._4121_ ),
    .X(\u_cpu.ALU.u_wallace._4145_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9624_  (.A(\u_cpu.ALU.u_wallace._4099_ ),
    .B(\u_cpu.ALU.u_wallace._4108_ ),
    .C(\u_cpu.ALU.u_wallace._4133_ ),
    .D(\u_cpu.ALU.u_wallace._4145_ ),
    .Y(\u_cpu.ALU.u_wallace._4146_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9625_  (.A1(\u_cpu.ALU.u_wallace._3750_ ),
    .A2(\u_cpu.ALU.u_wallace._4141_ ),
    .B1(\u_cpu.ALU.u_wallace._4144_ ),
    .C1(\u_cpu.ALU.u_wallace._4146_ ),
    .Y(\u_cpu.ALU.u_wallace._4147_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.ALU.u_wallace._9626_  (.A1(\u_cpu.ALU.u_wallace._4064_ ),
    .A2(\u_cpu.ALU.u_wallace._4070_ ),
    .B1(\u_cpu.ALU.u_wallace._4071_ ),
    .C1(\u_cpu.ALU.u_wallace._4136_ ),
    .D1(\u_cpu.ALU.u_wallace._4147_ ),
    .Y(\u_cpu.ALU.u_wallace._4148_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9627_  (.A(\u_cpu.ALU.u_wallace._4065_ ),
    .B(\u_cpu.ALU.u_wallace._4063_ ),
    .C(\u_cpu.ALU.u_wallace._4069_ ),
    .X(\u_cpu.ALU.u_wallace._4149_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9628_  (.A1(\u_cpu.ALU.u_wallace._4063_ ),
    .A2(\u_cpu.ALU.u_wallace._4069_ ),
    .B1(\u_cpu.ALU.u_wallace._4065_ ),
    .Y(\u_cpu.ALU.u_wallace._4151_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9629_  (.A1(\u_cpu.ALU.u_wallace._4144_ ),
    .A2(\u_cpu.ALU.u_wallace._4146_ ),
    .B1(\u_cpu.ALU.u_wallace._4135_ ),
    .Y(\u_cpu.ALU.u_wallace._4152_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9630_  (.A1(\u_cpu.ALU.u_wallace._3750_ ),
    .A2(\u_cpu.ALU.u_wallace._4141_ ),
    .B1(\u_cpu.ALU.u_wallace._4144_ ),
    .C1(\u_cpu.ALU.u_wallace._4146_ ),
    .X(\u_cpu.ALU.u_wallace._4153_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9631_  (.A1(\u_cpu.ALU.u_wallace._4149_ ),
    .A2(\u_cpu.ALU.u_wallace._4151_ ),
    .B1(\u_cpu.ALU.u_wallace._4152_ ),
    .B2(\u_cpu.ALU.u_wallace._4153_ ),
    .Y(\u_cpu.ALU.u_wallace._4154_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9632_  (.A1(\u_cpu.ALU.u_wallace._3808_ ),
    .A2(\u_cpu.ALU.u_wallace._3805_ ),
    .B1(\u_cpu.ALU.u_wallace._3793_ ),
    .Y(\u_cpu.ALU.u_wallace._4155_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9633_  (.A1(\u_cpu.ALU.u_wallace._4148_ ),
    .A2(\u_cpu.ALU.u_wallace._4154_ ),
    .B1(\u_cpu.ALU.u_wallace._4155_ ),
    .Y(\u_cpu.ALU.u_wallace._4156_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9634_  (.A1(\u_cpu.ALU.u_wallace._4064_ ),
    .A2(\u_cpu.ALU.u_wallace._4070_ ),
    .B1(\u_cpu.ALU.u_wallace._4071_ ),
    .C1(\u_cpu.ALU.u_wallace._4136_ ),
    .Y(\u_cpu.ALU.u_wallace._4157_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9635_  (.A1(\u_cpu.ALU.u_wallace._4153_ ),
    .A2(\u_cpu.ALU.u_wallace._4157_ ),
    .B1(\u_cpu.ALU.u_wallace._4154_ ),
    .C1(\u_cpu.ALU.u_wallace._4155_ ),
    .X(\u_cpu.ALU.u_wallace._4158_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9636_  (.A1(\u_cpu.ALU.u_wallace._4038_ ),
    .A2(\u_cpu.ALU.u_wallace._4041_ ),
    .B1(\u_cpu.ALU.u_wallace._4156_ ),
    .B2(\u_cpu.ALU.u_wallace._4158_ ),
    .Y(\u_cpu.ALU.u_wallace._4159_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9637_  (.A1(\u_cpu.ALU.u_wallace._4148_ ),
    .A2(\u_cpu.ALU.u_wallace._4154_ ),
    .B1(\u_cpu.ALU.u_wallace._4155_ ),
    .X(\u_cpu.ALU.u_wallace._4160_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9638_  (.A1(\u_cpu.ALU.u_wallace._4153_ ),
    .A2(\u_cpu.ALU.u_wallace._4157_ ),
    .B1(\u_cpu.ALU.u_wallace._4154_ ),
    .C1(\u_cpu.ALU.u_wallace._4155_ ),
    .Y(\u_cpu.ALU.u_wallace._4162_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9639_  (.A1(\u_cpu.ALU.u_wallace._4034_ ),
    .A2(\u_cpu.ALU.u_wallace._4035_ ),
    .B1(\u_cpu.ALU.u_wallace._4031_ ),
    .Y(\u_cpu.ALU.u_wallace._4163_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9640_  (.A(\u_cpu.ALU.u_wallace._4037_ ),
    .B(\u_cpu.ALU.u_wallace._4163_ ),
    .Y(\u_cpu.ALU.u_wallace._4164_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9641_  (.A1(\u_cpu.ALU.u_wallace._4164_ ),
    .A2(\u_cpu.ALU.u_wallace._4036_ ),
    .B1(\u_cpu.ALU.u_wallace._4038_ ),
    .Y(\u_cpu.ALU.u_wallace._4165_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9642_  (.A(\u_cpu.ALU.u_wallace._4160_ ),
    .B(\u_cpu.ALU.u_wallace._4162_ ),
    .C(\u_cpu.ALU.u_wallace._4165_ ),
    .Y(\u_cpu.ALU.u_wallace._4166_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9643_  (.A1(\u_cpu.ALU.u_wallace._3800_ ),
    .A2(\u_cpu.ALU.u_wallace._3806_ ),
    .B1(\u_cpu.ALU.u_wallace._3680_ ),
    .Y(\u_cpu.ALU.u_wallace._4167_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9644_  (.A1(\u_cpu.ALU.u_wallace._3817_ ),
    .A2(\u_cpu.ALU.u_wallace._4167_ ),
    .B1(\u_cpu.ALU.u_wallace._3807_ ),
    .Y(\u_cpu.ALU.u_wallace._4168_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9645_  (.A1(\u_cpu.ALU.u_wallace._4159_ ),
    .A2(\u_cpu.ALU.u_wallace._4166_ ),
    .B1(\u_cpu.ALU.u_wallace._4168_ ),
    .Y(\u_cpu.ALU.u_wallace._4169_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9646_  (.A1(\u_cpu.ALU.u_wallace._3660_ ),
    .A2(\u_cpu.ALU.u_wallace._4039_ ),
    .B1(\u_cpu.ALU.u_wallace._4032_ ),
    .Y(\u_cpu.ALU.u_wallace._4170_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._9647_  (.A(\u_cpu.ALU.u_wallace._4036_ ),
    .Y(\u_cpu.ALU.u_wallace._4171_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._9648_  (.A1(\u_cpu.ALU.u_wallace._4032_ ),
    .A2(\u_cpu.ALU.u_wallace._4036_ ),
    .B1(\u_cpu.ALU.u_wallace._3660_ ),
    .C1(\u_cpu.ALU.u_wallace._4039_ ),
    .X(\u_cpu.ALU.u_wallace._4173_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9649_  (.A1(\u_cpu.ALU.u_wallace._4170_ ),
    .A2(\u_cpu.ALU.u_wallace._4171_ ),
    .B1(\u_cpu.ALU.u_wallace._4173_ ),
    .C1(\u_cpu.ALU.u_wallace._4162_ ),
    .Y(\u_cpu.ALU.u_wallace._4174_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9650_  (.A(\u_cpu.ALU.u_wallace._3680_ ),
    .B(\u_cpu.ALU.u_wallace._3800_ ),
    .C(\u_cpu.ALU.u_wallace._3806_ ),
    .X(\u_cpu.ALU.u_wallace._4175_ ));
 sky130_fd_sc_hd__a311oi_2 \u_cpu.ALU.u_wallace._9651_  (.A1(\u_cpu.ALU.u_wallace._3809_ ),
    .A2(\u_cpu.ALU.u_wallace._3811_ ),
    .A3(\u_cpu.ALU.u_wallace._3812_ ),
    .B1(\u_cpu.ALU.u_wallace._3819_ ),
    .C1(\u_cpu.ALU.u_wallace._3820_ ),
    .Y(\u_cpu.ALU.u_wallace._4176_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._9652_  (.A1(\u_cpu.ALU.u_wallace._4156_ ),
    .A2(\u_cpu.ALU.u_wallace._4174_ ),
    .B1(\u_cpu.ALU.u_wallace._4175_ ),
    .B2(\u_cpu.ALU.u_wallace._4176_ ),
    .C1(\u_cpu.ALU.u_wallace._4159_ ),
    .X(\u_cpu.ALU.u_wallace._4177_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9653_  (.A1(\u_cpu.ALU.u_wallace._3980_ ),
    .A2(\u_cpu.ALU.u_wallace._3981_ ),
    .B1(\u_cpu.ALU.u_wallace._4169_ ),
    .B2(\u_cpu.ALU.u_wallace._4177_ ),
    .Y(\u_cpu.ALU.u_wallace._4178_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9654_  (.A1(\u_cpu.ALU.u_wallace._4159_ ),
    .A2(\u_cpu.ALU.u_wallace._4166_ ),
    .B1(\u_cpu.ALU.u_wallace._4168_ ),
    .X(\u_cpu.ALU.u_wallace._4179_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._9655_  (.A1(\u_cpu.ALU.u_wallace._4156_ ),
    .A2(\u_cpu.ALU.u_wallace._4174_ ),
    .B1(\u_cpu.ALU.u_wallace._4175_ ),
    .B2(\u_cpu.ALU.u_wallace._4176_ ),
    .C1(\u_cpu.ALU.u_wallace._4159_ ),
    .Y(\u_cpu.ALU.u_wallace._4180_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._9656_  (.A1(\u_cpu.ALU.u_wallace._3874_ ),
    .A2(\u_cpu.ALU.u_wallace._3978_ ),
    .B1(\u_cpu.ALU.u_wallace._3977_ ),
    .X(\u_cpu.ALU.u_wallace._4181_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9657_  (.A1(\u_cpu.ALU.u_wallace._4181_ ),
    .A2(\u_cpu.ALU.u_wallace._3972_ ),
    .B1(\u_cpu.ALU.u_wallace._3980_ ),
    .Y(\u_cpu.ALU.u_wallace._4182_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9658_  (.A(\u_cpu.ALU.u_wallace._4179_ ),
    .B(\u_cpu.ALU.u_wallace._4180_ ),
    .C(\u_cpu.ALU.u_wallace._4182_ ),
    .Y(\u_cpu.ALU.u_wallace._4184_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9659_  (.A1(\u_cpu.ALU.u_wallace._3880_ ),
    .A2(\u_cpu.ALU.u_wallace._3827_ ),
    .B1(\u_cpu.ALU.u_wallace._3885_ ),
    .X(\u_cpu.ALU.u_wallace._4185_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9660_  (.A1(\u_cpu.ALU.u_wallace._4178_ ),
    .A2(\u_cpu.ALU.u_wallace._4184_ ),
    .B1(\u_cpu.ALU.u_wallace._4185_ ),
    .X(\u_cpu.ALU.u_wallace._4186_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9661_  (.A(\u_cpu.ALU.u_wallace._4185_ ),
    .B(\u_cpu.ALU.u_wallace._4178_ ),
    .C(\u_cpu.ALU.u_wallace._4184_ ),
    .Y(\u_cpu.ALU.u_wallace._4187_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.ALU.u_wallace._9662_  (.A1(\u_cpu.ALU.u_wallace._3830_ ),
    .A2(\u_cpu.ALU.u_wallace._3867_ ),
    .A3(\u_cpu.ALU.u_wallace._3868_ ),
    .B1(\u_cpu.ALU.u_wallace._3875_ ),
    .B2(\u_cpu.ALU.u_wallace._3877_ ),
    .X(\u_cpu.ALU.u_wallace._4188_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9663_  (.A1(\u_cpu.ALU.u_wallace._4186_ ),
    .A2(\u_cpu.ALU.u_wallace._4187_ ),
    .B1(\u_cpu.ALU.u_wallace._4188_ ),
    .Y(\u_cpu.ALU.u_wallace._4189_ ));
 sky130_fd_sc_hd__a32oi_2 \u_cpu.ALU.u_wallace._9664_  (.A1(\u_cpu.ALU.u_wallace._3830_ ),
    .A2(\u_cpu.ALU.u_wallace._3867_ ),
    .A3(\u_cpu.ALU.u_wallace._3868_ ),
    .B1(\u_cpu.ALU.u_wallace._3875_ ),
    .B2(\u_cpu.ALU.u_wallace._3877_ ),
    .Y(\u_cpu.ALU.u_wallace._4190_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9665_  (.A1(\u_cpu.ALU.u_wallace._4178_ ),
    .A2(\u_cpu.ALU.u_wallace._4184_ ),
    .B1(\u_cpu.ALU.u_wallace._4185_ ),
    .Y(\u_cpu.ALU.u_wallace._4191_ ));
 sky130_fd_sc_hd__nor3b_2 \u_cpu.ALU.u_wallace._9666_  (.A(\u_cpu.ALU.u_wallace._4190_ ),
    .B(\u_cpu.ALU.u_wallace._4191_ ),
    .C_N(\u_cpu.ALU.u_wallace._4187_ ),
    .Y(\u_cpu.ALU.u_wallace._4192_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9667_  (.A1(\u_cpu.ALU.u_wallace._4189_ ),
    .A2(\u_cpu.ALU.u_wallace._4192_ ),
    .B1(\u_cpu.ALU.u_wallace._3889_ ),
    .C1(\u_cpu.ALU.u_wallace._3892_ ),
    .Y(\u_cpu.ALU.u_wallace._4193_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._9668_  (.A1(\u_cpu.ALU.u_wallace._3889_ ),
    .A2(\u_cpu.ALU.u_wallace._3892_ ),
    .B1(\u_cpu.ALU.u_wallace._4189_ ),
    .C1(\u_cpu.ALU.u_wallace._4192_ ),
    .X(\u_cpu.ALU.u_wallace._4195_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9669_  (.A(\u_cpu.ALU.u_wallace._4193_ ),
    .B(\u_cpu.ALU.u_wallace._4195_ ),
    .Y(\u_cpu.ALU.u_wallace._4196_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._9670_  (.A(\u_cpu.ALU.u_wallace._3910_ ),
    .B(\u_cpu.ALU.u_wallace._4196_ ),
    .X(\u_cpu.ALU.u_wallace._4197_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._9671_  (.A(\u_cpu.ALU.u_wallace._3909_ ),
    .B(\u_cpu.ALU.u_wallace._4197_ ),
    .X(\u_cpu.ALU.u_wallace._4198_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._9672_  (.A1(\u_cpu.ALU.u_wallace._3905_ ),
    .A2(\u_cpu.ALU.u_wallace._3907_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4198_ ),
    .Y(\u_cpu.ALU.u_wallace._4199_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9673_  (.A1(\u_cpu.ALU.u_wallace._3335_ ),
    .A2(\u_cpu.ALU.u_wallace._3607_ ),
    .B1(\u_cpu.ALU.u_wallace._3901_ ),
    .Y(\u_cpu.ALU.u_wallace._4200_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9674_  (.A(\u_cpu.ALU.u_wallace._3608_ ),
    .B(\u_cpu.ALU.u_wallace._3900_ ),
    .C(\u_cpu.ALU.u_wallace._3901_ ),
    .X(\u_cpu.ALU.u_wallace._4201_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9675_  (.A1(\u_cpu.ALU.u_wallace._3900_ ),
    .A2(\u_cpu.ALU.u_wallace._4200_ ),
    .B1(\u_cpu.ALU.u_wallace._4201_ ),
    .B2(\u_cpu.ALU.u_wallace._3614_ ),
    .Y(\u_cpu.ALU.u_wallace._4202_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9676_  (.A(\u_cpu.ALU.u_wallace._4202_ ),
    .B(\u_cpu.ALU.u_wallace._4198_ ),
    .Y(\u_cpu.ALU.u_wallace._4203_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._9677_  (.A(\u_cpu.ALU.u_wallace._4199_ ),
    .B(\u_cpu.ALU.u_wallace._4203_ ),
    .X(\u_cpu.ALU.u_wallace._4204_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._9678_  (.A(\u_cpu.ALU.u_wallace._4204_ ),
    .X(\u_cpu.ALU.Product_Wallace[30] ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9679_  (.A(\u_cpu.ALU.u_wallace._4198_ ),
    .B(\u_cpu.ALU.u_wallace._4202_ ),
    .Y(\u_cpu.ALU.u_wallace._4206_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.ALU.u_wallace._9680_  (.A(\u_cpu.ALU.u_wallace._3909_ ),
    .B_N(\u_cpu.ALU.u_wallace._4197_ ),
    .X(\u_cpu.ALU.u_wallace._4207_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._9681_  (.A1(\u_cpu.ALU.u_wallace._3912_ ),
    .A2(\u_cpu.ALU.u_wallace._2480_ ),
    .A3(\u_cpu.ALU.u_wallace._1333_ ),
    .B1(\u_cpu.ALU.u_wallace._3916_ ),
    .X(\u_cpu.ALU.u_wallace._4208_ ));
 sky130_fd_sc_hd__a21bo_2 \u_cpu.ALU.u_wallace._9682_  (.A1(\u_cpu.ALU.u_wallace._3858_ ),
    .A2(\u_cpu.ALU.u_wallace._3950_ ),
    .B1_N(\u_cpu.ALU.u_wallace._3957_ ),
    .X(\u_cpu.ALU.u_wallace._4209_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu.ALU.u_wallace._9683_  (.A(\u_cpu.ALU.u_wallace._3983_ ),
    .B(\u_cpu.ALU.u_wallace._4209_ ),
    .Y(\u_cpu.ALU.u_wallace._4210_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9684_  (.A(\u_cpu.ALU.u_wallace._0370_ ),
    .B(\u_cpu.ALU.SrcB[29] ),
    .Y(\u_cpu.ALU.u_wallace._4211_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._9685_  (.A1(\u_cpu.ALU.u_wallace._3982_ ),
    .A2(\u_cpu.ALU.u_wallace._3983_ ),
    .A3(\u_cpu.ALU.u_wallace._3991_ ),
    .B1(\u_cpu.ALU.u_wallace._3994_ ),
    .X(\u_cpu.ALU.u_wallace._4212_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu.ALU.u_wallace._9686_  (.A(\u_cpu.ALU.u_wallace._4211_ ),
    .B(\u_cpu.ALU.u_wallace._4212_ ),
    .Y(\u_cpu.ALU.u_wallace._4213_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9687_  (.A1(\u_cpu.ALU.u_wallace._0184_ ),
    .A2(\u_cpu.ALU.SrcB[30] ),
    .B1(\u_cpu.ALU.u_wallace._3934_ ),
    .Y(\u_cpu.ALU.u_wallace._4214_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9688_  (.A(\u_cpu.ALU.u_wallace._3934_ ),
    .B(\u_cpu.ALU.SrcB[30] ),
    .C(\u_cpu.ALU.u_wallace._0184_ ),
    .D(\u_cpu.ALU.u_wallace._3944_ ),
    .X(\u_cpu.ALU.u_wallace._4216_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU.u_wallace._9689_  (.A1(\u_cpu.ALU.u_wallace._3942_ ),
    .A2(\u_cpu.ALU.u_wallace._3955_ ),
    .B1(\u_cpu.ALU.u_wallace._0621_ ),
    .C1(\u_cpu.ALU.u_wallace._3549_ ),
    .Y(\u_cpu.ALU.u_wallace._4217_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9690_  (.A1(\u_cpu.ALU.u_wallace._0621_ ),
    .A2(\u_cpu.ALU.u_wallace._3549_ ),
    .B1(\u_cpu.ALU.u_wallace._3942_ ),
    .C1(\u_cpu.ALU.u_wallace._3955_ ),
    .X(\u_cpu.ALU.u_wallace._4218_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9691_  (.A(\u_cpu.ALU.u_wallace._4217_ ),
    .B(\u_cpu.ALU.u_wallace._4218_ ),
    .Y(\u_cpu.ALU.u_wallace._4219_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.ALU.u_wallace._9692_  (.A(\u_cpu.ALU.u_wallace._4214_ ),
    .B(\u_cpu.ALU.u_wallace._4216_ ),
    .C(\u_cpu.ALU.u_wallace._4219_ ),
    .Y(\u_cpu.ALU.u_wallace._4220_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._9693_  (.A1(\u_cpu.ALU.u_wallace._4214_ ),
    .A2(\u_cpu.ALU.u_wallace._4216_ ),
    .B1(\u_cpu.ALU.u_wallace._4219_ ),
    .X(\u_cpu.ALU.u_wallace._4221_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU.u_wallace._9694_  (.A(\u_cpu.ALU.u_wallace._4220_ ),
    .B(\u_cpu.ALU.u_wallace._4221_ ),
    .X(\u_cpu.ALU.u_wallace._4222_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu.ALU.u_wallace._9695_  (.A(\u_cpu.ALU.u_wallace._4213_ ),
    .B(\u_cpu.ALU.u_wallace._4222_ ),
    .Y(\u_cpu.ALU.u_wallace._4223_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu.ALU.u_wallace._9696_  (.A(\u_cpu.ALU.u_wallace._4210_ ),
    .B(\u_cpu.ALU.u_wallace._4223_ ),
    .Y(\u_cpu.ALU.u_wallace._4224_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._9697_  (.A(\u_cpu.ALU.u_wallace._4208_ ),
    .B(\u_cpu.ALU.u_wallace._4224_ ),
    .X(\u_cpu.ALU.u_wallace._4225_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9698_  (.A1(\u_cpu.ALU.u_wallace._4180_ ),
    .A2(\u_cpu.ALU.u_wallace._4184_ ),
    .B1(\u_cpu.ALU.u_wallace._4225_ ),
    .Y(\u_cpu.ALU.u_wallace._4227_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU.u_wallace._9699_  (.A1(\u_cpu.ALU.u_wallace._3980_ ),
    .A2(\u_cpu.ALU.u_wallace._3981_ ),
    .A3(\u_cpu.ALU.u_wallace._4169_ ),
    .B1(\u_cpu.ALU.u_wallace._4180_ ),
    .C1(\u_cpu.ALU.u_wallace._4225_ ),
    .X(\u_cpu.ALU.u_wallace._4228_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9700_  (.A(\u_cpu.ALU.u_wallace._4227_ ),
    .B(\u_cpu.ALU.u_wallace._4228_ ),
    .Y(\u_cpu.ALU.u_wallace._4229_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9701_  (.A1(\u_cpu.ALU.u_wallace._3910_ ),
    .A2(\u_cpu.ALU.u_wallace._4196_ ),
    .B1(\u_cpu.ALU.u_wallace._4195_ ),
    .Y(\u_cpu.ALU.u_wallace._4230_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu.ALU.u_wallace._9702_  (.A(\u_cpu.ALU.u_wallace._4229_ ),
    .B(\u_cpu.ALU.u_wallace._4230_ ),
    .Y(\u_cpu.ALU.u_wallace._4231_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9703_  (.A1(\u_cpu.ALU.u_wallace._1333_ ),
    .A2(\u_cpu.ALU.u_wallace._3258_ ),
    .B1(\u_cpu.ALU.u_wallace._3923_ ),
    .B2(\u_cpu.ALU.u_wallace._3924_ ),
    .X(\u_cpu.ALU.u_wallace._4232_ ));
 sky130_fd_sc_hd__or4b_2 \u_cpu.ALU.u_wallace._9704_  (.A(\u_cpu.ALU.u_wallace._4813_ ),
    .B(\u_cpu.ALU.u_wallace._3263_ ),
    .C(\u_cpu.ALU.u_wallace._3921_ ),
    .D_N(\u_cpu.ALU.u_wallace._3924_ ),
    .X(\u_cpu.ALU.u_wallace._4233_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9705_  (.A(\u_cpu.ALU.u_wallace._4232_ ),
    .B(\u_cpu.ALU.u_wallace._4233_ ),
    .Y(\u_cpu.ALU.u_wallace._4234_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._9706_  (.A(\u_cpu.ALU.u_wallace._3962_ ),
    .Y(\u_cpu.ALU.u_wallace._4235_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9707_  (.A1(\u_cpu.ALU.u_wallace._3966_ ),
    .A2(\u_cpu.ALU.u_wallace._3970_ ),
    .B1(\u_cpu.ALU.u_wallace._4235_ ),
    .X(\u_cpu.ALU.u_wallace._4236_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._9708_  (.A(\u_cpu.ALU.u_wallace._4234_ ),
    .B(\u_cpu.ALU.u_wallace._4236_ ),
    .X(\u_cpu.ALU.u_wallace._4238_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._9709_  (.A1(\u_cpu.ALU.u_wallace._4185_ ),
    .A2(\u_cpu.ALU.u_wallace._4178_ ),
    .A3(\u_cpu.ALU.u_wallace._4184_ ),
    .B1(\u_cpu.ALU.u_wallace._4192_ ),
    .X(\u_cpu.ALU.u_wallace._4239_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._9710_  (.A(\u_cpu.ALU.u_wallace._4238_ ),
    .B(\u_cpu.ALU.u_wallace._4239_ ),
    .X(\u_cpu.ALU.u_wallace._4240_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9711_  (.A(\u_cpu.ALU.u_wallace._3925_ ),
    .B(\u_cpu.ALU.u_wallace._3922_ ),
    .C(\u_cpu.ALU.u_wallace._3924_ ),
    .X(\u_cpu.ALU.u_wallace._4241_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._9712_  (.A1(\u_cpu.ALU.u_wallace._3926_ ),
    .A2(\u_cpu.ALU.u_wallace._2417_ ),
    .A3(\u_cpu.ALU.u_wallace._2343_ ),
    .B1(\u_cpu.ALU.u_wallace._4241_ ),
    .X(\u_cpu.ALU.u_wallace._4242_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9713_  (.A1(\u_cpu.ALU.u_wallace._4661_ ),
    .A2(\u_cpu.ALU.u_wallace._2417_ ),
    .B1(\u_cpu.ALU.u_wallace._2480_ ),
    .B2(\u_cpu.ALU.u_wallace._0198_ ),
    .X(\u_cpu.ALU.u_wallace._4243_ ));
 sky130_fd_sc_hd__or4_2 \u_cpu.ALU.u_wallace._9714_  (.A(\u_cpu.ALU.u_wallace._4677_ ),
    .B(\u_cpu.ALU.u_wallace._4454_ ),
    .C(\u_cpu.ALU.u_wallace._2131_ ),
    .D(\u_cpu.ALU.u_wallace._2482_ ),
    .X(\u_cpu.ALU.u_wallace._4244_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9715_  (.A(\u_cpu.ALU.u_wallace._3253_ ),
    .B(\u_cpu.ALU.u_wallace._3254_ ),
    .Y(\u_cpu.ALU.u_wallace._4245_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9716_  (.A1(\u_cpu.ALU.u_wallace._2343_ ),
    .A2(\u_cpu.ALU.u_wallace._2402_ ),
    .B1(\u_cpu.ALU.u_wallace._4245_ ),
    .Y(\u_cpu.ALU.u_wallace._4246_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9717_  (.A(\u_cpu.ALU.u_wallace._4245_ ),
    .B(\u_cpu.ALU.u_wallace._2402_ ),
    .C(\u_cpu.ALU.u_wallace._2343_ ),
    .X(\u_cpu.ALU.u_wallace._4247_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._9718_  (.A1(\u_cpu.ALU.u_wallace._4037_ ),
    .A2(\u_cpu.ALU.u_wallace._4163_ ),
    .B1(\u_cpu.ALU.u_wallace._4036_ ),
    .X(\u_cpu.ALU.u_wallace._4248_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.ALU.u_wallace._9719_  (.A(\u_cpu.ALU.u_wallace._4246_ ),
    .B(\u_cpu.ALU.u_wallace._4247_ ),
    .C(\u_cpu.ALU.u_wallace._4248_ ),
    .X(\u_cpu.ALU.u_wallace._4249_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9720_  (.A1(\u_cpu.ALU.u_wallace._4246_ ),
    .A2(\u_cpu.ALU.u_wallace._4247_ ),
    .B1(\u_cpu.ALU.u_wallace._4248_ ),
    .Y(\u_cpu.ALU.u_wallace._4250_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9721_  (.A(\u_cpu.ALU.u_wallace._4249_ ),
    .B(\u_cpu.ALU.u_wallace._4250_ ),
    .Y(\u_cpu.ALU.u_wallace._4251_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9722_  (.A(\u_cpu.ALU.u_wallace._4243_ ),
    .B(\u_cpu.ALU.u_wallace._4244_ ),
    .C(\u_cpu.ALU.u_wallace._4251_ ),
    .X(\u_cpu.ALU.u_wallace._4252_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9723_  (.A1(\u_cpu.ALU.u_wallace._4243_ ),
    .A2(\u_cpu.ALU.u_wallace._4244_ ),
    .B1(\u_cpu.ALU.u_wallace._4251_ ),
    .Y(\u_cpu.ALU.u_wallace._4253_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU.u_wallace._9724_  (.A(\u_cpu.ALU.u_wallace._4252_ ),
    .B(\u_cpu.ALU.u_wallace._4253_ ),
    .X(\u_cpu.ALU.u_wallace._4254_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._9725_  (.A(\u_cpu.ALU.u_wallace._4242_ ),
    .B(\u_cpu.ALU.u_wallace._4254_ ),
    .X(\u_cpu.ALU.u_wallace._4255_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._9726_  (.A1(\u_cpu.ALU.u_wallace._4110_ ),
    .A2(\u_cpu.ALU.u_wallace._4113_ ),
    .A3(\u_cpu.ALU.u_wallace._4116_ ),
    .B1(\u_cpu.ALU.u_wallace._4122_ ),
    .X(\u_cpu.ALU.u_wallace._4256_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._9727_  (.A1(\u_cpu.ALU.u_wallace._4733_ ),
    .A2(\u_cpu.ALU.u_wallace._3088_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4256_ ),
    .Y(\u_cpu.ALU.u_wallace._4257_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.ALU.u_wallace._9728_  (.A_N(\u_cpu.ALU.u_wallace._4122_ ),
    .B(\u_cpu.ALU.u_wallace._3088_ ),
    .C(\u_cpu.ALU.u_wallace._4733_ ),
    .D(\u_cpu.ALU.u_wallace._4118_ ),
    .X(\u_cpu.ALU.u_wallace._4259_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9729_  (.A(\u_cpu.ALU.u_wallace._0228_ ),
    .B(\u_cpu.ALU.SrcA[30] ),
    .Y(\u_cpu.ALU.u_wallace._4260_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.ALU.u_wallace._9730_  (.A1(\u_cpu.ALU.u_wallace._0097_ ),
    .A2(\u_cpu.ALU.SrcA[30] ),
    .A3(\u_cpu.ALU.u_wallace._4077_ ),
    .A4(\u_cpu.ALU.u_wallace._4078_ ),
    .B1(\u_cpu.ALU.u_wallace._4094_ ),
    .X(\u_cpu.ALU.u_wallace._4261_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9731_  (.A1(\u_cpu.ALU.u_wallace._4092_ ),
    .A2(\u_cpu.ALU.u_wallace._4087_ ),
    .B1(\u_cpu.ALU.u_wallace._4260_ ),
    .C1(\u_cpu.ALU.u_wallace._4261_ ),
    .Y(\u_cpu.ALU.u_wallace._4262_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9732_  (.A1(\u_cpu.ALU.u_wallace._4096_ ),
    .A2(\u_cpu.ALU.u_wallace._4094_ ),
    .B1(\u_cpu.ALU.u_wallace._4092_ ),
    .B2(\u_cpu.ALU.u_wallace._4087_ ),
    .Y(\u_cpu.ALU.u_wallace._4263_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._9733_  (.A(\u_cpu.ALU.u_wallace._0228_ ),
    .B(\u_cpu.ALU.SrcA[30] ),
    .X(\u_cpu.ALU.u_wallace._4264_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9734_  (.A(\u_cpu.ALU.u_wallace._4263_ ),
    .B(\u_cpu.ALU.u_wallace._4264_ ),
    .Y(\u_cpu.ALU.u_wallace._4265_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9735_  (.A(\u_cpu.ALU.u_wallace._0228_ ),
    .B(\u_cpu.ALU.u_wallace._0315_ ),
    .C(\u_cpu.ALU.u_wallace._3399_ ),
    .D(\u_cpu.ALU.SrcA[29] ),
    .X(\u_cpu.ALU.u_wallace._4266_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._9736_  (.A1(\u_cpu.ALU.u_wallace._4088_ ),
    .A2(\u_cpu.ALU.u_wallace._3058_ ),
    .A3(\u_cpu.ALU.u_wallace._4663_ ),
    .B1(\u_cpu.ALU.u_wallace._4266_ ),
    .X(\u_cpu.ALU.u_wallace._4267_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9737_  (.A1(\u_cpu.ALU.u_wallace._2198_ ),
    .A2(\u_cpu.ALU.u_wallace._4100_ ),
    .B1(\u_cpu.ALU.u_wallace._4267_ ),
    .Y(\u_cpu.ALU.u_wallace._4268_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9738_  (.A(\u_cpu.ALU.u_wallace._4267_ ),
    .B(\u_cpu.ALU.u_wallace._4100_ ),
    .C(\u_cpu.ALU.u_wallace._2198_ ),
    .Y(\u_cpu.ALU.u_wallace._4270_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.ALU.u_wallace._9739_  (.A(\u_cpu.ALU.u_wallace._4268_ ),
    .B_N(\u_cpu.ALU.u_wallace._4270_ ),
    .X(\u_cpu.ALU.u_wallace._4271_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9740_  (.A1(\u_cpu.ALU.u_wallace._4262_ ),
    .A2(\u_cpu.ALU.u_wallace._4265_ ),
    .B1(\u_cpu.ALU.u_wallace._4271_ ),
    .X(\u_cpu.ALU.u_wallace._4272_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9741_  (.A(\u_cpu.ALU.u_wallace._3719_ ),
    .B(\u_cpu.ALU.u_wallace._2569_ ),
    .Y(\u_cpu.ALU.u_wallace._4273_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9742_  (.A(\u_cpu.ALU.u_wallace._1578_ ),
    .B(\u_cpu.ALU.u_wallace._3718_ ),
    .Y(\u_cpu.ALU.u_wallace._4274_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9743_  (.A(\u_cpu.ALU.u_wallace._0884_ ),
    .B(\u_cpu.ALU.SrcA[30] ),
    .Y(\u_cpu.ALU.u_wallace._4275_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9744_  (.A1(\u_cpu.ALU.u_wallace._4273_ ),
    .A2(\u_cpu.ALU.u_wallace._4274_ ),
    .B1(\u_cpu.ALU.u_wallace._4275_ ),
    .Y(\u_cpu.ALU.u_wallace._4276_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9745_  (.A(\u_cpu.ALU.u_wallace._0315_ ),
    .B(\u_cpu.ALU.SrcA[29] ),
    .Y(\u_cpu.ALU.u_wallace._4277_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.ALU.u_wallace._9746_  (.A1(\u_cpu.ALU.u_wallace._4082_ ),
    .A2(\u_cpu.ALU.u_wallace._4276_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4277_ ),
    .X(\u_cpu.ALU.u_wallace._4278_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU.u_wallace._9747_  (.A1(\u_cpu.ALU.u_wallace._4934_ ),
    .A2(\u_cpu.ALU.u_wallace._4080_ ),
    .A3(\u_cpu.ALU.u_wallace._4081_ ),
    .B1(\u_cpu.ALU.u_wallace._4078_ ),
    .C1(\u_cpu.ALU.u_wallace._4277_ ),
    .X(\u_cpu.ALU.u_wallace._4279_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9748_  (.A(\u_cpu.ALU.u_wallace._3719_ ),
    .B(\u_cpu.ALU.u_wallace._3449_ ),
    .Y(\u_cpu.ALU.u_wallace._4281_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9749_  (.A1(\u_cpu.ALU.u_wallace._0884_ ),
    .A2(\u_cpu.ALU.SrcA[31] ),
    .B1(\u_cpu.ALU.u_wallace._4281_ ),
    .X(\u_cpu.ALU.u_wallace._4282_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9750_  (.A(\u_cpu.ALU.u_wallace._4281_ ),
    .B(\u_cpu.ALU.SrcA[31] ),
    .C(\u_cpu.ALU.u_wallace._0097_ ),
    .Y(\u_cpu.ALU.u_wallace._4283_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9751_  (.A(\u_cpu.ALU.u_wallace._0652_ ),
    .B(\u_cpu.ALU.u_wallace._3718_ ),
    .Y(\u_cpu.ALU.u_wallace._4284_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9752_  (.A1(\u_cpu.ALU.u_wallace._4282_ ),
    .A2(\u_cpu.ALU.u_wallace._4283_ ),
    .B1(\u_cpu.ALU.u_wallace._4284_ ),
    .X(\u_cpu.ALU.u_wallace._4285_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9753_  (.A(\u_cpu.ALU.u_wallace._4284_ ),
    .B(\u_cpu.ALU.u_wallace._4282_ ),
    .C(\u_cpu.ALU.u_wallace._4283_ ),
    .Y(\u_cpu.ALU.u_wallace._4286_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9754_  (.A(\u_cpu.ALU.u_wallace._4285_ ),
    .B(\u_cpu.ALU.u_wallace._4286_ ),
    .Y(\u_cpu.ALU.u_wallace._4287_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9755_  (.A(\u_cpu.ALU.u_wallace._4663_ ),
    .B(\u_cpu.ALU.u_wallace._3399_ ),
    .Y(\u_cpu.ALU.u_wallace._4288_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._9756_  (.A1(\u_cpu.ALU.u_wallace._4278_ ),
    .A2(\u_cpu.ALU.u_wallace._4279_ ),
    .A3(\u_cpu.ALU.u_wallace._4287_ ),
    .B1(\u_cpu.ALU.u_wallace._4288_ ),
    .X(\u_cpu.ALU.u_wallace._4289_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9757_  (.A1(\u_cpu.ALU.u_wallace._4278_ ),
    .A2(\u_cpu.ALU.u_wallace._4279_ ),
    .B1(\u_cpu.ALU.u_wallace._4287_ ),
    .Y(\u_cpu.ALU.u_wallace._4290_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9758_  (.A1(\u_cpu.ALU.u_wallace._4082_ ),
    .A2(\u_cpu.ALU.u_wallace._4276_ ),
    .B1(\u_cpu.ALU.u_wallace._0315_ ),
    .C1(\u_cpu.ALU.SrcA[29] ),
    .Y(\u_cpu.ALU.u_wallace._4292_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._9759_  (.A1(\u_cpu.ALU.u_wallace._0315_ ),
    .A2(\u_cpu.ALU.SrcA[29] ),
    .B1(\u_cpu.ALU.u_wallace._4082_ ),
    .C1(\u_cpu.ALU.u_wallace._4276_ ),
    .X(\u_cpu.ALU.u_wallace._4293_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9760_  (.A(\u_cpu.ALU.u_wallace._4285_ ),
    .B(\u_cpu.ALU.u_wallace._4286_ ),
    .C(\u_cpu.ALU.u_wallace._4292_ ),
    .D(\u_cpu.ALU.u_wallace._4293_ ),
    .Y(\u_cpu.ALU.u_wallace._4294_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9761_  (.A1(\u_cpu.ALU.u_wallace._4294_ ),
    .A2(\u_cpu.ALU.u_wallace._4290_ ),
    .B1(\u_cpu.ALU.u_wallace._4288_ ),
    .Y(\u_cpu.ALU.u_wallace._4295_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9762_  (.A1(\u_cpu.ALU.u_wallace._4289_ ),
    .A2(\u_cpu.ALU.u_wallace._4290_ ),
    .B1(\u_cpu.ALU.u_wallace._4295_ ),
    .Y(\u_cpu.ALU.u_wallace._4296_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9763_  (.A(\u_cpu.ALU.u_wallace._4267_ ),
    .B(\u_cpu.ALU.u_wallace._4100_ ),
    .C(\u_cpu.ALU.u_wallace._2198_ ),
    .X(\u_cpu.ALU.u_wallace._4297_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9764_  (.A1(\u_cpu.ALU.u_wallace._4268_ ),
    .A2(\u_cpu.ALU.u_wallace._4297_ ),
    .B1(\u_cpu.ALU.u_wallace._4262_ ),
    .C1(\u_cpu.ALU.u_wallace._4265_ ),
    .Y(\u_cpu.ALU.u_wallace._4298_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9765_  (.A(\u_cpu.ALU.u_wallace._4272_ ),
    .B(\u_cpu.ALU.u_wallace._4296_ ),
    .C(\u_cpu.ALU.u_wallace._4298_ ),
    .Y(\u_cpu.ALU.u_wallace._4299_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9766_  (.A(\u_cpu.ALU.u_wallace._4288_ ),
    .B(\u_cpu.ALU.u_wallace._4294_ ),
    .C(\u_cpu.ALU.u_wallace._4290_ ),
    .X(\u_cpu.ALU.u_wallace._4300_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9767_  (.A1(\u_cpu.ALU.u_wallace._4268_ ),
    .A2(\u_cpu.ALU.u_wallace._4297_ ),
    .B1(\u_cpu.ALU.u_wallace._4262_ ),
    .C1(\u_cpu.ALU.u_wallace._4265_ ),
    .X(\u_cpu.ALU.u_wallace._4301_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9768_  (.A1(\u_cpu.ALU.u_wallace._4262_ ),
    .A2(\u_cpu.ALU.u_wallace._4265_ ),
    .B1(\u_cpu.ALU.u_wallace._4271_ ),
    .Y(\u_cpu.ALU.u_wallace._4303_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9769_  (.A1(\u_cpu.ALU.u_wallace._4295_ ),
    .A2(\u_cpu.ALU.u_wallace._4300_ ),
    .B1(\u_cpu.ALU.u_wallace._4301_ ),
    .B2(\u_cpu.ALU.u_wallace._4303_ ),
    .Y(\u_cpu.ALU.u_wallace._4304_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._9770_  (.A1(\u_cpu.ALU.u_wallace._1037_ ),
    .A2(\u_cpu.ALU.u_wallace._3060_ ),
    .B1(\u_cpu.ALU.u_wallace._4123_ ),
    .B2(\u_cpu.ALU.u_wallace._4115_ ),
    .C1(\u_cpu.ALU.u_wallace._4112_ ),
    .X(\u_cpu.ALU.u_wallace._4305_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._9771_  (.A1(\u_cpu.ALU.u_wallace._4111_ ),
    .A2(\u_cpu.ALU.u_wallace._2882_ ),
    .A3(\u_cpu.ALU.u_wallace._2917_ ),
    .B1(\u_cpu.ALU.u_wallace._4114_ ),
    .X(\u_cpu.ALU.u_wallace._4306_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9772_  (.A(\u_cpu.ALU.u_wallace._4306_ ),
    .B(\u_cpu.ALU.u_wallace._3058_ ),
    .C(\u_cpu.ALU.u_wallace._2166_ ),
    .X(\u_cpu.ALU.u_wallace._4307_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU.u_wallace._9773_  (.A(\u_cpu.ALU.u_wallace._4305_ ),
    .B(\u_cpu.ALU.u_wallace._4307_ ),
    .X(\u_cpu.ALU.u_wallace._4308_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9774_  (.A1(\u_cpu.ALU.u_wallace._4299_ ),
    .A2(\u_cpu.ALU.u_wallace._4304_ ),
    .B1(\u_cpu.ALU.u_wallace._4308_ ),
    .X(\u_cpu.ALU.u_wallace._4309_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9775_  (.A1(\u_cpu.ALU.u_wallace._2284_ ),
    .A2(\u_cpu.ALU.u_wallace._2215_ ),
    .B1(\u_cpu.ALU.u_wallace._4108_ ),
    .C1(\u_cpu.ALU.u_wallace._4146_ ),
    .X(\u_cpu.ALU.u_wallace._4310_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9776_  (.A(\u_cpu.ALU.u_wallace._2917_ ),
    .B(\u_cpu.ALU.u_wallace._2569_ ),
    .Y(\u_cpu.ALU.u_wallace._4311_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9777_  (.A1(\u_cpu.ALU.u_wallace._4108_ ),
    .A2(\u_cpu.ALU.u_wallace._4146_ ),
    .B1(\u_cpu.ALU.u_wallace._4311_ ),
    .Y(\u_cpu.ALU.u_wallace._4312_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9778_  (.A(\u_cpu.ALU.u_wallace._4310_ ),
    .B(\u_cpu.ALU.u_wallace._4312_ ),
    .Y(\u_cpu.ALU.u_wallace._4314_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9779_  (.A1(\u_cpu.ALU.u_wallace._4305_ ),
    .A2(\u_cpu.ALU.u_wallace._4307_ ),
    .B1(\u_cpu.ALU.u_wallace._4299_ ),
    .C1(\u_cpu.ALU.u_wallace._4304_ ),
    .Y(\u_cpu.ALU.u_wallace._4315_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9780_  (.A(\u_cpu.ALU.u_wallace._4309_ ),
    .B(\u_cpu.ALU.u_wallace._4314_ ),
    .C(\u_cpu.ALU.u_wallace._4315_ ),
    .Y(\u_cpu.ALU.u_wallace._4316_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9781_  (.A1(\u_cpu.ALU.u_wallace._4305_ ),
    .A2(\u_cpu.ALU.u_wallace._4307_ ),
    .B1(\u_cpu.ALU.u_wallace._4299_ ),
    .C1(\u_cpu.ALU.u_wallace._4304_ ),
    .X(\u_cpu.ALU.u_wallace._4317_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9782_  (.A1(\u_cpu.ALU.u_wallace._4299_ ),
    .A2(\u_cpu.ALU.u_wallace._4304_ ),
    .B1(\u_cpu.ALU.u_wallace._4308_ ),
    .Y(\u_cpu.ALU.u_wallace._4318_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9783_  (.A1(\u_cpu.ALU.u_wallace._4310_ ),
    .A2(\u_cpu.ALU.u_wallace._4312_ ),
    .B1(\u_cpu.ALU.u_wallace._4317_ ),
    .B2(\u_cpu.ALU.u_wallace._4318_ ),
    .Y(\u_cpu.ALU.u_wallace._4319_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9784_  (.A1(\u_cpu.ALU.u_wallace._0124_ ),
    .A2(\u_cpu.ALU.u_wallace._0809_ ),
    .B1(\u_cpu.ALU.u_wallace._4316_ ),
    .C1(\u_cpu.ALU.u_wallace._4319_ ),
    .Y(\u_cpu.ALU.u_wallace._4320_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9785_  (.A(\u_cpu.ALU.u_wallace._0117_ ),
    .B(\u_cpu.ALU.u_wallace._2916_ ),
    .Y(\u_cpu.ALU.u_wallace._4321_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9786_  (.A1(\u_cpu.ALU.u_wallace._4316_ ),
    .A2(\u_cpu.ALU.u_wallace._4319_ ),
    .B1(\u_cpu.ALU.u_wallace._4321_ ),
    .X(\u_cpu.ALU.u_wallace._4322_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9787_  (.A1(\u_cpu.ALU.u_wallace._4257_ ),
    .A2(\u_cpu.ALU.u_wallace._4259_ ),
    .B1(\u_cpu.ALU.u_wallace._4320_ ),
    .C1(\u_cpu.ALU.u_wallace._4322_ ),
    .X(\u_cpu.ALU.u_wallace._4323_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9788_  (.A1(\u_cpu.ALU.u_wallace._0124_ ),
    .A2(\u_cpu.ALU.u_wallace._0809_ ),
    .B1(\u_cpu.ALU.u_wallace._4316_ ),
    .C1(\u_cpu.ALU.u_wallace._4319_ ),
    .X(\u_cpu.ALU.u_wallace._4325_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9789_  (.A1(\u_cpu.ALU.u_wallace._4316_ ),
    .A2(\u_cpu.ALU.u_wallace._4319_ ),
    .B1(\u_cpu.ALU.u_wallace._4321_ ),
    .Y(\u_cpu.ALU.u_wallace._4326_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9790_  (.A(\u_cpu.ALU.u_wallace._4257_ ),
    .B(\u_cpu.ALU.u_wallace._4259_ ),
    .Y(\u_cpu.ALU.u_wallace._4327_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9791_  (.A1(\u_cpu.ALU.u_wallace._4325_ ),
    .A2(\u_cpu.ALU.u_wallace._4326_ ),
    .B1(\u_cpu.ALU.u_wallace._4327_ ),
    .Y(\u_cpu.ALU.u_wallace._4328_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9792_  (.A(\u_cpu.ALU.u_wallace._4029_ ),
    .B(\u_cpu.ALU.u_wallace._4605_ ),
    .C(\u_cpu.ALU.u_wallace._2618_ ),
    .D(\u_cpu.ALU.u_wallace._2882_ ),
    .X(\u_cpu.ALU.u_wallace._4329_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9793_  (.A1(\u_cpu.ALU.u_wallace._4605_ ),
    .A2(\u_cpu.ALU.u_wallace._2618_ ),
    .B1(\u_cpu.ALU.u_wallace._2882_ ),
    .B2(\u_cpu.ALU.u_wallace._4029_ ),
    .Y(\u_cpu.ALU.u_wallace._4330_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU.u_wallace._9794_  (.A1_N(\u_cpu.ALU.u_wallace._4313_ ),
    .A2_N(\u_cpu.ALU.u_wallace._2598_ ),
    .B1(\u_cpu.ALU.u_wallace._4329_ ),
    .B2(\u_cpu.ALU.u_wallace._4330_ ),
    .X(\u_cpu.ALU.u_wallace._4331_ ));
 sky130_fd_sc_hd__and4bb_2 \u_cpu.ALU.u_wallace._9795_  (.A_N(\u_cpu.ALU.u_wallace._4329_ ),
    .B_N(\u_cpu.ALU.u_wallace._4330_ ),
    .C(\u_cpu.ALU.u_wallace._4313_ ),
    .D(\u_cpu.ALU.u_wallace._2598_ ),
    .X(\u_cpu.ALU.u_wallace._4332_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU.u_wallace._9796_  (.A1_N(\u_cpu.ALU.u_wallace._4054_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4061_ ),
    .B1(\u_cpu.ALU.u_wallace._4331_ ),
    .B2(\u_cpu.ALU.u_wallace._4332_ ),
    .X(\u_cpu.ALU.u_wallace._4333_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9797_  (.A(\u_cpu.ALU.u_wallace._4331_ ),
    .B(\u_cpu.ALU.u_wallace._4332_ ),
    .Y(\u_cpu.ALU.u_wallace._4334_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9798_  (.A(\u_cpu.ALU.u_wallace._4054_ ),
    .B(\u_cpu.ALU.u_wallace._4061_ ),
    .C(\u_cpu.ALU.u_wallace._4334_ ),
    .X(\u_cpu.ALU.u_wallace._4336_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9799_  (.A(\u_cpu.ALU.u_wallace._4333_ ),
    .B(\u_cpu.ALU.u_wallace._4336_ ),
    .Y(\u_cpu.ALU.u_wallace._4337_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9800_  (.A(\u_cpu.ALU.u_wallace._4328_ ),
    .B(\u_cpu.ALU.u_wallace._4337_ ),
    .Y(\u_cpu.ALU.u_wallace._4338_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._9801_  (.A1(\u_cpu.ALU.u_wallace._4325_ ),
    .A2(\u_cpu.ALU.u_wallace._4326_ ),
    .B1(\u_cpu.ALU.u_wallace._4327_ ),
    .X(\u_cpu.ALU.u_wallace._4339_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9802_  (.A1(\u_cpu.ALU.u_wallace._4333_ ),
    .A2(\u_cpu.ALU.u_wallace._4336_ ),
    .B1(\u_cpu.ALU.u_wallace._4323_ ),
    .B2(\u_cpu.ALU.u_wallace._4339_ ),
    .Y(\u_cpu.ALU.u_wallace._4340_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9803_  (.A1(\u_cpu.ALU.u_wallace._4323_ ),
    .A2(\u_cpu.ALU.u_wallace._4338_ ),
    .B1(\u_cpu.ALU.u_wallace._4340_ ),
    .Y(\u_cpu.ALU.u_wallace._4341_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9804_  (.A(\u_cpu.ALU.u_wallace._4894_ ),
    .B(\u_cpu.ALU.u_wallace._2907_ ),
    .Y(\u_cpu.ALU.u_wallace._4342_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU.u_wallace._9805_  (.A1_N(\u_cpu.ALU.u_wallace._4043_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4044_ ),
    .B1(\u_cpu.ALU.u_wallace._1737_ ),
    .B2(\u_cpu.ALU.u_wallace._3685_ ),
    .X(\u_cpu.ALU.u_wallace._4343_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._9806_  (.A(\u_cpu.ALU.u_wallace._4342_ ),
    .B(\u_cpu.ALU.u_wallace._4343_ ),
    .X(\u_cpu.ALU.u_wallace._4344_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._9807_  (.A(\u_cpu.ALU.u_wallace._4344_ ),
    .Y(\u_cpu.ALU.u_wallace._4345_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9808_  (.A1(\u_cpu.ALU.u_wallace._4147_ ),
    .A2(\u_cpu.ALU.u_wallace._4157_ ),
    .B1(\u_cpu.ALU.u_wallace._4345_ ),
    .Y(\u_cpu.ALU.u_wallace._4347_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU.u_wallace._9809_  (.A1(\u_cpu.ALU.u_wallace._4149_ ),
    .A2(\u_cpu.ALU.u_wallace._4151_ ),
    .A3(\u_cpu.ALU.u_wallace._4152_ ),
    .B1(\u_cpu.ALU.u_wallace._4345_ ),
    .C1(\u_cpu.ALU.u_wallace._4147_ ),
    .X(\u_cpu.ALU.u_wallace._4348_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9810_  (.A(\u_cpu.ALU.u_wallace._4347_ ),
    .B(\u_cpu.ALU.u_wallace._4348_ ),
    .Y(\u_cpu.ALU.u_wallace._4349_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._9811_  (.A(\u_cpu.ALU.u_wallace._4349_ ),
    .Y(\u_cpu.ALU.u_wallace._4350_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.ALU.u_wallace._9812_  (.A1(\u_cpu.ALU.u_wallace._0607_ ),
    .A2(\u_cpu.ALU.u_wallace._1855_ ),
    .B1(\u_cpu.ALU.u_wallace._3986_ ),
    .B2(\u_cpu.ALU.u_wallace._3987_ ),
    .Y(\u_cpu.ALU.u_wallace._4351_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9813_  (.A(\u_cpu.ALU.u_wallace._3987_ ),
    .B(\u_cpu.ALU.u_wallace._1855_ ),
    .C(\u_cpu.ALU.u_wallace._0607_ ),
    .D(\u_cpu.ALU.u_wallace._3986_ ),
    .X(\u_cpu.ALU.u_wallace._4352_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU.u_wallace._9814_  (.A(\u_cpu.ALU.u_wallace._4351_ ),
    .B(\u_cpu.ALU.u_wallace._4352_ ),
    .X(\u_cpu.ALU.u_wallace._4353_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9815_  (.A1(\u_cpu.ALU.u_wallace._4341_ ),
    .A2(\u_cpu.ALU.u_wallace._4350_ ),
    .B1(\u_cpu.ALU.u_wallace._4353_ ),
    .Y(\u_cpu.ALU.u_wallace._4354_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9816_  (.A1(\u_cpu.ALU.u_wallace._4147_ ),
    .A2(\u_cpu.ALU.u_wallace._4157_ ),
    .B1(\u_cpu.ALU.u_wallace._4344_ ),
    .Y(\u_cpu.ALU.u_wallace._4355_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU.u_wallace._9817_  (.A1(\u_cpu.ALU.u_wallace._4149_ ),
    .A2(\u_cpu.ALU.u_wallace._4151_ ),
    .A3(\u_cpu.ALU.u_wallace._4152_ ),
    .B1(\u_cpu.ALU.u_wallace._4344_ ),
    .C1(\u_cpu.ALU.u_wallace._4147_ ),
    .X(\u_cpu.ALU.u_wallace._4356_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.ALU.u_wallace._9818_  (.A1(\u_cpu.ALU.u_wallace._4355_ ),
    .A2(\u_cpu.ALU.u_wallace._4356_ ),
    .B1(\u_cpu.ALU.u_wallace._4323_ ),
    .B2(\u_cpu.ALU.u_wallace._4338_ ),
    .C1(\u_cpu.ALU.u_wallace._4340_ ),
    .Y(\u_cpu.ALU.u_wallace._4358_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9819_  (.A(\u_cpu.ALU.u_wallace._1129_ ),
    .B(\u_cpu.ALU.u_wallace._1578_ ),
    .C(\u_cpu.ALU.u_wallace._0959_ ),
    .D(\u_cpu.ALU.u_wallace._1615_ ),
    .X(\u_cpu.ALU.u_wallace._4359_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._9820_  (.A1(\u_cpu.ALU.u_wallace._0458_ ),
    .A2(\u_cpu.ALU.u_wallace._0973_ ),
    .B1(\u_cpu.ALU.u_wallace._2053_ ),
    .B2(\u_cpu.ALU.u_wallace._0169_ ),
    .X(\u_cpu.ALU.u_wallace._4360_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9821_  (.A1(\u_cpu.ALU.u_wallace._4359_ ),
    .A2(\u_cpu.ALU.u_wallace._4360_ ),
    .B1(\u_cpu.ALU.u_wallace._2658_ ),
    .C1(\u_cpu.ALU.u_wallace._1176_ ),
    .X(\u_cpu.ALU.u_wallace._4361_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU.u_wallace._9822_  (.A1(\u_cpu.ALU.u_wallace._2658_ ),
    .A2(\u_cpu.ALU.u_wallace._1176_ ),
    .B1(\u_cpu.ALU.u_wallace._4359_ ),
    .C1(\u_cpu.ALU.u_wallace._4360_ ),
    .Y(\u_cpu.ALU.u_wallace._4362_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.ALU.u_wallace._9823_  (.A1(\u_cpu.ALU.u_wallace._4063_ ),
    .A2(\u_cpu.ALU.u_wallace._4070_ ),
    .B1(\u_cpu.ALU.u_wallace._4361_ ),
    .C1(\u_cpu.ALU.u_wallace._4362_ ),
    .X(\u_cpu.ALU.u_wallace._4363_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9824_  (.A1(\u_cpu.ALU.u_wallace._4361_ ),
    .A2(\u_cpu.ALU.u_wallace._4362_ ),
    .B1(\u_cpu.ALU.u_wallace._4063_ ),
    .C1(\u_cpu.ALU.u_wallace._4070_ ),
    .Y(\u_cpu.ALU.u_wallace._4364_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9825_  (.A(\u_cpu.ALU.u_wallace._4363_ ),
    .B(\u_cpu.ALU.u_wallace._4364_ ),
    .Y(\u_cpu.ALU.u_wallace._4365_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.ALU.u_wallace._9826_  (.A(\u_cpu.ALU.u_wallace._4365_ ),
    .Y(\u_cpu.ALU.u_wallace._4366_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9827_  (.A(\u_cpu.ALU.u_wallace._0124_ ),
    .B(\u_cpu.ALU.u_wallace._0809_ ),
    .Y(\u_cpu.ALU.u_wallace._4367_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9828_  (.A(\u_cpu.ALU.u_wallace._4316_ ),
    .B(\u_cpu.ALU.u_wallace._4319_ ),
    .Y(\u_cpu.ALU.u_wallace._4369_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._9829_  (.A1_N(\u_cpu.ALU.u_wallace._4367_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4369_ ),
    .B1(\u_cpu.ALU.u_wallace._4257_ ),
    .B2(\u_cpu.ALU.u_wallace._4259_ ),
    .Y(\u_cpu.ALU.u_wallace._4370_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9830_  (.A1(\u_cpu.ALU.u_wallace._4325_ ),
    .A2(\u_cpu.ALU.u_wallace._4370_ ),
    .B1(\u_cpu.ALU.u_wallace._4337_ ),
    .C1(\u_cpu.ALU.u_wallace._4328_ ),
    .X(\u_cpu.ALU.u_wallace._4371_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9831_  (.A1(\u_cpu.ALU.u_wallace._4257_ ),
    .A2(\u_cpu.ALU.u_wallace._4259_ ),
    .B1(\u_cpu.ALU.u_wallace._4320_ ),
    .C1(\u_cpu.ALU.u_wallace._4322_ ),
    .Y(\u_cpu.ALU.u_wallace._4372_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9832_  (.A1(\u_cpu.ALU.u_wallace._4372_ ),
    .A2(\u_cpu.ALU.u_wallace._4328_ ),
    .B1(\u_cpu.ALU.u_wallace._4337_ ),
    .Y(\u_cpu.ALU.u_wallace._4373_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.ALU.u_wallace._9833_  (.A1(\u_cpu.ALU.u_wallace._4347_ ),
    .A2(\u_cpu.ALU.u_wallace._4348_ ),
    .B1(\u_cpu.ALU.u_wallace._4371_ ),
    .B2(\u_cpu.ALU.u_wallace._4373_ ),
    .Y(\u_cpu.ALU.u_wallace._4374_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._9834_  (.A1(\u_cpu.ALU.u_wallace._4358_ ),
    .A2(\u_cpu.ALU.u_wallace._4374_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4353_ ),
    .Y(\u_cpu.ALU.u_wallace._4375_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU.u_wallace._9835_  (.A1(\u_cpu.ALU.u_wallace._4354_ ),
    .A2(\u_cpu.ALU.u_wallace._4358_ ),
    .B1(\u_cpu.ALU.u_wallace._4366_ ),
    .C1(\u_cpu.ALU.u_wallace._4375_ ),
    .Y(\u_cpu.ALU.u_wallace._4376_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9836_  (.A1(\u_cpu.ALU.u_wallace._4350_ ),
    .A2(\u_cpu.ALU.u_wallace._4341_ ),
    .B1(\u_cpu.ALU.u_wallace._4354_ ),
    .Y(\u_cpu.ALU.u_wallace._4377_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.ALU.u_wallace._9837_  (.A1(\u_cpu.ALU.u_wallace._4355_ ),
    .A2(\u_cpu.ALU.u_wallace._4356_ ),
    .B1(\u_cpu.ALU.u_wallace._4323_ ),
    .B2(\u_cpu.ALU.u_wallace._4338_ ),
    .C1(\u_cpu.ALU.u_wallace._4340_ ),
    .X(\u_cpu.ALU.u_wallace._4378_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.ALU.u_wallace._9838_  (.A1(\u_cpu.ALU.u_wallace._4347_ ),
    .A2(\u_cpu.ALU.u_wallace._4348_ ),
    .B1(\u_cpu.ALU.u_wallace._4371_ ),
    .B2(\u_cpu.ALU.u_wallace._4373_ ),
    .X(\u_cpu.ALU.u_wallace._4380_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9839_  (.A1(\u_cpu.ALU.u_wallace._4378_ ),
    .A2(\u_cpu.ALU.u_wallace._4380_ ),
    .B1(\u_cpu.ALU.u_wallace._4353_ ),
    .Y(\u_cpu.ALU.u_wallace._4381_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9840_  (.A1(\u_cpu.ALU.u_wallace._4377_ ),
    .A2(\u_cpu.ALU.u_wallace._4381_ ),
    .B1(\u_cpu.ALU.u_wallace._4365_ ),
    .Y(\u_cpu.ALU.u_wallace._4382_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9841_  (.A1(\u_cpu.ALU.u_wallace._4894_ ),
    .A2(\u_cpu.ALU.u_wallace._2916_ ),
    .B1(\u_cpu.ALU.u_wallace._2907_ ),
    .B2(\u_cpu.ALU.u_wallace._4733_ ),
    .X(\u_cpu.ALU.u_wallace._4383_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.ALU.u_wallace._9842_  (.A1(\u_cpu.ALU.u_wallace._4383_ ),
    .A2(\u_cpu.ALU.u_wallace._2621_ ),
    .A3(\u_cpu.ALU.u_wallace._0117_ ),
    .B1(\u_cpu.ALU.u_wallace._4056_ ),
    .X(\u_cpu.ALU.u_wallace._4384_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.ALU.u_wallace._9843_  (.A1(\u_cpu.ALU.u_wallace._0122_ ),
    .A2(\u_cpu.ALU.u_wallace._2621_ ),
    .B1(\u_cpu.ALU.u_wallace._4001_ ),
    .B2(\u_cpu.ALU.u_wallace._4000_ ),
    .C1(\u_cpu.ALU.u_wallace._4004_ ),
    .X(\u_cpu.ALU.u_wallace._4385_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.ALU.u_wallace._9844_  (.A1(\u_cpu.ALU.u_wallace._4004_ ),
    .A2(\u_cpu.ALU.u_wallace._4002_ ),
    .B1(\u_cpu.ALU.u_wallace._0122_ ),
    .C1(\u_cpu.ALU.u_wallace._2621_ ),
    .Y(\u_cpu.ALU.u_wallace._4386_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.ALU.u_wallace._9845_  (.A1_N(\u_cpu.ALU.u_wallace._4385_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4386_ ),
    .B1(\u_cpu.ALU.u_wallace._1324_ ),
    .B2(\u_cpu.ALU.u_wallace._0554_ ),
    .X(\u_cpu.ALU.u_wallace._4387_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.ALU.u_wallace._9846_  (.A(\u_cpu.ALU.u_wallace._4386_ ),
    .B(\u_cpu.ALU.u_wallace._3204_ ),
    .C(\u_cpu.ALU.u_wallace._1974_ ),
    .D(\u_cpu.ALU.u_wallace._4385_ ),
    .X(\u_cpu.ALU.u_wallace._4388_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU.u_wallace._9847_  (.A(\u_cpu.ALU.u_wallace._4387_ ),
    .B(\u_cpu.ALU.u_wallace._4388_ ),
    .X(\u_cpu.ALU.u_wallace._4389_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9848_  (.A(\u_cpu.ALU.u_wallace._4384_ ),
    .B(\u_cpu.ALU.u_wallace._4389_ ),
    .Y(\u_cpu.ALU.u_wallace._4391_ ));
 sky130_fd_sc_hd__a311o_2 \u_cpu.ALU.u_wallace._9849_  (.A1(\u_cpu.ALU.u_wallace._0117_ ),
    .A2(\u_cpu.ALU.u_wallace._2621_ ),
    .A3(\u_cpu.ALU.u_wallace._4383_ ),
    .B1(\u_cpu.ALU.u_wallace._4056_ ),
    .C1(\u_cpu.ALU.u_wallace._4389_ ),
    .X(\u_cpu.ALU.u_wallace._4392_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9850_  (.A1(\u_cpu.ALU.u_wallace._4033_ ),
    .A2(\u_cpu.ALU.u_wallace._4030_ ),
    .B1(\u_cpu.ALU.u_wallace._4391_ ),
    .C1(\u_cpu.ALU.u_wallace._4392_ ),
    .X(\u_cpu.ALU.u_wallace._4393_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.ALU.u_wallace._9851_  (.A1(\u_cpu.ALU.u_wallace._4391_ ),
    .A2(\u_cpu.ALU.u_wallace._4392_ ),
    .B1(\u_cpu.ALU.u_wallace._4033_ ),
    .C1(\u_cpu.ALU.u_wallace._4030_ ),
    .Y(\u_cpu.ALU.u_wallace._4394_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9852_  (.A(\u_cpu.ALU.u_wallace._4393_ ),
    .B(\u_cpu.ALU.u_wallace._4394_ ),
    .Y(\u_cpu.ALU.u_wallace._4395_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._9853_  (.A1(\u_cpu.ALU.u_wallace._4376_ ),
    .A2(\u_cpu.ALU.u_wallace._4382_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4395_ ),
    .Y(\u_cpu.ALU.u_wallace._4396_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9854_  (.A1(\u_cpu.ALU.u_wallace._4377_ ),
    .A2(\u_cpu.ALU.u_wallace._4381_ ),
    .B1(\u_cpu.ALU.u_wallace._4365_ ),
    .X(\u_cpu.ALU.u_wallace._4397_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._9855_  (.A_N(\u_cpu.ALU.u_wallace._4376_ ),
    .B(\u_cpu.ALU.u_wallace._4397_ ),
    .C(\u_cpu.ALU.u_wallace._4395_ ),
    .Y(\u_cpu.ALU.u_wallace._4398_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.ALU.u_wallace._9856_  (.A1(\u_cpu.ALU.u_wallace._4038_ ),
    .A2(\u_cpu.ALU.u_wallace._4041_ ),
    .A3(\u_cpu.ALU.u_wallace._4156_ ),
    .B1(\u_cpu.ALU.u_wallace._4162_ ),
    .X(\u_cpu.ALU.u_wallace._4399_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.ALU.u_wallace._9857_  (.A1(\u_cpu.ALU.u_wallace._3911_ ),
    .A2(\u_cpu.ALU.u_wallace._3967_ ),
    .A3(\u_cpu.ALU.u_wallace._3971_ ),
    .B1(\u_cpu.ALU.u_wallace._4181_ ),
    .Y(\u_cpu.ALU.u_wallace._4400_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9858_  (.A1(\u_cpu.ALU.u_wallace._0847_ ),
    .A2(\u_cpu.ALU.u_wallace._1611_ ),
    .B1(\u_cpu.ALU.SrcB[31] ),
    .B2(\u_cpu.ALU.u_wallace._1886_ ),
    .X(\u_cpu.ALU.u_wallace._4402_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.ALU.u_wallace._9859_  (.A(\u_cpu.ALU.u_wallace._1886_ ),
    .B(\u_cpu.ALU.u_wallace._0847_ ),
    .C(\u_cpu.ALU.u_wallace._1611_ ),
    .D(\u_cpu.ALU.SrcB[31] ),
    .Y(\u_cpu.ALU.u_wallace._4403_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9860_  (.A(\u_cpu.ALU.u_wallace._4402_ ),
    .B(\u_cpu.ALU.u_wallace._4403_ ),
    .Y(\u_cpu.ALU.u_wallace._4404_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.ALU.u_wallace._9861_  (.A1(\u_cpu.ALU.u_wallace._4021_ ),
    .A2(\u_cpu.ALU.u_wallace._4015_ ),
    .B1(\u_cpu.ALU.u_wallace._0280_ ),
    .C1(\u_cpu.ALU.u_wallace._2248_ ),
    .X(\u_cpu.ALU.u_wallace._4405_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.ALU.u_wallace._9862_  (.A1(\u_cpu.ALU.u_wallace._4020_ ),
    .A2(\u_cpu.ALU.u_wallace._4002_ ),
    .A3(\u_cpu.ALU.u_wallace._4005_ ),
    .B1(\u_cpu.ALU.u_wallace._4023_ ),
    .C1(\u_cpu.ALU.u_wallace._3999_ ),
    .X(\u_cpu.ALU.u_wallace._4406_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9863_  (.A(\u_cpu.ALU.u_wallace._4405_ ),
    .B(\u_cpu.ALU.u_wallace._4406_ ),
    .Y(\u_cpu.ALU.u_wallace._4407_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._9864_  (.A(\u_cpu.ALU.u_wallace._4404_ ),
    .B(\u_cpu.ALU.u_wallace._4407_ ),
    .X(\u_cpu.ALU.u_wallace._4408_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu.ALU.u_wallace._9865_  (.A(\u_cpu.ALU.u_wallace._4400_ ),
    .B(\u_cpu.ALU.u_wallace._4408_ ),
    .Y(\u_cpu.ALU.u_wallace._4409_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._9866_  (.A(\u_cpu.ALU.u_wallace._4399_ ),
    .B(\u_cpu.ALU.u_wallace._4409_ ),
    .X(\u_cpu.ALU.u_wallace._4410_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9867_  (.A1(\u_cpu.ALU.u_wallace._4396_ ),
    .A2(\u_cpu.ALU.u_wallace._4398_ ),
    .B1(\u_cpu.ALU.u_wallace._4410_ ),
    .X(\u_cpu.ALU.u_wallace._4411_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9868_  (.A(\u_cpu.ALU.u_wallace._4396_ ),
    .B(\u_cpu.ALU.u_wallace._4398_ ),
    .C(\u_cpu.ALU.u_wallace._4410_ ),
    .Y(\u_cpu.ALU.u_wallace._4413_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9869_  (.A(\u_cpu.ALU.u_wallace._4255_ ),
    .B(\u_cpu.ALU.u_wallace._4411_ ),
    .C(\u_cpu.ALU.u_wallace._4413_ ),
    .Y(\u_cpu.ALU.u_wallace._4414_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.ALU.u_wallace._9870_  (.A1(\u_cpu.ALU.u_wallace._4411_ ),
    .A2(\u_cpu.ALU.u_wallace._4413_ ),
    .B1(\u_cpu.ALU.u_wallace._4255_ ),
    .X(\u_cpu.ALU.u_wallace._4415_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._9871_  (.A_N(\u_cpu.ALU.u_wallace._4240_ ),
    .B(\u_cpu.ALU.u_wallace._4414_ ),
    .C(\u_cpu.ALU.u_wallace._4415_ ),
    .Y(\u_cpu.ALU.u_wallace._4416_ ));
 sky130_fd_sc_hd__a21bo_2 \u_cpu.ALU.u_wallace._9872_  (.A1(\u_cpu.ALU.u_wallace._4414_ ),
    .A2(\u_cpu.ALU.u_wallace._4415_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4240_ ),
    .X(\u_cpu.ALU.u_wallace._4417_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.ALU.u_wallace._9873_  (.A_N(\u_cpu.ALU.u_wallace._4231_ ),
    .B(\u_cpu.ALU.u_wallace._4416_ ),
    .C(\u_cpu.ALU.u_wallace._4417_ ),
    .Y(\u_cpu.ALU.u_wallace._4418_ ));
 sky130_fd_sc_hd__a21bo_2 \u_cpu.ALU.u_wallace._9874_  (.A1(\u_cpu.ALU.u_wallace._4416_ ),
    .A2(\u_cpu.ALU.u_wallace._4417_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4231_ ),
    .X(\u_cpu.ALU.u_wallace._4419_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.ALU.u_wallace._9875_  (.A(\u_cpu.ALU.u_wallace._4207_ ),
    .B(\u_cpu.ALU.u_wallace._4418_ ),
    .C(\u_cpu.ALU.u_wallace._4419_ ),
    .Y(\u_cpu.ALU.u_wallace._4420_ ));
 sky130_fd_sc_hd__and3b_2 \u_cpu.ALU.u_wallace._9876_  (.A_N(\u_cpu.ALU.u_wallace._4231_ ),
    .B(\u_cpu.ALU.u_wallace._4416_ ),
    .C(\u_cpu.ALU.u_wallace._4417_ ),
    .X(\u_cpu.ALU.u_wallace._4421_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.ALU.u_wallace._9877_  (.A1(\u_cpu.ALU.u_wallace._4416_ ),
    .A2(\u_cpu.ALU.u_wallace._4417_ ),
    .B1_N(\u_cpu.ALU.u_wallace._4231_ ),
    .Y(\u_cpu.ALU.u_wallace._4422_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.ALU.u_wallace._9878_  (.A1_N(\u_cpu.ALU.u_wallace._4207_ ),
    .A2_N(\u_cpu.ALU.u_wallace._4199_ ),
    .B1(\u_cpu.ALU.u_wallace._4421_ ),
    .B2(\u_cpu.ALU.u_wallace._4422_ ),
    .Y(\u_cpu.ALU.u_wallace._4424_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.ALU.u_wallace._9879_  (.A1(\u_cpu.ALU.u_wallace._4206_ ),
    .A2(\u_cpu.ALU.u_wallace._4420_ ),
    .B1(\u_cpu.ALU.u_wallace._4424_ ),
    .X(\u_cpu.ALU.Product_Wallace[31] ));
 sky130_fd_sc_hd__xor2_2 \u_cpu.ALU.u_wallace._9880_  (.A(\u_cpu.ALU.u_wallace._2494_ ),
    .B(\u_cpu.ALU.u_wallace._3317_ ),
    .X(\u_cpu.ALU.Product_Wallace[7] ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9881_  (.A1(\u_cpu.ALU.u_wallace._1738_ ),
    .A2(\u_cpu.ALU.u_wallace._2451_ ),
    .B1(\u_cpu.ALU.u_wallace._2483_ ),
    .Y(\u_cpu.ALU.u_wallace._4425_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9882_  (.A1(\u_cpu.ALU.u_wallace._0720_ ),
    .A2(\u_cpu.ALU.u_wallace._1716_ ),
    .B1(\u_cpu.ALU.u_wallace._4425_ ),
    .Y(\u_cpu.ALU.u_wallace._4426_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.ALU.u_wallace._9883_  (.A_N(\u_cpu.ALU.u_wallace._2494_ ),
    .B(\u_cpu.ALU.u_wallace._4426_ ),
    .X(\u_cpu.ALU.u_wallace._4427_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._9884_  (.A(\u_cpu.ALU.u_wallace._4427_ ),
    .X(\u_cpu.ALU.Product_Wallace[6] ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9885_  (.A(\u_cpu.ALU.u_wallace._1694_ ),
    .B(\u_cpu.ALU.u_wallace._1705_ ),
    .Y(\u_cpu.ALU.u_wallace._4428_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.ALU.u_wallace._9886_  (.A(\u_cpu.ALU.u_wallace._1092_ ),
    .B(\u_cpu.ALU.u_wallace._1103_ ),
    .Y(\u_cpu.ALU.u_wallace._4429_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.ALU.u_wallace._9887_  (.A1(\u_cpu.ALU.u_wallace._0676_ ),
    .A2(\u_cpu.ALU.u_wallace._0720_ ),
    .B1(\u_cpu.ALU.u_wallace._4429_ ),
    .Y(\u_cpu.ALU.u_wallace._4430_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu.ALU.u_wallace._9888_  (.A(\u_cpu.ALU.u_wallace._4428_ ),
    .B(\u_cpu.ALU.u_wallace._4430_ ),
    .Y(\u_cpu.ALU.Product_Wallace[5] ));
 sky130_fd_sc_hd__and3_2 \u_cpu.ALU.u_wallace._9889_  (.A(\u_cpu.ALU.u_wallace._0676_ ),
    .B(\u_cpu.ALU.u_wallace._0720_ ),
    .C(\u_cpu.ALU.u_wallace._4429_ ),
    .X(\u_cpu.ALU.u_wallace._4432_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.ALU.u_wallace._9890_  (.A(\u_cpu.ALU.u_wallace._4430_ ),
    .B(\u_cpu.ALU.u_wallace._4432_ ),
    .Y(\u_cpu.ALU.Product_Wallace[4] ));
 sky130_fd_sc_hd__or2_2 \u_cpu.ALU.u_wallace._9891_  (.A(\u_cpu.ALU.u_wallace._0381_ ),
    .B(\u_cpu.ALU.u_wallace._0435_ ),
    .X(\u_cpu.ALU.u_wallace._4433_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.ALU.u_wallace._9892_  (.A1(\u_cpu.ALU.u_wallace._0239_ ),
    .A2(\u_cpu.ALU.u_wallace._4433_ ),
    .B1_N(\u_cpu.ALU.u_wallace._0709_ ),
    .Y(\u_cpu.ALU.u_wallace._4434_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._9893_  (.A(\u_cpu.ALU.u_wallace._0720_ ),
    .B(\u_cpu.ALU.u_wallace._4434_ ),
    .X(\u_cpu.ALU.u_wallace._4435_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._9894_  (.A(\u_cpu.ALU.u_wallace._4435_ ),
    .X(\u_cpu.ALU.Product_Wallace[3] ));
 sky130_fd_sc_hd__or3_2 \u_cpu.ALU.u_wallace._9895_  (.A(\u_cpu.ALU.u_wallace._0435_ ),
    .B(\u_cpu.ALU.u_wallace._0239_ ),
    .C(\u_cpu.ALU.u_wallace._0381_ ),
    .X(\u_cpu.ALU.u_wallace._4436_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.ALU.u_wallace._9896_  (.A1(\u_cpu.ALU.u_wallace._0381_ ),
    .A2(\u_cpu.ALU.u_wallace._0435_ ),
    .B1(\u_cpu.ALU.u_wallace._0239_ ),
    .Y(\u_cpu.ALU.u_wallace._4437_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._9897_  (.A(\u_cpu.ALU.u_wallace._4436_ ),
    .B(\u_cpu.ALU.u_wallace._4437_ ),
    .X(\u_cpu.ALU.u_wallace._4438_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._9898_  (.A(\u_cpu.ALU.u_wallace._4438_ ),
    .X(\u_cpu.ALU.Product_Wallace[2] ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.ALU.u_wallace._9899_  (.A1(\u_cpu.ALU.u_wallace._0097_ ),
    .A2(\u_cpu.ALU.u_wallace._0184_ ),
    .B1(\u_cpu.ALU.u_wallace._0228_ ),
    .B2(\u_cpu.ALU.u_wallace._1886_ ),
    .X(\u_cpu.ALU.u_wallace._4440_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.ALU.u_wallace._9900_  (.A(\u_cpu.ALU.u_wallace._0239_ ),
    .B(\u_cpu.ALU.u_wallace._4440_ ),
    .X(\u_cpu.ALU.u_wallace._4441_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.ALU.u_wallace._9901_  (.A(\u_cpu.ALU.u_wallace._4441_ ),
    .X(\u_cpu.ALU.Product_Wallace[1] ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0928_  (.A(\u_cpu.IMEM.a[8] ),
    .X(\u_cpu.IMEM._0295_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0929_  (.A(\u_cpu.IMEM._0295_ ),
    .X(\u_cpu.IMEM._0305_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0930_  (.A(\u_cpu.IMEM.a[9] ),
    .X(\u_cpu.IMEM._0316_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0931_  (.A(\u_cpu.IMEM.a[4] ),
    .X(\u_cpu.IMEM._0327_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.IMEM._0932_  (.A(\u_cpu.IMEM._0327_ ),
    .Y(\u_cpu.IMEM._0338_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.IMEM._0933_  (.A(\u_cpu.IMEM.a[3] ),
    .B_N(\u_cpu.IMEM.a[2] ),
    .X(\u_cpu.IMEM._0349_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0934_  (.A(\u_cpu.IMEM._0349_ ),
    .X(\u_cpu.IMEM._0359_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0935_  (.A(\u_cpu.IMEM.a[3] ),
    .X(\u_cpu.IMEM._0370_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.IMEM._0936_  (.A(\u_cpu.IMEM.a[2] ),
    .B_N(\u_cpu.IMEM._0370_ ),
    .X(\u_cpu.IMEM._0381_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0937_  (.A(\u_cpu.IMEM._0381_ ),
    .X(\u_cpu.IMEM._0392_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.IMEM._0938_  (.A(\u_cpu.IMEM._0338_ ),
    .B(\u_cpu.IMEM._0359_ ),
    .C(\u_cpu.IMEM._0392_ ),
    .Y(\u_cpu.IMEM._0403_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0939_  (.A(\u_cpu.IMEM._0403_ ),
    .X(\u_cpu.IMEM._0413_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0940_  (.A(\u_cpu.IMEM.a[5] ),
    .X(\u_cpu.IMEM._0424_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0941_  (.A(\u_cpu.IMEM._0424_ ),
    .X(\u_cpu.IMEM._0434_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0942_  (.A(\u_cpu.IMEM._0434_ ),
    .X(\u_cpu.IMEM._0445_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.IMEM._0943_  (.A(\u_cpu.IMEM._0370_ ),
    .B_N(\u_cpu.IMEM._0327_ ),
    .X(\u_cpu.IMEM._0456_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0944_  (.A(\u_cpu.IMEM._0456_ ),
    .X(\u_cpu.IMEM._0466_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0945_  (.A(\u_cpu.IMEM._0370_ ),
    .X(\u_cpu.IMEM._0477_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0946_  (.A(\u_cpu.IMEM.a[2] ),
    .X(\u_cpu.IMEM._0487_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._0947_  (.A1(\u_cpu.IMEM._0477_ ),
    .A2(\u_cpu.IMEM._0487_ ),
    .B1(\u_cpu.IMEM._0338_ ),
    .Y(\u_cpu.IMEM._0498_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0948_  (.A(\u_cpu.IMEM._0477_ ),
    .X(\u_cpu.IMEM._0509_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0949_  (.A(\u_cpu.IMEM._0327_ ),
    .X(\u_cpu.IMEM._0519_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0950_  (.A(\u_cpu.IMEM.a[5] ),
    .X(\u_cpu.IMEM._0530_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._0951_  (.A1(\u_cpu.IMEM._0509_ ),
    .A2(\u_cpu.IMEM._0519_ ),
    .B1(\u_cpu.IMEM._0530_ ),
    .Y(\u_cpu.IMEM._0540_ ));
 sky130_fd_sc_hd__a32oi_2 \u_cpu.IMEM._0952_  (.A1(\u_cpu.IMEM._0413_ ),
    .A2(\u_cpu.IMEM._0445_ ),
    .A3(\u_cpu.IMEM._0466_ ),
    .B1(\u_cpu.IMEM._0498_ ),
    .B2(\u_cpu.IMEM._0540_ ),
    .Y(\u_cpu.IMEM._0551_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0953_  (.A(\u_cpu.IMEM.a[2] ),
    .X(\u_cpu.IMEM._0562_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.IMEM._0954_  (.A_N(\u_cpu.IMEM._0562_ ),
    .B(\u_cpu.IMEM._0370_ ),
    .X(\u_cpu.IMEM._0572_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0955_  (.A(\u_cpu.IMEM._0572_ ),
    .X(\u_cpu.IMEM._0583_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.IMEM._0956_  (.A(\u_cpu.IMEM.a[6] ),
    .Y(\u_cpu.IMEM._0594_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0957_  (.A(\u_cpu.IMEM._0594_ ),
    .X(\u_cpu.IMEM._0604_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0958_  (.A(\u_cpu.IMEM._0604_ ),
    .X(\u_cpu.IMEM._0615_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0959_  (.A(\u_cpu.IMEM._0327_ ),
    .X(\u_cpu.IMEM._0626_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0960_  (.A(\u_cpu.IMEM._0626_ ),
    .X(\u_cpu.IMEM._0636_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0961_  (.A(\u_cpu.IMEM._0636_ ),
    .X(\u_cpu.IMEM._0646_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0962_  (.A(\u_cpu.IMEM.a[7] ),
    .X(\u_cpu.IMEM._0657_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0963_  (.A(\u_cpu.IMEM._0657_ ),
    .X(\u_cpu.IMEM._0667_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._0964_  (.A1(\u_cpu.IMEM._0583_ ),
    .A2(\u_cpu.IMEM._0615_ ),
    .A3(\u_cpu.IMEM._0646_ ),
    .B1(\u_cpu.IMEM._0667_ ),
    .X(\u_cpu.IMEM._0678_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.IMEM._0965_  (.A(\u_cpu.IMEM.a[7] ),
    .Y(\u_cpu.IMEM._0689_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0966_  (.A(\u_cpu.IMEM._0689_ ),
    .X(\u_cpu.IMEM._0699_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0967_  (.A(\u_cpu.IMEM._0699_ ),
    .X(\u_cpu.IMEM._0710_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0968_  (.A(\u_cpu.IMEM._0594_ ),
    .X(\u_cpu.IMEM._0721_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0969_  (.A(\u_cpu.IMEM._0721_ ),
    .X(\u_cpu.IMEM._0731_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.IMEM._0970_  (.A(\u_cpu.IMEM.a[5] ),
    .Y(\u_cpu.IMEM._0742_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0971_  (.A(\u_cpu.IMEM._0742_ ),
    .X(\u_cpu.IMEM._0753_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0972_  (.A(\u_cpu.IMEM._0753_ ),
    .X(\u_cpu.IMEM._0763_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.IMEM._0973_  (.A(\u_cpu.IMEM._0477_ ),
    .B(\u_cpu.IMEM._0562_ ),
    .X(\u_cpu.IMEM._0774_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0974_  (.A(\u_cpu.IMEM.a[4] ),
    .X(\u_cpu.IMEM._0785_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0975_  (.A(\u_cpu.IMEM._0785_ ),
    .X(\u_cpu.IMEM._0795_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._0976_  (.A(\u_cpu.IMEM._0370_ ),
    .B(\u_cpu.IMEM._0562_ ),
    .Y(\u_cpu.IMEM._0806_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0977_  (.A(\u_cpu.IMEM._0806_ ),
    .X(\u_cpu.IMEM._0816_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.IMEM._0978_  (.A(\u_cpu.IMEM._0477_ ),
    .B(\u_cpu.IMEM._0327_ ),
    .Y(\u_cpu.IMEM._0827_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.IMEM._0979_  (.A1(\u_cpu.IMEM._0774_ ),
    .A2(\u_cpu.IMEM._0795_ ),
    .A3(\u_cpu.IMEM._0816_ ),
    .B1(\u_cpu.IMEM._0827_ ),
    .Y(\u_cpu.IMEM._0837_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0980_  (.A(\u_cpu.IMEM._0338_ ),
    .X(\u_cpu.IMEM._0848_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0981_  (.A(\u_cpu.IMEM._0848_ ),
    .X(\u_cpu.IMEM._0858_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.IMEM._0982_  (.A(\u_cpu.IMEM._0370_ ),
    .B(\u_cpu.IMEM._0562_ ),
    .Y(\u_cpu.IMEM._0868_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0983_  (.A(\u_cpu.IMEM._0868_ ),
    .X(\u_cpu.IMEM._0879_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0984_  (.A(\u_cpu.IMEM._0530_ ),
    .X(\u_cpu.IMEM._0889_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._0985_  (.A1(\u_cpu.IMEM._0848_ ),
    .A2(\u_cpu.IMEM._0816_ ),
    .B1(\u_cpu.IMEM._0889_ ),
    .Y(\u_cpu.IMEM._0899_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._0986_  (.A1(\u_cpu.IMEM._0858_ ),
    .A2(\u_cpu.IMEM._0879_ ),
    .B1(\u_cpu.IMEM._0899_ ),
    .Y(\u_cpu.IMEM._0910_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0987_  (.A(\u_cpu.IMEM._0848_ ),
    .X(\u_cpu.IMEM._0920_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0988_  (.A(\u_cpu.IMEM._0477_ ),
    .X(\u_cpu.IMEM._0927_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0989_  (.A(\u_cpu.IMEM._0927_ ),
    .X(\u_cpu.IMEM._0000_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0990_  (.A(\u_cpu.IMEM._0530_ ),
    .X(\u_cpu.IMEM._0001_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0991_  (.A(\u_cpu.IMEM._0001_ ),
    .X(\u_cpu.IMEM._0002_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0992_  (.A(\u_cpu.IMEM._0594_ ),
    .X(\u_cpu.IMEM._0003_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.IMEM._0993_  (.A1(\u_cpu.IMEM._0920_ ),
    .A2(\u_cpu.IMEM._0000_ ),
    .B1(\u_cpu.IMEM._0002_ ),
    .C1(\u_cpu.IMEM._0003_ ),
    .D1(\u_cpu.IMEM._0413_ ),
    .Y(\u_cpu.IMEM._0004_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._0994_  (.A1(\u_cpu.IMEM._0731_ ),
    .A2(\u_cpu.IMEM._0763_ ),
    .A3(\u_cpu.IMEM._0837_ ),
    .B1(\u_cpu.IMEM._0910_ ),
    .C1(\u_cpu.IMEM._0004_ ),
    .X(\u_cpu.IMEM._0005_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.IMEM._0995_  (.A1(\u_cpu.IMEM._0551_ ),
    .A2(\u_cpu.IMEM._0678_ ),
    .B1(\u_cpu.IMEM._0710_ ),
    .B2(\u_cpu.IMEM._0005_ ),
    .Y(\u_cpu.IMEM._0006_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0996_  (.A(\u_cpu.IMEM.a[6] ),
    .X(\u_cpu.IMEM._0007_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0997_  (.A(\u_cpu.IMEM._0007_ ),
    .X(\u_cpu.IMEM._0008_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._0998_  (.A(\u_cpu.IMEM._0530_ ),
    .X(\u_cpu.IMEM._0009_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._0999_  (.A(\u_cpu.IMEM._0008_ ),
    .B(\u_cpu.IMEM._0009_ ),
    .Y(\u_cpu.IMEM._0010_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1000_  (.A(\u_cpu.IMEM._0424_ ),
    .X(\u_cpu.IMEM._0011_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1001_  (.A(\u_cpu.IMEM._0785_ ),
    .X(\u_cpu.IMEM._0012_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1002_  (.A(\u_cpu.IMEM._0012_ ),
    .X(\u_cpu.IMEM._0013_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1003_  (.A(\u_cpu.IMEM._0392_ ),
    .X(\u_cpu.IMEM._0014_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1004_  (.A(\u_cpu.IMEM._0007_ ),
    .X(\u_cpu.IMEM._0015_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1005_  (.A1(\u_cpu.IMEM._0011_ ),
    .A2(\u_cpu.IMEM._0013_ ),
    .A3(\u_cpu.IMEM._0014_ ),
    .B1(\u_cpu.IMEM._0015_ ),
    .X(\u_cpu.IMEM._0016_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1006_  (.A(\u_cpu.IMEM._0370_ ),
    .X(\u_cpu.IMEM._0017_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1007_  (.A(\u_cpu.IMEM._0017_ ),
    .B(\u_cpu.IMEM._0785_ ),
    .Y(\u_cpu.IMEM._0018_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1008_  (.A(\u_cpu.IMEM._0562_ ),
    .X(\u_cpu.IMEM._0019_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1009_  (.A(\u_cpu.IMEM._0019_ ),
    .X(\u_cpu.IMEM._0020_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.IMEM._1010_  (.A(\u_cpu.IMEM._0370_ ),
    .Y(\u_cpu.IMEM._0021_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.IMEM._1011_  (.A(\u_cpu.IMEM.a[2] ),
    .Y(\u_cpu.IMEM._0022_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1012_  (.A(\u_cpu.IMEM._0022_ ),
    .X(\u_cpu.IMEM._0023_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1013_  (.A(\u_cpu.IMEM._0785_ ),
    .X(\u_cpu.IMEM._0024_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.IMEM._1014_  (.A(\u_cpu.IMEM._0021_ ),
    .B(\u_cpu.IMEM._0023_ ),
    .C(\u_cpu.IMEM._0024_ ),
    .D(\u_cpu.IMEM._0889_ ),
    .Y(\u_cpu.IMEM._0025_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1015_  (.A1(\u_cpu.IMEM._0011_ ),
    .A2(\u_cpu.IMEM._0018_ ),
    .A3(\u_cpu.IMEM._0020_ ),
    .B1(\u_cpu.IMEM._0604_ ),
    .C1(\u_cpu.IMEM._0025_ ),
    .X(\u_cpu.IMEM._0026_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.IMEM._1016_  (.A1(\u_cpu.IMEM._0413_ ),
    .A2(\u_cpu.IMEM._0010_ ),
    .B1(\u_cpu.IMEM._0016_ ),
    .B2(\u_cpu.IMEM._0026_ ),
    .Y(\u_cpu.IMEM._0027_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1017_  (.A(\u_cpu.IMEM._0667_ ),
    .X(\u_cpu.IMEM._0028_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1018_  (.A(\u_cpu.IMEM._0027_ ),
    .B(\u_cpu.IMEM._0028_ ),
    .Y(\u_cpu.IMEM._0029_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1019_  (.A(\u_cpu.IMEM._0795_ ),
    .X(\u_cpu.IMEM._0030_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.IMEM._1020_  (.A(\u_cpu.IMEM._0370_ ),
    .B(\u_cpu.IMEM._0562_ ),
    .X(\u_cpu.IMEM._0031_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1021_  (.A(\u_cpu.IMEM._0031_ ),
    .X(\u_cpu.IMEM._0032_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1022_  (.A(\u_cpu.IMEM._0032_ ),
    .X(\u_cpu.IMEM._0033_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1023_  (.A(\u_cpu.IMEM._0487_ ),
    .X(\u_cpu.IMEM._0034_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.IMEM._1024_  (.A1(\u_cpu.IMEM._0509_ ),
    .A2(\u_cpu.IMEM._0034_ ),
    .A3(\u_cpu.IMEM._0012_ ),
    .B1(\u_cpu.IMEM._0889_ ),
    .Y(\u_cpu.IMEM._0035_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1025_  (.A1(\u_cpu.IMEM._0030_ ),
    .A2(\u_cpu.IMEM._0033_ ),
    .B1(\u_cpu.IMEM._0035_ ),
    .Y(\u_cpu.IMEM._0036_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1026_  (.A(\u_cpu.IMEM._0689_ ),
    .X(\u_cpu.IMEM._0037_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1027_  (.A(\u_cpu.IMEM._0007_ ),
    .X(\u_cpu.IMEM._0038_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1028_  (.A(\u_cpu.IMEM._0037_ ),
    .B(\u_cpu.IMEM._0038_ ),
    .Y(\u_cpu.IMEM._0039_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1029_  (.A(\u_cpu.IMEM._0795_ ),
    .X(\u_cpu.IMEM._0040_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1030_  (.A(\u_cpu.IMEM._0827_ ),
    .X(\u_cpu.IMEM._0041_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1031_  (.A(\u_cpu.IMEM._0034_ ),
    .X(\u_cpu.IMEM._0042_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1032_  (.A(\u_cpu.IMEM._0530_ ),
    .X(\u_cpu.IMEM._0043_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1033_  (.A(\u_cpu.IMEM._0043_ ),
    .X(\u_cpu.IMEM._0044_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.IMEM._1034_  (.A1(\u_cpu.IMEM._0040_ ),
    .A2(\u_cpu.IMEM._0879_ ),
    .B1(\u_cpu.IMEM._0041_ ),
    .B2(\u_cpu.IMEM._0042_ ),
    .C1(\u_cpu.IMEM._0044_ ),
    .Y(\u_cpu.IMEM._0045_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1035_  (.A(\u_cpu.IMEM._0007_ ),
    .X(\u_cpu.IMEM._0046_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.IMEM._1036_  (.A(\u_cpu.IMEM._0657_ ),
    .B(\u_cpu.IMEM._0046_ ),
    .X(\u_cpu.IMEM._0047_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1037_  (.A(\u_cpu.IMEM._0774_ ),
    .X(\u_cpu.IMEM._0048_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1038_  (.A(\u_cpu.IMEM._0019_ ),
    .X(\u_cpu.IMEM._0049_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1039_  (.A1(\u_cpu.IMEM._0049_ ),
    .A2(\u_cpu.IMEM._0848_ ),
    .B1(\u_cpu.IMEM._0001_ ),
    .Y(\u_cpu.IMEM._0050_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1040_  (.A(\u_cpu.IMEM._0519_ ),
    .X(\u_cpu.IMEM._0051_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1041_  (.A1(\u_cpu.IMEM._0023_ ),
    .A2(\u_cpu.IMEM._0927_ ),
    .B1(\u_cpu.IMEM._0051_ ),
    .Y(\u_cpu.IMEM._0052_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.IMEM._1042_  (.A1(\u_cpu.IMEM._0011_ ),
    .A2(\u_cpu.IMEM._0013_ ),
    .A3(\u_cpu.IMEM._0048_ ),
    .B1(\u_cpu.IMEM._0050_ ),
    .B2(\u_cpu.IMEM._0052_ ),
    .X(\u_cpu.IMEM._0053_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.IMEM._1043_  (.A1(\u_cpu.IMEM._0036_ ),
    .A2(\u_cpu.IMEM._0039_ ),
    .A3(\u_cpu.IMEM._0045_ ),
    .B1(\u_cpu.IMEM._0047_ ),
    .B2(\u_cpu.IMEM._0053_ ),
    .X(\u_cpu.IMEM._0054_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1044_  (.A(\u_cpu.IMEM.a[9] ),
    .X(\u_cpu.IMEM._0055_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1045_  (.A1(\u_cpu.IMEM._0029_ ),
    .A2(\u_cpu.IMEM._0054_ ),
    .B1(\u_cpu.IMEM._0055_ ),
    .Y(\u_cpu.IMEM._0056_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1046_  (.A1(\u_cpu.IMEM._0316_ ),
    .A2(\u_cpu.IMEM._0006_ ),
    .B1(\u_cpu.IMEM._0056_ ),
    .Y(\u_cpu.IMEM._0057_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1047_  (.A(\u_cpu.IMEM._0015_ ),
    .X(\u_cpu.IMEM._0058_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1048_  (.A(\u_cpu.IMEM._0338_ ),
    .X(\u_cpu.IMEM._0059_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1049_  (.A(\u_cpu.IMEM._0017_ ),
    .X(\u_cpu.IMEM._0060_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1050_  (.A(\u_cpu.IMEM._0742_ ),
    .X(\u_cpu.IMEM._0061_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1051_  (.A1(\u_cpu.IMEM._0059_ ),
    .A2(\u_cpu.IMEM._0060_ ),
    .B1(\u_cpu.IMEM._0061_ ),
    .C1(\u_cpu.IMEM._0403_ ),
    .Y(\u_cpu.IMEM._0062_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1052_  (.A1(\u_cpu.IMEM._0017_ ),
    .A2(\u_cpu.IMEM._0487_ ),
    .B1(\u_cpu.IMEM._0519_ ),
    .X(\u_cpu.IMEM._0063_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1053_  (.A(\u_cpu.IMEM._0043_ ),
    .X(\u_cpu.IMEM._0064_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1054_  (.A1(\u_cpu.IMEM._0509_ ),
    .A2(\u_cpu.IMEM._0019_ ),
    .B1(\u_cpu.IMEM._0012_ ),
    .Y(\u_cpu.IMEM._0065_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1055_  (.A(\u_cpu.IMEM.a[7] ),
    .X(\u_cpu.IMEM._0066_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.IMEM._1056_  (.A1(\u_cpu.IMEM._0063_ ),
    .A2(\u_cpu.IMEM._0064_ ),
    .A3(\u_cpu.IMEM._0065_ ),
    .B1(\u_cpu.IMEM._0066_ ),
    .Y(\u_cpu.IMEM._0067_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.IMEM._1057_  (.A_N(\u_cpu.IMEM._0868_ ),
    .B(\u_cpu.IMEM._0012_ ),
    .C(\u_cpu.IMEM._0816_ ),
    .Y(\u_cpu.IMEM._0068_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.IMEM._1058_  (.A(\u_cpu.IMEM._0477_ ),
    .B(\u_cpu.IMEM._0785_ ),
    .X(\u_cpu.IMEM._0069_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1059_  (.A(\u_cpu.IMEM._0742_ ),
    .X(\u_cpu.IMEM._0070_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1060_  (.A(\u_cpu.IMEM._0070_ ),
    .B(\u_cpu.IMEM._0007_ ),
    .Y(\u_cpu.IMEM._0071_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1061_  (.A1(\u_cpu.IMEM._0068_ ),
    .A2(\u_cpu.IMEM._0069_ ),
    .B1(\u_cpu.IMEM._0071_ ),
    .X(\u_cpu.IMEM._0072_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.IMEM._1062_  (.A1(\u_cpu.IMEM._0058_ ),
    .A2(\u_cpu.IMEM._0062_ ),
    .B1(\u_cpu.IMEM._0067_ ),
    .C1(\u_cpu.IMEM._0072_ ),
    .X(\u_cpu.IMEM._0073_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1063_  (.A(\u_cpu.IMEM._0022_ ),
    .B(\u_cpu.IMEM._0785_ ),
    .Y(\u_cpu.IMEM._0074_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1064_  (.A(\u_cpu.IMEM._0017_ ),
    .X(\u_cpu.IMEM._0075_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.IMEM._1065_  (.A(\u_cpu.IMEM._0074_ ),
    .B(\u_cpu.IMEM._0075_ ),
    .C(\u_cpu.IMEM._0043_ ),
    .X(\u_cpu.IMEM._0076_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1066_  (.A(\u_cpu.IMEM._0037_ ),
    .X(\u_cpu.IMEM._0077_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1067_  (.A(\u_cpu.IMEM._0359_ ),
    .X(\u_cpu.IMEM._0078_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.IMEM._1068_  (.A1(\u_cpu.IMEM._0509_ ),
    .A2(\u_cpu.IMEM._0019_ ),
    .B1_N(\u_cpu.IMEM._0519_ ),
    .X(\u_cpu.IMEM._0079_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1069_  (.A(\u_cpu.IMEM._0889_ ),
    .X(\u_cpu.IMEM._0080_ ));
 sky130_fd_sc_hd__a311oi_2 \u_cpu.IMEM._1070_  (.A1(\u_cpu.IMEM._0078_ ),
    .A2(\u_cpu.IMEM._0014_ ),
    .A3(\u_cpu.IMEM._0040_ ),
    .B1(\u_cpu.IMEM._0079_ ),
    .C1(\u_cpu.IMEM._0080_ ),
    .Y(\u_cpu.IMEM._0081_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1071_  (.A(\u_cpu.IMEM._0530_ ),
    .X(\u_cpu.IMEM._0082_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1072_  (.A(\u_cpu.IMEM._0626_ ),
    .X(\u_cpu.IMEM._0083_ ));
 sky130_fd_sc_hd__or4_2 \u_cpu.IMEM._1073_  (.A(\u_cpu.IMEM._0007_ ),
    .B(\u_cpu.IMEM._0082_ ),
    .C(\u_cpu.IMEM._0060_ ),
    .D(\u_cpu.IMEM._0083_ ),
    .X(\u_cpu.IMEM._0084_ ));
 sky130_fd_sc_hd__nor4b_2 \u_cpu.IMEM._1074_  (.A(\u_cpu.IMEM._0076_ ),
    .B(\u_cpu.IMEM._0077_ ),
    .C(\u_cpu.IMEM._0081_ ),
    .D_N(\u_cpu.IMEM._0084_ ),
    .Y(\u_cpu.IMEM._0085_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1075_  (.A(\u_cpu.IMEM._0021_ ),
    .X(\u_cpu.IMEM._0086_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.IMEM._1076_  (.A_N(\u_cpu.IMEM._0562_ ),
    .B(\u_cpu.IMEM._0327_ ),
    .X(\u_cpu.IMEM._0087_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1077_  (.A(\u_cpu.IMEM._0087_ ),
    .X(\u_cpu.IMEM._0088_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.IMEM._1078_  (.A(\u_cpu.IMEM._0001_ ),
    .B(\u_cpu.IMEM._0086_ ),
    .C(\u_cpu.IMEM._0088_ ),
    .X(\u_cpu.IMEM._0089_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1079_  (.A(\u_cpu.IMEM._0066_ ),
    .X(\u_cpu.IMEM._0090_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.IMEM._1080_  (.A(\u_cpu.IMEM.a[9] ),
    .Y(\u_cpu.IMEM._0091_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1081_  (.A1(\u_cpu.IMEM._0089_ ),
    .A2(\u_cpu.IMEM._0090_ ),
    .B1(\u_cpu.IMEM._0091_ ),
    .X(\u_cpu.IMEM._0092_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1082_  (.A(\u_cpu.IMEM._0007_ ),
    .X(\u_cpu.IMEM._0093_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1083_  (.A(\u_cpu.IMEM._0093_ ),
    .X(\u_cpu.IMEM._0094_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1084_  (.A(\u_cpu.IMEM._0742_ ),
    .X(\u_cpu.IMEM._0095_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1085_  (.A(\u_cpu.IMEM._0095_ ),
    .X(\u_cpu.IMEM._0096_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.IMEM._1086_  (.A1_N(\u_cpu.IMEM._0065_ ),
    .A2_N(\u_cpu.IMEM._0899_ ),
    .B1(\u_cpu.IMEM._0096_ ),
    .B2(\u_cpu.IMEM._0837_ ),
    .X(\u_cpu.IMEM._0097_ ));
 sky130_fd_sc_hd__nor2b_2 \u_cpu.IMEM._1087_  (.A(\u_cpu.IMEM._0519_ ),
    .B_N(\u_cpu.IMEM._0017_ ),
    .Y(\u_cpu.IMEM._0098_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1088_  (.A1(\u_cpu.IMEM._0509_ ),
    .A2(\u_cpu.IMEM._0019_ ),
    .A3(\u_cpu.IMEM._0626_ ),
    .B1(\u_cpu.IMEM._0530_ ),
    .X(\u_cpu.IMEM._0099_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1089_  (.A1(\u_cpu.IMEM._0098_ ),
    .A2(\u_cpu.IMEM._0099_ ),
    .B1(\u_cpu.IMEM._0015_ ),
    .Y(\u_cpu.IMEM._0100_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1090_  (.A(\u_cpu.IMEM._0359_ ),
    .B(\u_cpu.IMEM._0392_ ),
    .Y(\u_cpu.IMEM._0101_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1091_  (.A1(\u_cpu.IMEM._0101_ ),
    .A2(\u_cpu.IMEM._0040_ ),
    .B1(\u_cpu.IMEM._0035_ ),
    .Y(\u_cpu.IMEM._0102_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1092_  (.A(\u_cpu.IMEM._0689_ ),
    .X(\u_cpu.IMEM._0103_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.IMEM._1093_  (.A1(\u_cpu.IMEM._0100_ ),
    .A2(\u_cpu.IMEM._0102_ ),
    .B1(\u_cpu.IMEM._0103_ ),
    .X(\u_cpu.IMEM._0104_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.IMEM._1094_  (.A1(\u_cpu.IMEM._0094_ ),
    .A2(\u_cpu.IMEM._0097_ ),
    .B1(\u_cpu.IMEM._0104_ ),
    .X(\u_cpu.IMEM._0105_ ));
 sky130_fd_sc_hd__o32ai_2 \u_cpu.IMEM._1095_  (.A1(\u_cpu.IMEM._0055_ ),
    .A2(\u_cpu.IMEM._0073_ ),
    .A3(\u_cpu.IMEM._0085_ ),
    .B1(\u_cpu.IMEM._0092_ ),
    .B2(\u_cpu.IMEM._0105_ ),
    .Y(\u_cpu.IMEM._0106_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1096_  (.A(\u_cpu.IMEM._0106_ ),
    .B(\u_cpu.IMEM._0305_ ),
    .Y(\u_cpu.IMEM._0107_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1097_  (.A1(\u_cpu.IMEM._0305_ ),
    .A2(\u_cpu.IMEM._0057_ ),
    .B1(\u_cpu.IMEM._0107_ ),
    .Y(\u_cpu.IMEM.rd[2] ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1098_  (.A(\u_cpu.IMEM._0055_ ),
    .X(\u_cpu.IMEM._0108_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.IMEM._1099_  (.A(\u_cpu.IMEM.a[8] ),
    .Y(\u_cpu.IMEM._0109_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.IMEM._1100_  (.A(\u_cpu.IMEM._0109_ ),
    .B(\u_cpu.IMEM._0037_ ),
    .Y(\u_cpu.IMEM._0110_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.IMEM._1101_  (.A(\u_cpu.IMEM._0562_ ),
    .B(\u_cpu.IMEM._0327_ ),
    .X(\u_cpu.IMEM._0111_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1102_  (.A(\u_cpu.IMEM._0742_ ),
    .X(\u_cpu.IMEM._0112_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.IMEM._1103_  (.A(\u_cpu.IMEM._0111_ ),
    .B(\u_cpu.IMEM._0112_ ),
    .C(\u_cpu.IMEM._0927_ ),
    .X(\u_cpu.IMEM._0113_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1104_  (.A(\u_cpu.IMEM._0090_ ),
    .X(\u_cpu.IMEM._0114_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1105_  (.A(\u_cpu.IMEM._0001_ ),
    .B(\u_cpu.IMEM._0051_ ),
    .Y(\u_cpu.IMEM._0115_ ));
 sky130_fd_sc_hd__or4_2 \u_cpu.IMEM._1106_  (.A(\u_cpu.IMEM._0038_ ),
    .B(\u_cpu.IMEM._0000_ ),
    .C(\u_cpu.IMEM._0042_ ),
    .D(\u_cpu.IMEM._0115_ ),
    .X(\u_cpu.IMEM._0116_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1107_  (.A(\u_cpu.IMEM._0295_ ),
    .X(\u_cpu.IMEM._0117_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1108_  (.A(\u_cpu.IMEM._0019_ ),
    .B(\u_cpu.IMEM._0827_ ),
    .Y(\u_cpu.IMEM._0118_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1109_  (.A(\u_cpu.IMEM._0118_ ),
    .X(\u_cpu.IMEM._0119_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.IMEM._1110_  (.A(\u_cpu.IMEM._0021_ ),
    .B(\u_cpu.IMEM._0626_ ),
    .C(\u_cpu.IMEM._0424_ ),
    .Y(\u_cpu.IMEM._0120_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1111_  (.A(\u_cpu.IMEM._0023_ ),
    .X(\u_cpu.IMEM._0121_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.IMEM._1112_  (.A1(\u_cpu.IMEM._0044_ ),
    .A2(\u_cpu.IMEM._0030_ ),
    .A3(\u_cpu.IMEM._0048_ ),
    .B1(\u_cpu.IMEM._0120_ ),
    .B2(\u_cpu.IMEM._0121_ ),
    .X(\u_cpu.IMEM._0122_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1113_  (.A(\u_cpu.IMEM._0008_ ),
    .X(\u_cpu.IMEM._0123_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1114_  (.A(\u_cpu.IMEM._0123_ ),
    .X(\u_cpu.IMEM._0124_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1115_  (.A(\u_cpu.IMEM._0103_ ),
    .X(\u_cpu.IMEM._0125_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.IMEM._1116_  (.A1(\u_cpu.IMEM._0119_ ),
    .A2(\u_cpu.IMEM._0071_ ),
    .B1(\u_cpu.IMEM._0122_ ),
    .B2(\u_cpu.IMEM._0124_ ),
    .C1(\u_cpu.IMEM._0125_ ),
    .X(\u_cpu.IMEM._0126_ ));
 sky130_fd_sc_hd__a2111oi_2 \u_cpu.IMEM._1117_  (.A1(\u_cpu.IMEM._0114_ ),
    .A2(\u_cpu.IMEM._0116_ ),
    .B1(\u_cpu.IMEM._0055_ ),
    .C1(\u_cpu.IMEM._0117_ ),
    .D1(\u_cpu.IMEM._0126_ ),
    .Y(\u_cpu.IMEM._0127_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1118_  (.A1(\u_cpu.IMEM._0108_ ),
    .A2(\u_cpu.IMEM._0110_ ),
    .A3(\u_cpu.IMEM._0113_ ),
    .B1(\u_cpu.IMEM._0127_ ),
    .X(\u_cpu.IMEM.rd[3] ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1119_  (.A(\u_cpu.IMEM._0091_ ),
    .X(\u_cpu.IMEM._0128_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1120_  (.A(\u_cpu.IMEM._0657_ ),
    .X(\u_cpu.IMEM._0129_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1121_  (.A(\u_cpu.IMEM._0129_ ),
    .X(\u_cpu.IMEM._0130_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1122_  (.A(\u_cpu.IMEM._0123_ ),
    .X(\u_cpu.IMEM._0131_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1123_  (.A(\u_cpu.IMEM._0061_ ),
    .X(\u_cpu.IMEM._0132_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1124_  (.A(\u_cpu.IMEM._0024_ ),
    .B(\u_cpu.IMEM._0032_ ),
    .Y(\u_cpu.IMEM._0133_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1125_  (.A(\u_cpu.IMEM._0742_ ),
    .X(\u_cpu.IMEM._0134_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1126_  (.A1(\u_cpu.IMEM._0040_ ),
    .A2(\u_cpu.IMEM._0879_ ),
    .B1(\u_cpu.IMEM._0134_ ),
    .Y(\u_cpu.IMEM._0135_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1127_  (.A1(\u_cpu.IMEM._0132_ ),
    .A2(\u_cpu.IMEM._0133_ ),
    .A3(\u_cpu.IMEM._0118_ ),
    .B1(\u_cpu.IMEM._0135_ ),
    .X(\u_cpu.IMEM._0136_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1128_  (.A(\u_cpu.IMEM._0689_ ),
    .X(\u_cpu.IMEM._0137_ ));
 sky130_fd_sc_hd__nor2b_2 \u_cpu.IMEM._1129_  (.A(\u_cpu.IMEM._0017_ ),
    .B_N(\u_cpu.IMEM._0519_ ),
    .Y(\u_cpu.IMEM._0138_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1130_  (.A1(\u_cpu.IMEM._0858_ ),
    .A2(\u_cpu.IMEM._0078_ ),
    .B1(\u_cpu.IMEM._0138_ ),
    .C1(\u_cpu.IMEM._0080_ ),
    .X(\u_cpu.IMEM._0139_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.IMEM._1131_  (.A1(\u_cpu.IMEM._0137_ ),
    .A2(\u_cpu.IMEM._0139_ ),
    .B1(\u_cpu.IMEM._0295_ ),
    .X(\u_cpu.IMEM._0140_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.IMEM._1132_  (.A1(\u_cpu.IMEM._0020_ ),
    .A2(\u_cpu.IMEM._0636_ ),
    .B1(\u_cpu.IMEM._0466_ ),
    .C1(\u_cpu.IMEM._0816_ ),
    .D1(\u_cpu.IMEM._0753_ ),
    .Y(\u_cpu.IMEM._0141_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.IMEM._1133_  (.A(\u_cpu.IMEM._0626_ ),
    .B(\u_cpu.IMEM._0806_ ),
    .Y(\u_cpu.IMEM._0142_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1134_  (.A(\u_cpu.IMEM._0082_ ),
    .B(\u_cpu.IMEM._0142_ ),
    .Y(\u_cpu.IMEM._0143_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1135_  (.A(\u_cpu.IMEM._0657_ ),
    .X(\u_cpu.IMEM._0144_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1136_  (.A(\u_cpu.IMEM._0003_ ),
    .X(\u_cpu.IMEM._0145_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1137_  (.A1(\u_cpu.IMEM._0141_ ),
    .A2(\u_cpu.IMEM._0143_ ),
    .B1(\u_cpu.IMEM._0144_ ),
    .C1(\u_cpu.IMEM._0145_ ),
    .X(\u_cpu.IMEM._0146_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1138_  (.A1(\u_cpu.IMEM._0130_ ),
    .A2(\u_cpu.IMEM._0131_ ),
    .A3(\u_cpu.IMEM._0136_ ),
    .B1(\u_cpu.IMEM._0140_ ),
    .C1(\u_cpu.IMEM._0146_ ),
    .X(\u_cpu.IMEM._0147_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1139_  (.A(\u_cpu.IMEM._0021_ ),
    .X(\u_cpu.IMEM._0148_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.IMEM._1140_  (.A(\u_cpu.IMEM._0562_ ),
    .B(\u_cpu.IMEM._0327_ ),
    .Y(\u_cpu.IMEM._0149_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1141_  (.A1(\u_cpu.IMEM._0149_ ),
    .A2(\u_cpu.IMEM._0111_ ),
    .B1(\u_cpu.IMEM._0112_ ),
    .Y(\u_cpu.IMEM._0150_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.IMEM._1142_  (.A1(\u_cpu.IMEM._0120_ ),
    .A2(\u_cpu.IMEM._0131_ ),
    .B1(\u_cpu.IMEM._0148_ ),
    .B2(\u_cpu.IMEM._0150_ ),
    .C1(\u_cpu.IMEM._0025_ ),
    .Y(\u_cpu.IMEM._0151_ ));
 sky130_fd_sc_hd__nor2b_2 \u_cpu.IMEM._1143_  (.A(\u_cpu.IMEM._0477_ ),
    .B_N(\u_cpu.IMEM._0487_ ),
    .Y(\u_cpu.IMEM._0152_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1144_  (.A1(\u_cpu.IMEM._0848_ ),
    .A2(\u_cpu.IMEM._0152_ ),
    .B1(\u_cpu.IMEM._0498_ ),
    .C1(\u_cpu.IMEM._0889_ ),
    .Y(\u_cpu.IMEM._0153_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.IMEM._1145_  (.A(\u_cpu.IMEM._0095_ ),
    .B(\u_cpu.IMEM._0848_ ),
    .C(\u_cpu.IMEM._0049_ ),
    .D(\u_cpu.IMEM._0075_ ),
    .Y(\u_cpu.IMEM._0154_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1146_  (.A1(\u_cpu.IMEM._0153_ ),
    .A2(\u_cpu.IMEM._0154_ ),
    .B1(\u_cpu.IMEM._0130_ ),
    .Y(\u_cpu.IMEM._0155_ ));
 sky130_fd_sc_hd__a311oi_2 \u_cpu.IMEM._1147_  (.A1(\u_cpu.IMEM._0151_ ),
    .A2(\u_cpu.IMEM._0114_ ),
    .A3(\u_cpu.IMEM._0116_ ),
    .B1(\u_cpu.IMEM._0155_ ),
    .C1(\u_cpu.IMEM._0117_ ),
    .Y(\u_cpu.IMEM._0156_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1148_  (.A(\u_cpu.IMEM._0051_ ),
    .X(\u_cpu.IMEM._0157_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1149_  (.A1(\u_cpu.IMEM._0338_ ),
    .A2(\u_cpu.IMEM._0806_ ),
    .B1(\u_cpu.IMEM._0112_ ),
    .X(\u_cpu.IMEM._0158_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1150_  (.A1(\u_cpu.IMEM._0157_ ),
    .A2(\u_cpu.IMEM._0048_ ),
    .B1(\u_cpu.IMEM._0093_ ),
    .C1(\u_cpu.IMEM._0158_ ),
    .X(\u_cpu.IMEM._0159_ ));
 sky130_fd_sc_hd__and3b_2 \u_cpu.IMEM._1151_  (.A_N(\u_cpu.IMEM._0487_ ),
    .B(\u_cpu.IMEM._0785_ ),
    .C(\u_cpu.IMEM._0477_ ),
    .X(\u_cpu.IMEM._0160_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1152_  (.A(\u_cpu.IMEM._0160_ ),
    .X(\u_cpu.IMEM._0161_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.IMEM._1153_  (.A(\u_cpu.IMEM._0509_ ),
    .B(\u_cpu.IMEM._0034_ ),
    .C(\u_cpu.IMEM._0012_ ),
    .Y(\u_cpu.IMEM._0162_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.IMEM._1154_  (.A(\u_cpu.IMEM._0434_ ),
    .B(\u_cpu.IMEM._0604_ ),
    .Y(\u_cpu.IMEM._0163_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1155_  (.A1(\u_cpu.IMEM._0161_ ),
    .A2(\u_cpu.IMEM._0162_ ),
    .B1(\u_cpu.IMEM._0163_ ),
    .Y(\u_cpu.IMEM._0164_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1156_  (.A(\u_cpu.IMEM._0359_ ),
    .X(\u_cpu.IMEM._0165_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1157_  (.A1(\u_cpu.IMEM._0165_ ),
    .A2(\u_cpu.IMEM._0014_ ),
    .B1(\u_cpu.IMEM._0040_ ),
    .Y(\u_cpu.IMEM._0166_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1158_  (.A1(\u_cpu.IMEM._0075_ ),
    .A2(\u_cpu.IMEM._0848_ ),
    .B1(\u_cpu.IMEM._0043_ ),
    .Y(\u_cpu.IMEM._0167_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1159_  (.A(\u_cpu.IMEM._0111_ ),
    .X(\u_cpu.IMEM._0168_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1160_  (.A1(\u_cpu.IMEM._0059_ ),
    .A2(\u_cpu.IMEM._0359_ ),
    .A3(\u_cpu.IMEM._0392_ ),
    .B1(\u_cpu.IMEM._0082_ ),
    .X(\u_cpu.IMEM._0169_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.IMEM._1161_  (.A1(\u_cpu.IMEM._0166_ ),
    .A2(\u_cpu.IMEM._0167_ ),
    .B1(\u_cpu.IMEM._0168_ ),
    .B2(\u_cpu.IMEM._0169_ ),
    .C1(\u_cpu.IMEM._0615_ ),
    .Y(\u_cpu.IMEM._0170_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1162_  (.A1(\u_cpu.IMEM._0646_ ),
    .A2(\u_cpu.IMEM._0583_ ),
    .A3(\u_cpu.IMEM._0071_ ),
    .B1(\u_cpu.IMEM._0137_ ),
    .X(\u_cpu.IMEM._0171_ ));
 sky130_fd_sc_hd__a32oi_2 \u_cpu.IMEM._1163_  (.A1(\u_cpu.IMEM._0130_ ),
    .A2(\u_cpu.IMEM._0159_ ),
    .A3(\u_cpu.IMEM._0164_ ),
    .B1(\u_cpu.IMEM._0170_ ),
    .B2(\u_cpu.IMEM._0171_ ),
    .Y(\u_cpu.IMEM._0172_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1164_  (.A(\u_cpu.IMEM._0144_ ),
    .X(\u_cpu.IMEM._0173_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1165_  (.A(\u_cpu.IMEM._0509_ ),
    .X(\u_cpu.IMEM._0174_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1166_  (.A(\u_cpu.IMEM._0487_ ),
    .B(\u_cpu.IMEM._0327_ ),
    .Y(\u_cpu.IMEM._0175_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1167_  (.A(\u_cpu.IMEM._0175_ ),
    .X(\u_cpu.IMEM._0176_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1168_  (.A(\u_cpu.IMEM._0530_ ),
    .B(\u_cpu.IMEM._0017_ ),
    .Y(\u_cpu.IMEM._0177_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.IMEM._1169_  (.A1(\u_cpu.IMEM._0149_ ),
    .A2(\u_cpu.IMEM._0111_ ),
    .B1_N(\u_cpu.IMEM._0177_ ),
    .Y(\u_cpu.IMEM._0178_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.IMEM._1170_  (.A1(\u_cpu.IMEM._0011_ ),
    .A2(\u_cpu.IMEM._0174_ ),
    .A3(\u_cpu.IMEM._0176_ ),
    .B1(\u_cpu.IMEM._0178_ ),
    .Y(\u_cpu.IMEM._0179_ ));
 sky130_fd_sc_hd__nor3b_2 \u_cpu.IMEM._1171_  (.A(\u_cpu.IMEM._0477_ ),
    .B(\u_cpu.IMEM._0487_ ),
    .C_N(\u_cpu.IMEM._0785_ ),
    .Y(\u_cpu.IMEM._0180_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1172_  (.A1(\u_cpu.IMEM._0001_ ),
    .A2(\u_cpu.IMEM._0180_ ),
    .B1(\u_cpu.IMEM._0008_ ),
    .Y(\u_cpu.IMEM._0181_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.IMEM._1173_  (.A1(\u_cpu.IMEM._0064_ ),
    .A2(\u_cpu.IMEM._0133_ ),
    .A3(\u_cpu.IMEM._0118_ ),
    .B1(\u_cpu.IMEM._0181_ ),
    .Y(\u_cpu.IMEM._0182_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1174_  (.A1(\u_cpu.IMEM._0145_ ),
    .A2(\u_cpu.IMEM._0179_ ),
    .B1(\u_cpu.IMEM._0182_ ),
    .Y(\u_cpu.IMEM._0183_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1175_  (.A(\u_cpu.IMEM._0487_ ),
    .X(\u_cpu.IMEM._0184_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1176_  (.A(\u_cpu.IMEM._0184_ ),
    .X(\u_cpu.IMEM._0185_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1177_  (.A1(\u_cpu.IMEM._0000_ ),
    .A2(\u_cpu.IMEM._0185_ ),
    .A3(\u_cpu.IMEM._0920_ ),
    .B1(\u_cpu.IMEM._0132_ ),
    .C1(\u_cpu.IMEM._0731_ ),
    .X(\u_cpu.IMEM._0186_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1178_  (.A(\u_cpu.IMEM._0424_ ),
    .X(\u_cpu.IMEM._0187_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1179_  (.A(\u_cpu.IMEM._0187_ ),
    .X(\u_cpu.IMEM._0188_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.IMEM._1180_  (.A_N(\u_cpu.IMEM._0487_ ),
    .B(\u_cpu.IMEM._0519_ ),
    .C(\u_cpu.IMEM._0017_ ),
    .Y(\u_cpu.IMEM._0189_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1181_  (.A(\u_cpu.IMEM._0021_ ),
    .X(\u_cpu.IMEM._0190_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1182_  (.A(\u_cpu.IMEM._0112_ ),
    .X(\u_cpu.IMEM._0191_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1183_  (.A1(\u_cpu.IMEM._0083_ ),
    .A2(\u_cpu.IMEM._0023_ ),
    .A3(\u_cpu.IMEM._0190_ ),
    .B1(\u_cpu.IMEM._0046_ ),
    .C1(\u_cpu.IMEM._0191_ ),
    .X(\u_cpu.IMEM._0192_ ));
 sky130_fd_sc_hd__a311o_2 \u_cpu.IMEM._1184_  (.A1(\u_cpu.IMEM._0188_ ),
    .A2(\u_cpu.IMEM._0189_ ),
    .A3(\u_cpu.IMEM._0119_ ),
    .B1(\u_cpu.IMEM._0699_ ),
    .C1(\u_cpu.IMEM._0192_ ),
    .X(\u_cpu.IMEM._0193_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1185_  (.A(\u_cpu.IMEM.a[8] ),
    .X(\u_cpu.IMEM._0194_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.IMEM._1186_  (.A1(\u_cpu.IMEM._0173_ ),
    .A2(\u_cpu.IMEM._0183_ ),
    .B1(\u_cpu.IMEM._0186_ ),
    .B2(\u_cpu.IMEM._0193_ ),
    .C1(\u_cpu.IMEM._0194_ ),
    .Y(\u_cpu.IMEM._0195_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1187_  (.A1(\u_cpu.IMEM._0305_ ),
    .A2(\u_cpu.IMEM._0172_ ),
    .B1(\u_cpu.IMEM._0195_ ),
    .C1(\u_cpu.IMEM._0128_ ),
    .Y(\u_cpu.IMEM._0196_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1188_  (.A1(\u_cpu.IMEM._0128_ ),
    .A2(\u_cpu.IMEM._0147_ ),
    .A3(\u_cpu.IMEM._0156_ ),
    .B1(\u_cpu.IMEM._0196_ ),
    .X(\u_cpu.IMEM.rd[4] ));
 sky130_fd_sc_hd__and3_2 \u_cpu.IMEM._1189_  (.A(\u_cpu.IMEM._0927_ ),
    .B(\u_cpu.IMEM._0034_ ),
    .C(\u_cpu.IMEM._0012_ ),
    .X(\u_cpu.IMEM._0197_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.IMEM._1190_  (.A1(\u_cpu.IMEM._0445_ ),
    .A2(\u_cpu.IMEM._0098_ ),
    .A3(\u_cpu.IMEM._0197_ ),
    .B1(\u_cpu.IMEM._0167_ ),
    .B2(\u_cpu.IMEM._0162_ ),
    .X(\u_cpu.IMEM._0198_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1191_  (.A(\u_cpu.IMEM._0066_ ),
    .X(\u_cpu.IMEM._0199_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1192_  (.A1(\u_cpu.IMEM._0774_ ),
    .A2(\u_cpu.IMEM._0013_ ),
    .B1(\u_cpu.IMEM._0721_ ),
    .C1(\u_cpu.IMEM._0158_ ),
    .X(\u_cpu.IMEM._0200_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.IMEM._1193_  (.A1(\u_cpu.IMEM._0120_ ),
    .A2(\u_cpu.IMEM._0124_ ),
    .B1(\u_cpu.IMEM._0199_ ),
    .C1(\u_cpu.IMEM._0062_ ),
    .D1(\u_cpu.IMEM._0200_ ),
    .Y(\u_cpu.IMEM._0201_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.IMEM._1194_  (.A1(\u_cpu.IMEM._0173_ ),
    .A2(\u_cpu.IMEM._0198_ ),
    .B1(\u_cpu.IMEM._0055_ ),
    .C1(\u_cpu.IMEM._0201_ ),
    .X(\u_cpu.IMEM._0202_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1195_  (.A1(\u_cpu.IMEM._0190_ ),
    .A2(\u_cpu.IMEM._0083_ ),
    .B1(\u_cpu.IMEM._0753_ ),
    .C1(\u_cpu.IMEM._0079_ ),
    .X(\u_cpu.IMEM._0203_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.IMEM._1196_  (.A1(\u_cpu.IMEM._0188_ ),
    .A2(\u_cpu.IMEM._0185_ ),
    .A3(\u_cpu.IMEM._0041_ ),
    .B1(\u_cpu.IMEM._0203_ ),
    .C1(\u_cpu.IMEM._0145_ ),
    .Y(\u_cpu.IMEM._0204_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1197_  (.A(\u_cpu.IMEM._0149_ ),
    .X(\u_cpu.IMEM._0205_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1198_  (.A1(\u_cpu.IMEM._0174_ ),
    .A2(\u_cpu.IMEM._0205_ ),
    .B1(\u_cpu.IMEM._0753_ ),
    .C1(\u_cpu.IMEM._0088_ ),
    .X(\u_cpu.IMEM._0206_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1199_  (.A1(\u_cpu.IMEM._0043_ ),
    .A2(\u_cpu.IMEM._0075_ ),
    .A3(\u_cpu.IMEM._0059_ ),
    .B1(\u_cpu.IMEM._0008_ ),
    .X(\u_cpu.IMEM._0207_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1200_  (.A(\u_cpu.IMEM._0667_ ),
    .X(\u_cpu.IMEM._0208_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1201_  (.A1(\u_cpu.IMEM._0206_ ),
    .A2(\u_cpu.IMEM._0207_ ),
    .B1(\u_cpu.IMEM._0208_ ),
    .Y(\u_cpu.IMEM._0209_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.IMEM._1202_  (.A(\u_cpu.IMEM._0370_ ),
    .B(\u_cpu.IMEM._0327_ ),
    .X(\u_cpu.IMEM._0210_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1203_  (.A(\u_cpu.IMEM._0210_ ),
    .X(\u_cpu.IMEM._0211_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1204_  (.A(\u_cpu.IMEM._0046_ ),
    .X(\u_cpu.IMEM._0212_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1205_  (.A1(\u_cpu.IMEM._0445_ ),
    .A2(\u_cpu.IMEM._0211_ ),
    .A3(\u_cpu.IMEM._0121_ ),
    .B1(\u_cpu.IMEM._0212_ ),
    .X(\u_cpu.IMEM._0213_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1206_  (.A1(\u_cpu.IMEM._0024_ ),
    .A2(\u_cpu.IMEM._0868_ ),
    .B1(\u_cpu.IMEM._0070_ ),
    .Y(\u_cpu.IMEM._0214_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.IMEM._1207_  (.A1_N(\u_cpu.IMEM._0180_ ),
    .A2_N(\u_cpu.IMEM._0214_ ),
    .B1(\u_cpu.IMEM._0413_ ),
    .B2(\u_cpu.IMEM._0188_ ),
    .Y(\u_cpu.IMEM._0215_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1208_  (.A(\u_cpu.IMEM._0174_ ),
    .X(\u_cpu.IMEM._0216_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1209_  (.A(\u_cpu.IMEM._0149_ ),
    .X(\u_cpu.IMEM._0217_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1210_  (.A(\u_cpu.IMEM._0008_ ),
    .X(\u_cpu.IMEM._0218_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1211_  (.A1(\u_cpu.IMEM._0064_ ),
    .A2(\u_cpu.IMEM._0098_ ),
    .B1(\u_cpu.IMEM._0218_ ),
    .Y(\u_cpu.IMEM._0219_ ));
 sky130_fd_sc_hd__a2111o_2 \u_cpu.IMEM._1212_  (.A1(\u_cpu.IMEM._0216_ ),
    .A2(\u_cpu.IMEM._0121_ ),
    .B1(\u_cpu.IMEM._0217_ ),
    .C1(\u_cpu.IMEM._0168_ ),
    .D1(\u_cpu.IMEM._0219_ ),
    .X(\u_cpu.IMEM._0220_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1213_  (.A1(\u_cpu.IMEM._0213_ ),
    .A2(\u_cpu.IMEM._0215_ ),
    .B1(\u_cpu.IMEM._0220_ ),
    .Y(\u_cpu.IMEM._0221_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.IMEM._1214_  (.A1(\u_cpu.IMEM._0204_ ),
    .A2(\u_cpu.IMEM._0209_ ),
    .B1(\u_cpu.IMEM._0221_ ),
    .B2(\u_cpu.IMEM._0114_ ),
    .C1(\u_cpu.IMEM._0316_ ),
    .Y(\u_cpu.IMEM._0222_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1215_  (.A1(\u_cpu.IMEM._0041_ ),
    .A2(\u_cpu.IMEM._0211_ ),
    .B1(\u_cpu.IMEM._0080_ ),
    .Y(\u_cpu.IMEM._0223_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1216_  (.A(\u_cpu.IMEM._0910_ ),
    .B(\u_cpu.IMEM._0223_ ),
    .Y(\u_cpu.IMEM._0224_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1217_  (.A(\u_cpu.IMEM._0604_ ),
    .X(\u_cpu.IMEM._0225_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.IMEM._1218_  (.A1(\u_cpu.IMEM._0445_ ),
    .A2(\u_cpu.IMEM._0138_ ),
    .B1(\u_cpu.IMEM._0413_ ),
    .C1(\u_cpu.IMEM._0120_ ),
    .D1(\u_cpu.IMEM._0225_ ),
    .X(\u_cpu.IMEM._0226_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.IMEM._1219_  (.A1(\u_cpu.IMEM._0224_ ),
    .A2(\u_cpu.IMEM._0131_ ),
    .B1(\u_cpu.IMEM._0208_ ),
    .C1(\u_cpu.IMEM._0226_ ),
    .Y(\u_cpu.IMEM._0227_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1220_  (.A(\u_cpu.IMEM._0191_ ),
    .X(\u_cpu.IMEM._0228_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1221_  (.A(\u_cpu.IMEM._0721_ ),
    .X(\u_cpu.IMEM._0229_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1222_  (.A(\u_cpu.IMEM._0082_ ),
    .X(\u_cpu.IMEM._0230_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1223_  (.A(\u_cpu.IMEM._0338_ ),
    .B(\u_cpu.IMEM._0017_ ),
    .Y(\u_cpu.IMEM._0231_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1224_  (.A1(\u_cpu.IMEM._0229_ ),
    .A2(\u_cpu.IMEM._0230_ ),
    .A3(\u_cpu.IMEM._0231_ ),
    .B1(\u_cpu.IMEM._0667_ ),
    .X(\u_cpu.IMEM._0232_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.IMEM._1225_  (.A1(\u_cpu.IMEM._0094_ ),
    .A2(\u_cpu.IMEM._0910_ ),
    .B1(\u_cpu.IMEM._0228_ ),
    .B2(\u_cpu.IMEM._0837_ ),
    .C1(\u_cpu.IMEM._0232_ ),
    .X(\u_cpu.IMEM._0233_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1226_  (.A1(\u_cpu.IMEM._0068_ ),
    .A2(\u_cpu.IMEM._0069_ ),
    .B1(\u_cpu.IMEM._0445_ ),
    .Y(\u_cpu.IMEM._0234_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.IMEM._1227_  (.A1(\u_cpu.IMEM._0060_ ),
    .A2(\u_cpu.IMEM._0049_ ),
    .B1(\u_cpu.IMEM._0001_ ),
    .X(\u_cpu.IMEM._0235_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1228_  (.A(\u_cpu.IMEM._0594_ ),
    .X(\u_cpu.IMEM._0236_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1229_  (.A(\u_cpu.IMEM._0236_ ),
    .X(\u_cpu.IMEM._0237_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1230_  (.A(\u_cpu.IMEM._0519_ ),
    .X(\u_cpu.IMEM._0238_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.IMEM._1231_  (.A(\u_cpu.IMEM._0238_ ),
    .B(\u_cpu.IMEM._0086_ ),
    .C(\u_cpu.IMEM._0061_ ),
    .X(\u_cpu.IMEM._0239_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1232_  (.A1(\u_cpu.IMEM._0848_ ),
    .A2(\u_cpu.IMEM._0879_ ),
    .B1(\u_cpu.IMEM._0063_ ),
    .C1(\u_cpu.IMEM._0082_ ),
    .Y(\u_cpu.IMEM._0240_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1233_  (.A1(\u_cpu.IMEM._0827_ ),
    .A2(\u_cpu.IMEM._0211_ ),
    .B1(\u_cpu.IMEM._0134_ ),
    .Y(\u_cpu.IMEM._0241_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1234_  (.A1(\u_cpu.IMEM._0240_ ),
    .A2(\u_cpu.IMEM._0241_ ),
    .B1(\u_cpu.IMEM._0218_ ),
    .X(\u_cpu.IMEM._0242_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.IMEM._1235_  (.A1(\u_cpu.IMEM._0237_ ),
    .A2(\u_cpu.IMEM._0239_ ),
    .B1(\u_cpu.IMEM._0242_ ),
    .C1(\u_cpu.IMEM._0072_ ),
    .D1(\u_cpu.IMEM._0077_ ),
    .Y(\u_cpu.IMEM._0243_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.IMEM._1236_  (.A1(\u_cpu.IMEM._0710_ ),
    .A2(\u_cpu.IMEM._0234_ ),
    .A3(\u_cpu.IMEM._0235_ ),
    .B1(\u_cpu.IMEM.a[9] ),
    .C1(\u_cpu.IMEM._0243_ ),
    .Y(\u_cpu.IMEM._0244_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.IMEM._1237_  (.A1(\u_cpu.IMEM._0316_ ),
    .A2(\u_cpu.IMEM._0227_ ),
    .A3(\u_cpu.IMEM._0233_ ),
    .B1(\u_cpu.IMEM._0244_ ),
    .C1(\u_cpu.IMEM._0305_ ),
    .Y(\u_cpu.IMEM._0245_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1238_  (.A1(\u_cpu.IMEM._0305_ ),
    .A2(\u_cpu.IMEM._0202_ ),
    .A3(\u_cpu.IMEM._0222_ ),
    .B1(\u_cpu.IMEM._0245_ ),
    .X(\u_cpu.IMEM.rd[5] ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1239_  (.A(\u_cpu.IMEM._0055_ ),
    .X(\u_cpu.IMEM._0246_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1240_  (.A1(\u_cpu.IMEM._0011_ ),
    .A2(\u_cpu.IMEM._0079_ ),
    .A3(\u_cpu.IMEM._0211_ ),
    .B1(\u_cpu.IMEM._0015_ ),
    .X(\u_cpu.IMEM._0247_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1241_  (.A1(\u_cpu.IMEM._0247_ ),
    .A2(\u_cpu.IMEM._0206_ ),
    .B1(\u_cpu.IMEM._0144_ ),
    .Y(\u_cpu.IMEM._0248_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.IMEM._1242_  (.A1(\u_cpu.IMEM._0248_ ),
    .A2(\u_cpu.IMEM._0204_ ),
    .B1(\u_cpu.IMEM._0316_ ),
    .C1(\u_cpu.IMEM._0117_ ),
    .Y(\u_cpu.IMEM._0249_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.IMEM._1243_  (.A(\u_cpu.IMEM._0213_ ),
    .B(\u_cpu.IMEM._0215_ ),
    .Y(\u_cpu.IMEM._0250_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1244_  (.A(\u_cpu.IMEM._0868_ ),
    .X(\u_cpu.IMEM._0251_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1245_  (.A1(\u_cpu.IMEM._0012_ ),
    .A2(\u_cpu.IMEM._0022_ ),
    .B1(\u_cpu.IMEM._0424_ ),
    .Y(\u_cpu.IMEM._0252_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.IMEM._1246_  (.A1(\u_cpu.IMEM._0188_ ),
    .A2(\u_cpu.IMEM._0098_ ),
    .B1(\u_cpu.IMEM._0251_ ),
    .B2(\u_cpu.IMEM._0252_ ),
    .C1(\u_cpu.IMEM._0131_ ),
    .X(\u_cpu.IMEM._0253_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1247_  (.A1(\u_cpu.IMEM._0250_ ),
    .A2(\u_cpu.IMEM._0253_ ),
    .B1(\u_cpu.IMEM._0114_ ),
    .Y(\u_cpu.IMEM._0254_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.IMEM._1248_  (.A1(\u_cpu.IMEM._0246_ ),
    .A2(\u_cpu.IMEM._0110_ ),
    .A3(\u_cpu.IMEM._0235_ ),
    .B1(\u_cpu.IMEM._0249_ ),
    .B2(\u_cpu.IMEM._0254_ ),
    .X(\u_cpu.IMEM.rd[6] ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1249_  (.A(\u_cpu.IMEM.a[8] ),
    .X(\u_cpu.IMEM._0255_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1250_  (.A(\u_cpu.IMEM._0206_ ),
    .B(\u_cpu.IMEM._0207_ ),
    .Y(\u_cpu.IMEM._0256_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1251_  (.A(\u_cpu.IMEM._0009_ ),
    .X(\u_cpu.IMEM._0257_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1252_  (.A1(\u_cpu.IMEM._0184_ ),
    .A2(\u_cpu.IMEM._0018_ ),
    .A3(\u_cpu.IMEM._0095_ ),
    .B1(\u_cpu.IMEM._0721_ ),
    .X(\u_cpu.IMEM._0258_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.IMEM._1253_  (.A1(\u_cpu.IMEM._0257_ ),
    .A2(\u_cpu.IMEM._0185_ ),
    .A3(\u_cpu.IMEM._0041_ ),
    .B1(\u_cpu.IMEM._0258_ ),
    .Y(\u_cpu.IMEM._0259_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1254_  (.A1(\u_cpu.IMEM._0256_ ),
    .A2(\u_cpu.IMEM._0259_ ),
    .B1(\u_cpu.IMEM._0028_ ),
    .Y(\u_cpu.IMEM._0260_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1255_  (.A1(\u_cpu.IMEM._0020_ ),
    .A2(\u_cpu.IMEM._0083_ ),
    .B1(\u_cpu.IMEM._0009_ ),
    .C1(\u_cpu.IMEM._0190_ ),
    .X(\u_cpu.IMEM._0261_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1256_  (.A(\u_cpu.IMEM._0015_ ),
    .X(\u_cpu.IMEM._0262_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.IMEM._1257_  (.A(\u_cpu.IMEM._0240_ ),
    .B(\u_cpu.IMEM._0261_ ),
    .C(\u_cpu.IMEM._0262_ ),
    .Y(\u_cpu.IMEM._0263_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.IMEM._1258_  (.A1(\u_cpu.IMEM._0763_ ),
    .A2(\u_cpu.IMEM._0176_ ),
    .B1(\u_cpu.IMEM._0180_ ),
    .B2(\u_cpu.IMEM._0214_ ),
    .C1(\u_cpu.IMEM._0225_ ),
    .Y(\u_cpu.IMEM._0264_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1259_  (.A1(\u_cpu.IMEM._0263_ ),
    .A2(\u_cpu.IMEM._0264_ ),
    .B1(\u_cpu.IMEM._0125_ ),
    .Y(\u_cpu.IMEM._0265_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.IMEM._1260_  (.A(\u_cpu.IMEM._0165_ ),
    .B(\u_cpu.IMEM._0014_ ),
    .C(\u_cpu.IMEM._0540_ ),
    .X(\u_cpu.IMEM._0266_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1261_  (.A1(\u_cpu.IMEM._0188_ ),
    .A2(\u_cpu.IMEM._0101_ ),
    .B1(\u_cpu.IMEM._0266_ ),
    .Y(\u_cpu.IMEM._0267_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1262_  (.A(\u_cpu.IMEM._0236_ ),
    .B(\u_cpu.IMEM._0657_ ),
    .Y(\u_cpu.IMEM._0268_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1263_  (.A(\u_cpu.IMEM._0059_ ),
    .B(\u_cpu.IMEM._0020_ ),
    .Y(\u_cpu.IMEM._0269_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.IMEM._1264_  (.A1(\u_cpu.IMEM._0075_ ),
    .A2(\u_cpu.IMEM._0184_ ),
    .B1(\u_cpu.IMEM._0043_ ),
    .C1(\u_cpu.IMEM._0018_ ),
    .X(\u_cpu.IMEM._0270_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1265_  (.A1(\u_cpu.IMEM._0051_ ),
    .A2(\u_cpu.IMEM._0023_ ),
    .A3(\u_cpu.IMEM._0086_ ),
    .B1(\u_cpu.IMEM._0061_ ),
    .X(\u_cpu.IMEM._0271_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1266_  (.A(\u_cpu.IMEM._0657_ ),
    .B(\u_cpu.IMEM._0008_ ),
    .Y(\u_cpu.IMEM._0272_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.IMEM._1267_  (.A1(\u_cpu.IMEM._0269_ ),
    .A2(\u_cpu.IMEM._0270_ ),
    .B1(\u_cpu.IMEM._0271_ ),
    .B2(\u_cpu.IMEM._0065_ ),
    .C1(\u_cpu.IMEM._0272_ ),
    .X(\u_cpu.IMEM._0273_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.IMEM._1268_  (.A(\u_cpu.IMEM._0043_ ),
    .B(\u_cpu.IMEM._0075_ ),
    .C(\u_cpu.IMEM._0149_ ),
    .X(\u_cpu.IMEM._0274_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1269_  (.A1(\u_cpu.IMEM._0187_ ),
    .A2(\u_cpu.IMEM._0174_ ),
    .B1(\u_cpu.IMEM._0015_ ),
    .Y(\u_cpu.IMEM._0275_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1270_  (.A1(\u_cpu.IMEM._0238_ ),
    .A2(\u_cpu.IMEM._0816_ ),
    .B1(\u_cpu.IMEM._0070_ ),
    .C1(\u_cpu.IMEM._0098_ ),
    .X(\u_cpu.IMEM._0276_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.IMEM._1271_  (.A1(\u_cpu.IMEM._0274_ ),
    .A2(\u_cpu.IMEM._0275_ ),
    .B1(\u_cpu.IMEM._0207_ ),
    .B2(\u_cpu.IMEM._0276_ ),
    .C1(\u_cpu.IMEM._0667_ ),
    .X(\u_cpu.IMEM._0277_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.IMEM._1272_  (.A1(\u_cpu.IMEM._0267_ ),
    .A2(\u_cpu.IMEM._0268_ ),
    .B1(\u_cpu.IMEM._0295_ ),
    .C1(\u_cpu.IMEM._0273_ ),
    .D1(\u_cpu.IMEM._0277_ ),
    .Y(\u_cpu.IMEM._0278_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1273_  (.A1(\u_cpu.IMEM._0255_ ),
    .A2(\u_cpu.IMEM._0260_ ),
    .A3(\u_cpu.IMEM._0265_ ),
    .B1(\u_cpu.IMEM._0278_ ),
    .X(\u_cpu.IMEM._0279_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.IMEM._1274_  (.A(\u_cpu.IMEM._0021_ ),
    .B(\u_cpu.IMEM._0019_ ),
    .C(\u_cpu.IMEM._0626_ ),
    .D(\u_cpu.IMEM._0530_ ),
    .Y(\u_cpu.IMEM._0280_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1275_  (.A(\u_cpu.IMEM._0280_ ),
    .X(\u_cpu.IMEM._0281_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1276_  (.A1(\u_cpu.IMEM._0281_ ),
    .A2(\u_cpu.IMEM._0261_ ),
    .B1(\u_cpu.IMEM._0262_ ),
    .Y(\u_cpu.IMEM._0282_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1277_  (.A1(\u_cpu.IMEM._0019_ ),
    .A2(\u_cpu.IMEM._0519_ ),
    .B1(\u_cpu.IMEM._0806_ ),
    .Y(\u_cpu.IMEM._0283_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.IMEM._1278_  (.A(\u_cpu.IMEM._0231_ ),
    .B(\u_cpu.IMEM._0007_ ),
    .C(\u_cpu.IMEM._0095_ ),
    .D(\u_cpu.IMEM._0283_ ),
    .X(\u_cpu.IMEM._0284_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.IMEM._1279_  (.A(\u_cpu.IMEM._0594_ ),
    .B(\u_cpu.IMEM._0095_ ),
    .Y(\u_cpu.IMEM._0285_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1280_  (.A1(\u_cpu.IMEM._0216_ ),
    .A2(\u_cpu.IMEM._0285_ ),
    .A3(\u_cpu.IMEM._0217_ ),
    .B1(\u_cpu.IMEM._0066_ ),
    .X(\u_cpu.IMEM._0286_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1281_  (.A(\u_cpu.IMEM._0074_ ),
    .X(\u_cpu.IMEM._0287_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.IMEM._1282_  (.A(\u_cpu.IMEM._0070_ ),
    .B(\u_cpu.IMEM._0816_ ),
    .C(\u_cpu.IMEM._0069_ ),
    .D(\u_cpu.IMEM._0287_ ),
    .X(\u_cpu.IMEM._0288_ ));
 sky130_fd_sc_hd__a311o_2 \u_cpu.IMEM._1283_  (.A1(\u_cpu.IMEM._0257_ ),
    .A2(\u_cpu.IMEM._0148_ ),
    .A3(\u_cpu.IMEM._0121_ ),
    .B1(\u_cpu.IMEM._0103_ ),
    .C1(\u_cpu.IMEM._0288_ ),
    .X(\u_cpu.IMEM._0289_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1284_  (.A1(\u_cpu.IMEM._0282_ ),
    .A2(\u_cpu.IMEM._0284_ ),
    .A3(\u_cpu.IMEM._0286_ ),
    .B1(\u_cpu.IMEM._0295_ ),
    .C1(\u_cpu.IMEM._0289_ ),
    .X(\u_cpu.IMEM._0290_ ));
 sky130_fd_sc_hd__nor3b_2 \u_cpu.IMEM._1285_  (.A(\u_cpu.IMEM._0477_ ),
    .B(\u_cpu.IMEM._0785_ ),
    .C_N(\u_cpu.IMEM._0562_ ),
    .Y(\u_cpu.IMEM._0291_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1286_  (.A1(\u_cpu.IMEM._0180_ ),
    .A2(\u_cpu.IMEM._0291_ ),
    .B1(\u_cpu.IMEM._0009_ ),
    .Y(\u_cpu.IMEM._0292_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.IMEM._1287_  (.A1(\u_cpu.IMEM._0033_ ),
    .A2(\u_cpu.IMEM._0251_ ),
    .B1(\u_cpu.IMEM._0646_ ),
    .C1(\u_cpu.IMEM._0292_ ),
    .D1(\u_cpu.IMEM._0229_ ),
    .X(\u_cpu.IMEM._0293_ ));
 sky130_fd_sc_hd__or4b_2 \u_cpu.IMEM._1288_  (.A(\u_cpu.IMEM._0889_ ),
    .B(\u_cpu.IMEM._0184_ ),
    .C(\u_cpu.IMEM._0051_ ),
    .D_N(\u_cpu.IMEM._0075_ ),
    .X(\u_cpu.IMEM._0294_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1289_  (.A1(\u_cpu.IMEM._0294_ ),
    .A2(\u_cpu.IMEM._0292_ ),
    .B1(\u_cpu.IMEM._0237_ ),
    .Y(\u_cpu.IMEM._0296_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1290_  (.A1(\u_cpu.IMEM._0049_ ),
    .A2(\u_cpu.IMEM._0086_ ),
    .B1(\u_cpu.IMEM._0238_ ),
    .Y(\u_cpu.IMEM._0297_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1291_  (.A(\u_cpu.IMEM._0291_ ),
    .X(\u_cpu.IMEM._0298_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.IMEM._1292_  (.A1_N(\u_cpu.IMEM._0899_ ),
    .A2_N(\u_cpu.IMEM._0297_ ),
    .B1(\u_cpu.IMEM._0167_ ),
    .B2(\u_cpu.IMEM._0298_ ),
    .Y(\u_cpu.IMEM._0299_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.IMEM._1293_  (.A1(\u_cpu.IMEM._0009_ ),
    .A2(\u_cpu.IMEM._0190_ ),
    .B1(\u_cpu.IMEM._0008_ ),
    .C1(\u_cpu.IMEM._0120_ ),
    .X(\u_cpu.IMEM._0300_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1294_  (.A1(\u_cpu.IMEM._0615_ ),
    .A2(\u_cpu.IMEM._0299_ ),
    .B1(\u_cpu.IMEM._0300_ ),
    .C1(\u_cpu.IMEM._0699_ ),
    .X(\u_cpu.IMEM._0301_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1295_  (.A(\u_cpu.IMEM._0109_ ),
    .X(\u_cpu.IMEM._0302_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1296_  (.A1(\u_cpu.IMEM._0199_ ),
    .A2(\u_cpu.IMEM._0293_ ),
    .A3(\u_cpu.IMEM._0296_ ),
    .B1(\u_cpu.IMEM._0301_ ),
    .C1(\u_cpu.IMEM._0302_ ),
    .X(\u_cpu.IMEM._0303_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1297_  (.A1(\u_cpu.IMEM._0290_ ),
    .A2(\u_cpu.IMEM._0303_ ),
    .B1(\u_cpu.IMEM._0246_ ),
    .Y(\u_cpu.IMEM._0304_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1298_  (.A1(\u_cpu.IMEM._0108_ ),
    .A2(\u_cpu.IMEM._0279_ ),
    .B1(\u_cpu.IMEM._0304_ ),
    .Y(\u_cpu.IMEM.rd[7] ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1299_  (.A(\u_cpu.IMEM._0295_ ),
    .X(\u_cpu.IMEM._0306_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1300_  (.A(\u_cpu.IMEM._0112_ ),
    .X(\u_cpu.IMEM._0307_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1301_  (.A1(\u_cpu.IMEM._0307_ ),
    .A2(\u_cpu.IMEM._0138_ ),
    .B1(\u_cpu.IMEM._0093_ ),
    .Y(\u_cpu.IMEM._0308_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1302_  (.A(\u_cpu.IMEM._0059_ ),
    .X(\u_cpu.IMEM._0309_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1303_  (.A1(\u_cpu.IMEM._0309_ ),
    .A2(\u_cpu.IMEM._0101_ ),
    .B1(\u_cpu.IMEM._0099_ ),
    .Y(\u_cpu.IMEM._0310_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1304_  (.A1(\u_cpu.IMEM._0086_ ),
    .A2(\u_cpu.IMEM._0083_ ),
    .B1(\u_cpu.IMEM._0205_ ),
    .C1(\u_cpu.IMEM._0011_ ),
    .X(\u_cpu.IMEM._0311_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1305_  (.A1(\u_cpu.IMEM._0061_ ),
    .A2(\u_cpu.IMEM._0190_ ),
    .A3(\u_cpu.IMEM._0088_ ),
    .B1(\u_cpu.IMEM._0604_ ),
    .X(\u_cpu.IMEM._0312_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1306_  (.A1(\u_cpu.IMEM._0168_ ),
    .A2(\u_cpu.IMEM._0311_ ),
    .B1(\u_cpu.IMEM._0312_ ),
    .Y(\u_cpu.IMEM._0313_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.IMEM._1307_  (.A1(\u_cpu.IMEM._0308_ ),
    .A2(\u_cpu.IMEM._0310_ ),
    .B1(\u_cpu.IMEM._0090_ ),
    .C1(\u_cpu.IMEM._0313_ ),
    .X(\u_cpu.IMEM._0314_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1308_  (.A(\u_cpu.IMEM._0594_ ),
    .B(\u_cpu.IMEM._0889_ ),
    .Y(\u_cpu.IMEM._0315_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1309_  (.A1(\u_cpu.IMEM._0165_ ),
    .A2(\u_cpu.IMEM._0013_ ),
    .B1(\u_cpu.IMEM._0298_ ),
    .Y(\u_cpu.IMEM._0317_ ));
 sky130_fd_sc_hd__nor4b_2 \u_cpu.IMEM._1310_  (.A(\u_cpu.IMEM._0889_ ),
    .B(\u_cpu.IMEM._0184_ ),
    .C(\u_cpu.IMEM._0024_ ),
    .D_N(\u_cpu.IMEM._0927_ ),
    .Y(\u_cpu.IMEM._0318_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.IMEM._1311_  (.A_N(\u_cpu.IMEM._0034_ ),
    .B(\u_cpu.IMEM._0626_ ),
    .C(\u_cpu.IMEM._0424_ ),
    .D(\u_cpu.IMEM._0509_ ),
    .X(\u_cpu.IMEM._0319_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1312_  (.A1(\u_cpu.IMEM._0318_ ),
    .A2(\u_cpu.IMEM._0319_ ),
    .B1(\u_cpu.IMEM._0093_ ),
    .Y(\u_cpu.IMEM._0320_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1313_  (.A1(\u_cpu.IMEM._0315_ ),
    .A2(\u_cpu.IMEM._0317_ ),
    .B1(\u_cpu.IMEM._0320_ ),
    .Y(\u_cpu.IMEM._0321_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu.IMEM._1314_  (.A(\u_cpu.IMEM._0077_ ),
    .B(\u_cpu.IMEM._0321_ ),
    .X(\u_cpu.IMEM._0322_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1315_  (.A(\u_cpu.IMEM._0152_ ),
    .X(\u_cpu.IMEM._0323_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1316_  (.A1(\u_cpu.IMEM._0017_ ),
    .A2(\u_cpu.IMEM._0149_ ),
    .B1(\u_cpu.IMEM._0742_ ),
    .Y(\u_cpu.IMEM._0324_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.IMEM._1317_  (.A1(\u_cpu.IMEM._0309_ ),
    .A2(\u_cpu.IMEM._0323_ ),
    .B1(\u_cpu.IMEM._0119_ ),
    .C1(\u_cpu.IMEM._0225_ ),
    .D1(\u_cpu.IMEM._0324_ ),
    .Y(\u_cpu.IMEM._0325_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1318_  (.A1(\u_cpu.IMEM._0060_ ),
    .A2(\u_cpu.IMEM._0049_ ),
    .A3(\u_cpu.IMEM._0238_ ),
    .B1(\u_cpu.IMEM._0753_ ),
    .X(\u_cpu.IMEM._0326_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1319_  (.A1(\u_cpu.IMEM._0257_ ),
    .A2(\u_cpu.IMEM._0466_ ),
    .B1(\u_cpu.IMEM._0731_ ),
    .C1(\u_cpu.IMEM._0326_ ),
    .X(\u_cpu.IMEM._0328_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1320_  (.A1(\u_cpu.IMEM._0216_ ),
    .A2(\u_cpu.IMEM._0185_ ),
    .A3(\u_cpu.IMEM._0763_ ),
    .B1(\u_cpu.IMEM._0129_ ),
    .X(\u_cpu.IMEM._0329_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.IMEM._1321_  (.A1(\u_cpu.IMEM._0710_ ),
    .A2(\u_cpu.IMEM._0325_ ),
    .A3(\u_cpu.IMEM._0328_ ),
    .B1(\u_cpu.IMEM._0329_ ),
    .Y(\u_cpu.IMEM._0330_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1322_  (.A(\u_cpu.IMEM._0134_ ),
    .B(\u_cpu.IMEM._0657_ ),
    .Y(\u_cpu.IMEM._0331_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1323_  (.A1(\u_cpu.IMEM._0040_ ),
    .A2(\u_cpu.IMEM._0152_ ),
    .B1(\u_cpu.IMEM._0217_ ),
    .Y(\u_cpu.IMEM._0332_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1324_  (.A(\u_cpu.IMEM.a[8] ),
    .X(\u_cpu.IMEM._0333_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1325_  (.A1(\u_cpu.IMEM._0331_ ),
    .A2(\u_cpu.IMEM._0332_ ),
    .B1(\u_cpu.IMEM._0333_ ),
    .Y(\u_cpu.IMEM._0334_ ));
 sky130_fd_sc_hd__o32ai_2 \u_cpu.IMEM._1326_  (.A1(\u_cpu.IMEM._0306_ ),
    .A2(\u_cpu.IMEM._0314_ ),
    .A3(\u_cpu.IMEM._0322_ ),
    .B1(\u_cpu.IMEM._0330_ ),
    .B2(\u_cpu.IMEM._0334_ ),
    .Y(\u_cpu.IMEM._0335_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1327_  (.A1(\u_cpu.IMEM._0294_ ),
    .A2(\u_cpu.IMEM._0212_ ),
    .B1(\u_cpu.IMEM._0129_ ),
    .Y(\u_cpu.IMEM._0336_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1328_  (.A1(\u_cpu.IMEM._0075_ ),
    .A2(\u_cpu.IMEM._0051_ ),
    .B1(\u_cpu.IMEM._0189_ ),
    .Y(\u_cpu.IMEM._0337_ ));
 sky130_fd_sc_hd__and4bb_2 \u_cpu.IMEM._1329_  (.A_N(\u_cpu.IMEM._0424_ ),
    .B_N(\u_cpu.IMEM._0927_ ),
    .C(\u_cpu.IMEM._0034_ ),
    .D(\u_cpu.IMEM._0012_ ),
    .X(\u_cpu.IMEM._0339_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1330_  (.A1(\u_cpu.IMEM._0337_ ),
    .A2(\u_cpu.IMEM._0080_ ),
    .B1(\u_cpu.IMEM._0339_ ),
    .Y(\u_cpu.IMEM._0340_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.IMEM._1331_  (.A(\u_cpu.IMEM._0021_ ),
    .B(\u_cpu.IMEM._0184_ ),
    .C(\u_cpu.IMEM._0024_ ),
    .X(\u_cpu.IMEM._0341_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.IMEM._1332_  (.A1(\u_cpu.IMEM._0101_ ),
    .A2(\u_cpu.IMEM._0044_ ),
    .A3(\u_cpu.IMEM._0920_ ),
    .B1(\u_cpu.IMEM._0341_ ),
    .Y(\u_cpu.IMEM._0342_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.IMEM._1333_  (.A1(\u_cpu.IMEM._0340_ ),
    .A2(\u_cpu.IMEM._0272_ ),
    .B1(\u_cpu.IMEM._0268_ ),
    .B2(\u_cpu.IMEM._0342_ ),
    .Y(\u_cpu.IMEM._0343_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1334_  (.A1(\u_cpu.IMEM._0170_ ),
    .A2(\u_cpu.IMEM._0336_ ),
    .B1(\u_cpu.IMEM._0343_ ),
    .Y(\u_cpu.IMEM._0344_ ));
 sky130_fd_sc_hd__nor4_2 \u_cpu.IMEM._1335_  (.A(\u_cpu.IMEM._0082_ ),
    .B(\u_cpu.IMEM._0636_ ),
    .C(\u_cpu.IMEM._0032_ ),
    .D(\u_cpu.IMEM._0879_ ),
    .Y(\u_cpu.IMEM._0345_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.IMEM._1336_  (.A1(\u_cpu.IMEM._0257_ ),
    .A2(\u_cpu.IMEM._0119_ ),
    .B1(\u_cpu.IMEM._0332_ ),
    .B2(\u_cpu.IMEM._0345_ ),
    .Y(\u_cpu.IMEM._0346_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1337_  (.A1(\u_cpu.IMEM._0034_ ),
    .A2(\u_cpu.IMEM._0795_ ),
    .B1(\u_cpu.IMEM._0112_ ),
    .Y(\u_cpu.IMEM._0347_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.IMEM._1338_  (.A1(\u_cpu.IMEM._0033_ ),
    .A2(\u_cpu.IMEM._0251_ ),
    .B1(\u_cpu.IMEM._0236_ ),
    .C1(\u_cpu.IMEM._0347_ ),
    .X(\u_cpu.IMEM._0348_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.IMEM._1339_  (.A1(\u_cpu.IMEM._0346_ ),
    .A2(\u_cpu.IMEM._0094_ ),
    .B1(\u_cpu.IMEM._0348_ ),
    .C1(\u_cpu.IMEM._0186_ ),
    .Y(\u_cpu.IMEM._0350_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1340_  (.A(\u_cpu.IMEM.a[8] ),
    .B(\u_cpu.IMEM._0667_ ),
    .Y(\u_cpu.IMEM._0351_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.IMEM._1341_  (.A1(\u_cpu.IMEM._0763_ ),
    .A2(\u_cpu.IMEM._0197_ ),
    .A3(\u_cpu.IMEM._0166_ ),
    .B1(\u_cpu.IMEM._0089_ ),
    .C1(\u_cpu.IMEM._0225_ ),
    .Y(\u_cpu.IMEM._0352_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1342_  (.A1(\u_cpu.IMEM._0086_ ),
    .A2(\u_cpu.IMEM._0238_ ),
    .B1(\u_cpu.IMEM._0009_ ),
    .Y(\u_cpu.IMEM._0353_ ));
 sky130_fd_sc_hd__or3b_2 \u_cpu.IMEM._1343_  (.A(\u_cpu.IMEM._0353_ ),
    .B(\u_cpu.IMEM._0236_ ),
    .C_N(\u_cpu.IMEM._0120_ ),
    .X(\u_cpu.IMEM._0354_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.IMEM._1344_  (.A(\u_cpu.IMEM._0129_ ),
    .B(\u_cpu.IMEM._0109_ ),
    .Y(\u_cpu.IMEM._0355_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.IMEM._1345_  (.A1(\u_cpu.IMEM._0352_ ),
    .A2(\u_cpu.IMEM._0354_ ),
    .A3(\u_cpu.IMEM._0355_ ),
    .B1(\u_cpu.IMEM.a[9] ),
    .Y(\u_cpu.IMEM._0356_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.IMEM._1346_  (.A1(\u_cpu.IMEM._0194_ ),
    .A2(\u_cpu.IMEM._0344_ ),
    .B1(\u_cpu.IMEM._0350_ ),
    .B2(\u_cpu.IMEM._0351_ ),
    .C1(\u_cpu.IMEM._0356_ ),
    .X(\u_cpu.IMEM._0357_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1347_  (.A1(\u_cpu.IMEM._0108_ ),
    .A2(\u_cpu.IMEM._0335_ ),
    .B1(\u_cpu.IMEM._0357_ ),
    .Y(\u_cpu.IMEM.rd[8] ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1348_  (.A1(\u_cpu.IMEM._0030_ ),
    .A2(\u_cpu.IMEM._0148_ ),
    .B1(\u_cpu.IMEM._0044_ ),
    .Y(\u_cpu.IMEM._0358_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.IMEM._1349_  (.A(\u_cpu.IMEM._0868_ ),
    .B(\u_cpu.IMEM._0848_ ),
    .C(\u_cpu.IMEM._0032_ ),
    .Y(\u_cpu.IMEM._0360_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.IMEM._1350_  (.A(\u_cpu.IMEM._0191_ ),
    .B(\u_cpu.IMEM._0165_ ),
    .C(\u_cpu.IMEM._0014_ ),
    .D(\u_cpu.IMEM._0040_ ),
    .Y(\u_cpu.IMEM._0361_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1351_  (.A1(\u_cpu.IMEM._0358_ ),
    .A2(\u_cpu.IMEM._0360_ ),
    .B1(\u_cpu.IMEM._0294_ ),
    .C1(\u_cpu.IMEM._0361_ ),
    .Y(\u_cpu.IMEM._0362_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.IMEM._1352_  (.A(\u_cpu.IMEM._0359_ ),
    .B(\u_cpu.IMEM._0392_ ),
    .C(\u_cpu.IMEM._0012_ ),
    .Y(\u_cpu.IMEM._0363_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1353_  (.A(\u_cpu.IMEM._0032_ ),
    .B(\u_cpu.IMEM._0059_ ),
    .Y(\u_cpu.IMEM._0364_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1354_  (.A1(\u_cpu.IMEM._0283_ ),
    .A2(\u_cpu.IMEM._0082_ ),
    .A3(\u_cpu.IMEM._0008_ ),
    .B1(\u_cpu.IMEM.a[7] ),
    .X(\u_cpu.IMEM._0365_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1355_  (.A1(\u_cpu.IMEM._0163_ ),
    .A2(\u_cpu.IMEM._0363_ ),
    .A3(\u_cpu.IMEM._0364_ ),
    .B1(\u_cpu.IMEM._0365_ ),
    .X(\u_cpu.IMEM._0366_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1356_  (.A1(\u_cpu.IMEM._0145_ ),
    .A2(\u_cpu.IMEM._0362_ ),
    .B1(\u_cpu.IMEM._0366_ ),
    .Y(\u_cpu.IMEM._0367_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.IMEM._1357_  (.A(\u_cpu.IMEM._0134_ ),
    .B(\u_cpu.IMEM._0088_ ),
    .C(\u_cpu.IMEM._0298_ ),
    .X(\u_cpu.IMEM._0368_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1358_  (.A1(\u_cpu.IMEM._0187_ ),
    .A2(\u_cpu.IMEM._0138_ ),
    .A3(\u_cpu.IMEM._0217_ ),
    .B1(\u_cpu.IMEM._0003_ ),
    .X(\u_cpu.IMEM._0369_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1359_  (.A(\u_cpu.IMEM._0392_ ),
    .X(\u_cpu.IMEM._0371_ ));
 sky130_fd_sc_hd__a311o_2 \u_cpu.IMEM._1360_  (.A1(\u_cpu.IMEM._0920_ ),
    .A2(\u_cpu.IMEM._0078_ ),
    .A3(\u_cpu.IMEM._0371_ ),
    .B1(\u_cpu.IMEM._0180_ ),
    .C1(\u_cpu.IMEM._0096_ ),
    .X(\u_cpu.IMEM._0372_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1361_  (.A1(\u_cpu.IMEM._0000_ ),
    .A2(\u_cpu.IMEM._0042_ ),
    .B1(\u_cpu.IMEM._0176_ ),
    .Y(\u_cpu.IMEM._0373_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1362_  (.A1(\u_cpu.IMEM._0763_ ),
    .A2(\u_cpu.IMEM._0373_ ),
    .B1(\u_cpu.IMEM._0731_ ),
    .Y(\u_cpu.IMEM._0374_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.IMEM._1363_  (.A1(\u_cpu.IMEM._0368_ ),
    .A2(\u_cpu.IMEM._0369_ ),
    .B1(\u_cpu.IMEM._0372_ ),
    .B2(\u_cpu.IMEM._0374_ ),
    .C1(\u_cpu.IMEM._0077_ ),
    .Y(\u_cpu.IMEM._0375_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1364_  (.A1(\u_cpu.IMEM._0148_ ),
    .A2(\u_cpu.IMEM._0042_ ),
    .A3(\u_cpu.IMEM._0858_ ),
    .B1(\u_cpu.IMEM._0099_ ),
    .X(\u_cpu.IMEM._0376_ ));
 sky130_fd_sc_hd__nor2b_2 \u_cpu.IMEM._1365_  (.A(\u_cpu.IMEM._0519_ ),
    .B_N(\u_cpu.IMEM._0019_ ),
    .Y(\u_cpu.IMEM._0377_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.IMEM._1366_  (.A(\u_cpu.IMEM._0604_ ),
    .B(\u_cpu.IMEM._0879_ ),
    .C(\u_cpu.IMEM._0377_ ),
    .X(\u_cpu.IMEM._0378_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1367_  (.A1(\u_cpu.IMEM._0115_ ),
    .A2(\u_cpu.IMEM._0046_ ),
    .A3(\u_cpu.IMEM._0048_ ),
    .B1(\u_cpu.IMEM._0689_ ),
    .X(\u_cpu.IMEM._0379_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.IMEM._1368_  (.A1(\u_cpu.IMEM._0144_ ),
    .A2(\u_cpu.IMEM._0376_ ),
    .B1(\u_cpu.IMEM._0378_ ),
    .B2(\u_cpu.IMEM._0379_ ),
    .C1(\u_cpu.IMEM._0109_ ),
    .X(\u_cpu.IMEM._0380_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1369_  (.A1(\u_cpu.IMEM._0255_ ),
    .A2(\u_cpu.IMEM._0367_ ),
    .A3(\u_cpu.IMEM._0375_ ),
    .B1(\u_cpu.IMEM._0380_ ),
    .X(\u_cpu.IMEM._0382_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1370_  (.A1(\u_cpu.IMEM._0174_ ),
    .A2(\u_cpu.IMEM._0636_ ),
    .B1(\u_cpu.IMEM._0721_ ),
    .X(\u_cpu.IMEM._0383_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1371_  (.A1(\u_cpu.IMEM._0161_ ),
    .A2(\u_cpu.IMEM._0162_ ),
    .A3(\u_cpu.IMEM._0315_ ),
    .B1(\u_cpu.IMEM._0383_ ),
    .C1(\u_cpu.IMEM._0062_ ),
    .X(\u_cpu.IMEM._0384_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1372_  (.A1(\u_cpu.IMEM._0086_ ),
    .A2(\u_cpu.IMEM._0238_ ),
    .B1(\u_cpu.IMEM._0070_ ),
    .C1(\u_cpu.IMEM._0205_ ),
    .X(\u_cpu.IMEM._0385_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1373_  (.A1(\u_cpu.IMEM._0060_ ),
    .A2(\u_cpu.IMEM._0049_ ),
    .B1(\u_cpu.IMEM._0205_ ),
    .C1(\u_cpu.IMEM._0082_ ),
    .X(\u_cpu.IMEM._0386_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1374_  (.A1(\u_cpu.IMEM._0731_ ),
    .A2(\u_cpu.IMEM._0385_ ),
    .A3(\u_cpu.IMEM._0386_ ),
    .B1(\u_cpu.IMEM._0667_ ),
    .X(\u_cpu.IMEM._0387_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.IMEM._1375_  (.A(\u_cpu.IMEM._0920_ ),
    .B(\u_cpu.IMEM._0078_ ),
    .C(\u_cpu.IMEM._0371_ ),
    .D(\u_cpu.IMEM._0187_ ),
    .Y(\u_cpu.IMEM._0388_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.IMEM._1376_  (.A1(\u_cpu.IMEM._0189_ ),
    .A2(\u_cpu.IMEM._0169_ ),
    .A3(\u_cpu.IMEM._0388_ ),
    .B1(\u_cpu.IMEM._0237_ ),
    .Y(\u_cpu.IMEM._0389_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.IMEM._1377_  (.A1(\u_cpu.IMEM._0077_ ),
    .A2(\u_cpu.IMEM._0384_ ),
    .B1(\u_cpu.IMEM._0387_ ),
    .B2(\u_cpu.IMEM._0389_ ),
    .C1(\u_cpu.IMEM._0333_ ),
    .X(\u_cpu.IMEM._0390_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1378_  (.A1(\u_cpu.IMEM._0132_ ),
    .A2(\u_cpu.IMEM._0413_ ),
    .A3(\u_cpu.IMEM._0176_ ),
    .B1(\u_cpu.IMEM._0123_ ),
    .X(\u_cpu.IMEM._0391_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.IMEM._1379_  (.A1(\u_cpu.IMEM._0920_ ),
    .A2(\u_cpu.IMEM._0185_ ),
    .B1(\u_cpu.IMEM._0251_ ),
    .B2(\u_cpu.IMEM._0033_ ),
    .C1(\u_cpu.IMEM._0257_ ),
    .X(\u_cpu.IMEM._0393_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1380_  (.A1(\u_cpu.IMEM._0391_ ),
    .A2(\u_cpu.IMEM._0393_ ),
    .B1(\u_cpu.IMEM._0248_ ),
    .Y(\u_cpu.IMEM._0394_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.IMEM._1381_  (.A(\u_cpu.IMEM._0046_ ),
    .B(\u_cpu.IMEM._0187_ ),
    .Y(\u_cpu.IMEM._0395_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.IMEM._1382_  (.A(\u_cpu.IMEM._0007_ ),
    .B(\u_cpu.IMEM._0095_ ),
    .Y(\u_cpu.IMEM._0396_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.IMEM._1383_  (.A1(\u_cpu.IMEM._0466_ ),
    .A2(\u_cpu.IMEM._0498_ ),
    .A3(\u_cpu.IMEM._0395_ ),
    .B1(\u_cpu.IMEM._0396_ ),
    .B2(\u_cpu.IMEM._0197_ ),
    .X(\u_cpu.IMEM._0397_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1384_  (.A1(\u_cpu.IMEM._0858_ ),
    .A2(\u_cpu.IMEM._0323_ ),
    .B1(\u_cpu.IMEM._0118_ ),
    .C1(\u_cpu.IMEM._0096_ ),
    .Y(\u_cpu.IMEM._0398_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1385_  (.A1(\u_cpu.IMEM._0240_ ),
    .A2(\u_cpu.IMEM._0398_ ),
    .B1(\u_cpu.IMEM._0237_ ),
    .Y(\u_cpu.IMEM._0399_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1386_  (.A1(\u_cpu.IMEM._0397_ ),
    .A2(\u_cpu.IMEM._0399_ ),
    .B1(\u_cpu.IMEM._0028_ ),
    .Y(\u_cpu.IMEM._0400_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1387_  (.A1(\u_cpu.IMEM._0394_ ),
    .A2(\u_cpu.IMEM._0400_ ),
    .B1(\u_cpu.IMEM._0306_ ),
    .Y(\u_cpu.IMEM._0401_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.IMEM._1388_  (.A1(\u_cpu.IMEM._0390_ ),
    .A2(\u_cpu.IMEM._0401_ ),
    .B1_N(\u_cpu.IMEM._0055_ ),
    .Y(\u_cpu.IMEM._0402_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1389_  (.A1(\u_cpu.IMEM._0128_ ),
    .A2(\u_cpu.IMEM._0382_ ),
    .B1(\u_cpu.IMEM._0402_ ),
    .Y(\u_cpu.IMEM.rd[9] ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.IMEM._1390_  (.A1(\u_cpu.IMEM._0174_ ),
    .A2(\u_cpu.IMEM._0636_ ),
    .B1(\u_cpu.IMEM._0011_ ),
    .C1(\u_cpu.IMEM._0189_ ),
    .X(\u_cpu.IMEM._0404_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1391_  (.A1(\u_cpu.IMEM._0165_ ),
    .A2(\u_cpu.IMEM._0014_ ),
    .B1(\u_cpu.IMEM._0030_ ),
    .C1(\u_cpu.IMEM._0315_ ),
    .X(\u_cpu.IMEM._0405_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1392_  (.A1(\u_cpu.IMEM._0731_ ),
    .A2(\u_cpu.IMEM._0326_ ),
    .A3(\u_cpu.IMEM._0404_ ),
    .B1(\u_cpu.IMEM._0129_ ),
    .C1(\u_cpu.IMEM._0405_ ),
    .X(\u_cpu.IMEM._0406_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1393_  (.A(\u_cpu.IMEM._0174_ ),
    .B(\u_cpu.IMEM._0205_ ),
    .Y(\u_cpu.IMEM._0407_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1394_  (.A1(\u_cpu.IMEM._0466_ ),
    .A2(\u_cpu.IMEM._0049_ ),
    .B1(\u_cpu.IMEM._0070_ ),
    .C1(\u_cpu.IMEM._0879_ ),
    .X(\u_cpu.IMEM._0408_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.IMEM._1395_  (.A1(\u_cpu.IMEM._0044_ ),
    .A2(\u_cpu.IMEM._0088_ ),
    .A3(\u_cpu.IMEM._0101_ ),
    .B1(\u_cpu.IMEM._0229_ ),
    .C1(\u_cpu.IMEM._0408_ ),
    .Y(\u_cpu.IMEM._0409_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1396_  (.A1(\u_cpu.IMEM._0615_ ),
    .A2(\u_cpu.IMEM._0407_ ),
    .A3(\u_cpu.IMEM._0188_ ),
    .B1(\u_cpu.IMEM._0699_ ),
    .C1(\u_cpu.IMEM._0409_ ),
    .X(\u_cpu.IMEM._0410_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1397_  (.A(\u_cpu.IMEM._0022_ ),
    .X(\u_cpu.IMEM._0411_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1398_  (.A1(\u_cpu.IMEM._0030_ ),
    .A2(\u_cpu.IMEM._0411_ ),
    .B1(\u_cpu.IMEM._0307_ ),
    .Y(\u_cpu.IMEM._0412_ ));
 sky130_fd_sc_hd__o32ai_2 \u_cpu.IMEM._1399_  (.A1(\u_cpu.IMEM._0298_ ),
    .A2(\u_cpu.IMEM._0763_ ),
    .A3(\u_cpu.IMEM._0161_ ),
    .B1(\u_cpu.IMEM._0412_ ),
    .B2(\u_cpu.IMEM._0251_ ),
    .Y(\u_cpu.IMEM._0414_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1400_  (.A(\u_cpu.IMEM._0816_ ),
    .X(\u_cpu.IMEM._0415_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.IMEM._1401_  (.A1(\u_cpu.IMEM._0646_ ),
    .A2(\u_cpu.IMEM._0415_ ),
    .B1(\u_cpu.IMEM._0048_ ),
    .C1(\u_cpu.IMEM._0396_ ),
    .X(\u_cpu.IMEM._0416_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.IMEM._1402_  (.A1(\u_cpu.IMEM._0414_ ),
    .A2(\u_cpu.IMEM._0124_ ),
    .B1(\u_cpu.IMEM._0125_ ),
    .C1(\u_cpu.IMEM._0416_ ),
    .Y(\u_cpu.IMEM._0417_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.IMEM._1403_  (.A(\u_cpu.IMEM._0218_ ),
    .B(\u_cpu.IMEM._0251_ ),
    .C(\u_cpu.IMEM._0096_ ),
    .D(\u_cpu.IMEM._0157_ ),
    .X(\u_cpu.IMEM._0418_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1404_  (.A1(\u_cpu.IMEM._0197_ ),
    .A2(\u_cpu.IMEM._0003_ ),
    .A3(\u_cpu.IMEM._0230_ ),
    .B1(\u_cpu.IMEM._0066_ ),
    .X(\u_cpu.IMEM._0419_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1405_  (.A1(\u_cpu.IMEM._0418_ ),
    .A2(\u_cpu.IMEM._0419_ ),
    .B1(\u_cpu.IMEM._0333_ ),
    .Y(\u_cpu.IMEM._0420_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.IMEM._1406_  (.A1(\u_cpu.IMEM._0255_ ),
    .A2(\u_cpu.IMEM._0406_ ),
    .A3(\u_cpu.IMEM._0410_ ),
    .B1(\u_cpu.IMEM._0417_ ),
    .B2(\u_cpu.IMEM._0420_ ),
    .X(\u_cpu.IMEM._0421_ ));
 sky130_fd_sc_hd__or4_2 \u_cpu.IMEM._1407_  (.A(\u_cpu.IMEM._0604_ ),
    .B(\u_cpu.IMEM._0217_ ),
    .C(\u_cpu.IMEM._0191_ ),
    .D(\u_cpu.IMEM._0323_ ),
    .X(\u_cpu.IMEM._0422_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1408_  (.A1(\u_cpu.IMEM._0094_ ),
    .A2(\u_cpu.IMEM._0135_ ),
    .A3(\u_cpu.IMEM._0310_ ),
    .B1(\u_cpu.IMEM._0422_ ),
    .C1(\u_cpu.IMEM._0125_ ),
    .X(\u_cpu.IMEM._0423_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.IMEM._1409_  (.A(\u_cpu.IMEM._0742_ ),
    .B(\u_cpu.IMEM._0509_ ),
    .C(\u_cpu.IMEM._0034_ ),
    .D(\u_cpu.IMEM._0012_ ),
    .Y(\u_cpu.IMEM._0425_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1410_  (.A1(\u_cpu.IMEM._0425_ ),
    .A2(\u_cpu.IMEM._0120_ ),
    .B1(\u_cpu.IMEM._0721_ ),
    .X(\u_cpu.IMEM._0426_ ));
 sky130_fd_sc_hd__o41a_2 \u_cpu.IMEM._1411_  (.A1(\u_cpu.IMEM._0038_ ),
    .A2(\u_cpu.IMEM._0064_ ),
    .A3(\u_cpu.IMEM._0185_ ),
    .A4(\u_cpu.IMEM._0231_ ),
    .B1(\u_cpu.IMEM._0426_ ),
    .X(\u_cpu.IMEM._0427_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1412_  (.A1(\u_cpu.IMEM._0258_ ),
    .A2(\u_cpu.IMEM._0281_ ),
    .B1(\u_cpu.IMEM._0318_ ),
    .C1(\u_cpu.IMEM._0066_ ),
    .X(\u_cpu.IMEM._0428_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.IMEM._1413_  (.A(\u_cpu.IMEM._0281_ ),
    .B(\u_cpu.IMEM._0258_ ),
    .Y(\u_cpu.IMEM._0429_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.IMEM._1414_  (.A1_N(\u_cpu.IMEM._0199_ ),
    .A2_N(\u_cpu.IMEM._0427_ ),
    .B1(\u_cpu.IMEM._0428_ ),
    .B2(\u_cpu.IMEM._0429_ ),
    .X(\u_cpu.IMEM._0430_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1415_  (.A(\u_cpu.IMEM.a[9] ),
    .X(\u_cpu.IMEM._0431_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.IMEM._1416_  (.A1(\u_cpu.IMEM._0423_ ),
    .A2(\u_cpu.IMEM._0334_ ),
    .B1(\u_cpu.IMEM._0305_ ),
    .B2(\u_cpu.IMEM._0430_ ),
    .C1(\u_cpu.IMEM._0431_ ),
    .Y(\u_cpu.IMEM._0432_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1417_  (.A1(\u_cpu.IMEM._0108_ ),
    .A2(\u_cpu.IMEM._0421_ ),
    .B1(\u_cpu.IMEM._0432_ ),
    .Y(\u_cpu.IMEM.rd[10] ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1418_  (.A1(\u_cpu.IMEM._0858_ ),
    .A2(\u_cpu.IMEM._0042_ ),
    .B1(\u_cpu.IMEM._0191_ ),
    .C1(\u_cpu.IMEM._0498_ ),
    .Y(\u_cpu.IMEM._0433_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1419_  (.A(\u_cpu.IMEM._0038_ ),
    .X(\u_cpu.IMEM._0435_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1420_  (.A1(\u_cpu.IMEM._0121_ ),
    .A2(\u_cpu.IMEM._0030_ ),
    .A3(\u_cpu.IMEM._0080_ ),
    .B1(\u_cpu.IMEM._0066_ ),
    .X(\u_cpu.IMEM._0436_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.IMEM._1421_  (.A1(\u_cpu.IMEM._0101_ ),
    .A2(\u_cpu.IMEM._0188_ ),
    .B1(\u_cpu.IMEM._0435_ ),
    .C1(\u_cpu.IMEM._0436_ ),
    .Y(\u_cpu.IMEM._0437_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.IMEM._1422_  (.A(\u_cpu.IMEM._0487_ ),
    .B(\u_cpu.IMEM._0785_ ),
    .X(\u_cpu.IMEM._0438_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1423_  (.A(\u_cpu.IMEM._0438_ ),
    .X(\u_cpu.IMEM._0439_ ));
 sky130_fd_sc_hd__or4_2 \u_cpu.IMEM._1424_  (.A(\u_cpu.IMEM._0007_ ),
    .B(\u_cpu.IMEM._0024_ ),
    .C(\u_cpu.IMEM._0816_ ),
    .D(\u_cpu.IMEM._0095_ ),
    .X(\u_cpu.IMEM._0440_ ));
 sky130_fd_sc_hd__o41ai_2 \u_cpu.IMEM._1425_  (.A1(\u_cpu.IMEM._0229_ ),
    .A2(\u_cpu.IMEM._0257_ ),
    .A3(\u_cpu.IMEM._0216_ ),
    .A4(\u_cpu.IMEM._0439_ ),
    .B1(\u_cpu.IMEM._0440_ ),
    .Y(\u_cpu.IMEM._0441_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.IMEM._1426_  (.A1(\u_cpu.IMEM._0433_ ),
    .A2(\u_cpu.IMEM._0437_ ),
    .B1(\u_cpu.IMEM._0441_ ),
    .B2(\u_cpu.IMEM._0173_ ),
    .C1(\u_cpu.IMEM._0194_ ),
    .Y(\u_cpu.IMEM._0442_ ));
 sky130_fd_sc_hd__or4_2 \u_cpu.IMEM._1427_  (.A(\u_cpu.IMEM._0230_ ),
    .B(\u_cpu.IMEM._0157_ ),
    .C(\u_cpu.IMEM._0415_ ),
    .D(\u_cpu.IMEM._0272_ ),
    .X(\u_cpu.IMEM._0443_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1428_  (.A1(\u_cpu.IMEM._0228_ ),
    .A2(\u_cpu.IMEM._0119_ ),
    .A3(\u_cpu.IMEM._0039_ ),
    .B1(\u_cpu.IMEM._0333_ ),
    .C1(\u_cpu.IMEM._0443_ ),
    .X(\u_cpu.IMEM._0444_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1429_  (.A1(\u_cpu.IMEM._0075_ ),
    .A2(\u_cpu.IMEM._0023_ ),
    .B1(\u_cpu.IMEM._0051_ ),
    .Y(\u_cpu.IMEM._0446_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1430_  (.A(\u_cpu.IMEM._0038_ ),
    .X(\u_cpu.IMEM._0447_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.IMEM._1431_  (.A1(\u_cpu.IMEM._0060_ ),
    .A2(\u_cpu.IMEM._0205_ ),
    .B1(\u_cpu.IMEM._0014_ ),
    .B2(\u_cpu.IMEM._0636_ ),
    .C1(\u_cpu.IMEM._0011_ ),
    .Y(\u_cpu.IMEM._0448_ ));
 sky130_fd_sc_hd__a311oi_2 \u_cpu.IMEM._1432_  (.A1(\u_cpu.IMEM._0119_ ),
    .A2(\u_cpu.IMEM._0324_ ),
    .A3(\u_cpu.IMEM._0446_ ),
    .B1(\u_cpu.IMEM._0447_ ),
    .C1(\u_cpu.IMEM._0448_ ),
    .Y(\u_cpu.IMEM._0449_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1433_  (.A1(\u_cpu.IMEM._0060_ ),
    .A2(\u_cpu.IMEM._0238_ ),
    .B1(\u_cpu.IMEM._0061_ ),
    .X(\u_cpu.IMEM._0450_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1434_  (.A1(\u_cpu.IMEM._0251_ ),
    .A2(\u_cpu.IMEM._0041_ ),
    .A3(\u_cpu.IMEM._0450_ ),
    .B1(\u_cpu.IMEM._0150_ ),
    .C1(\u_cpu.IMEM._0262_ ),
    .X(\u_cpu.IMEM._0451_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.IMEM._1435_  (.A(\u_cpu.IMEM._0103_ ),
    .B(\u_cpu.IMEM._0445_ ),
    .C(\u_cpu.IMEM._0332_ ),
    .X(\u_cpu.IMEM._0452_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1436_  (.A1(\u_cpu.IMEM._0208_ ),
    .A2(\u_cpu.IMEM._0449_ ),
    .A3(\u_cpu.IMEM._0451_ ),
    .B1(\u_cpu.IMEM._0452_ ),
    .C1(\u_cpu.IMEM._0194_ ),
    .X(\u_cpu.IMEM._0453_ ));
 sky130_fd_sc_hd__or4_2 \u_cpu.IMEM._1437_  (.A(\u_cpu.IMEM._0015_ ),
    .B(\u_cpu.IMEM._0115_ ),
    .C(\u_cpu.IMEM._0000_ ),
    .D(\u_cpu.IMEM._0411_ ),
    .X(\u_cpu.IMEM._0454_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1438_  (.A1(\u_cpu.IMEM._0040_ ),
    .A2(\u_cpu.IMEM._0323_ ),
    .B1(\u_cpu.IMEM._0347_ ),
    .Y(\u_cpu.IMEM._0455_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1439_  (.A1(\u_cpu.IMEM._0361_ ),
    .A2(\u_cpu.IMEM._0455_ ),
    .B1(\u_cpu.IMEM._0615_ ),
    .X(\u_cpu.IMEM._0457_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1440_  (.A1(\u_cpu.IMEM._0454_ ),
    .A2(\u_cpu.IMEM._0457_ ),
    .B1(\u_cpu.IMEM._0208_ ),
    .Y(\u_cpu.IMEM._0458_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.IMEM._1441_  (.A1(\u_cpu.IMEM._0184_ ),
    .A2(\u_cpu.IMEM._0024_ ),
    .B1(\u_cpu.IMEM._0466_ ),
    .C1(\u_cpu.IMEM._0095_ ),
    .X(\u_cpu.IMEM._0459_ ));
 sky130_fd_sc_hd__a32oi_2 \u_cpu.IMEM._1442_  (.A1(\u_cpu.IMEM._0324_ ),
    .A2(\u_cpu.IMEM._0446_ ),
    .A3(\u_cpu.IMEM._0119_ ),
    .B1(\u_cpu.IMEM._0459_ ),
    .B2(\u_cpu.IMEM._0176_ ),
    .Y(\u_cpu.IMEM._0460_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.IMEM._1443_  (.A1(\u_cpu.IMEM._0369_ ),
    .A2(\u_cpu.IMEM._0455_ ),
    .B1(\u_cpu.IMEM._0460_ ),
    .B2(\u_cpu.IMEM._0131_ ),
    .C1(\u_cpu.IMEM._0125_ ),
    .Y(\u_cpu.IMEM._0461_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.IMEM._1444_  (.A1(\u_cpu.IMEM._0306_ ),
    .A2(\u_cpu.IMEM._0458_ ),
    .A3(\u_cpu.IMEM._0461_ ),
    .B1(\u_cpu.IMEM._0316_ ),
    .Y(\u_cpu.IMEM._0462_ ));
 sky130_fd_sc_hd__o32ai_2 \u_cpu.IMEM._1445_  (.A1(\u_cpu.IMEM._0431_ ),
    .A2(\u_cpu.IMEM._0442_ ),
    .A3(\u_cpu.IMEM._0444_ ),
    .B1(\u_cpu.IMEM._0453_ ),
    .B2(\u_cpu.IMEM._0462_ ),
    .Y(\u_cpu.IMEM.rd[11] ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.IMEM._1446_  (.A(\u_cpu.IMEM._0594_ ),
    .B(\u_cpu.IMEM._0021_ ),
    .C(\u_cpu.IMEM._0023_ ),
    .D(\u_cpu.IMEM._0795_ ),
    .Y(\u_cpu.IMEM._0463_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.IMEM._1447_  (.A1_N(\u_cpu.IMEM._0434_ ),
    .A2_N(\u_cpu.IMEM._0463_ ),
    .B1(\u_cpu.IMEM._0161_ ),
    .B2(\u_cpu.IMEM._0285_ ),
    .X(\u_cpu.IMEM._0464_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1448_  (.A1(\u_cpu.IMEM._0434_ ),
    .A2(\u_cpu.IMEM._0013_ ),
    .A3(\u_cpu.IMEM._0415_ ),
    .B1(\u_cpu.IMEM._0236_ ),
    .X(\u_cpu.IMEM._0465_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1449_  (.A1(\u_cpu.IMEM._0153_ ),
    .A2(\u_cpu.IMEM._0262_ ),
    .B1(\u_cpu.IMEM._0465_ ),
    .Y(\u_cpu.IMEM._0467_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.IMEM._1450_  (.A1(\u_cpu.IMEM._0419_ ),
    .A2(\u_cpu.IMEM._0464_ ),
    .B1(\u_cpu.IMEM._0467_ ),
    .B2(\u_cpu.IMEM._0125_ ),
    .X(\u_cpu.IMEM._0468_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1451_  (.A(\u_cpu.IMEM._0109_ ),
    .X(\u_cpu.IMEM._0469_ ));
 sky130_fd_sc_hd__o41a_2 \u_cpu.IMEM._1452_  (.A1(\u_cpu.IMEM._0009_ ),
    .A2(\u_cpu.IMEM._0086_ ),
    .A3(\u_cpu.IMEM._0176_ ),
    .A4(\u_cpu.IMEM._0721_ ),
    .B1(\u_cpu.IMEM._0689_ ),
    .X(\u_cpu.IMEM._0470_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1453_  (.A1(\u_cpu.IMEM._0002_ ),
    .A2(\u_cpu.IMEM._0142_ ),
    .B1(\u_cpu.IMEM._0035_ ),
    .C1(\u_cpu.IMEM._0229_ ),
    .Y(\u_cpu.IMEM._0471_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.IMEM._1454_  (.A1(\u_cpu.IMEM._0144_ ),
    .A2(\u_cpu.IMEM._0294_ ),
    .B1(\u_cpu.IMEM._0470_ ),
    .B2(\u_cpu.IMEM._0471_ ),
    .C1(\u_cpu.IMEM._0109_ ),
    .X(\u_cpu.IMEM._0472_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.IMEM._1455_  (.A1(\u_cpu.IMEM._0468_ ),
    .A2(\u_cpu.IMEM._0469_ ),
    .B1_N(\u_cpu.IMEM._0472_ ),
    .Y(\u_cpu.IMEM._0473_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.IMEM._1456_  (.A1(\u_cpu.IMEM._0020_ ),
    .A2(\u_cpu.IMEM._0083_ ),
    .B1(\u_cpu.IMEM._0008_ ),
    .C1(\u_cpu.IMEM._0466_ ),
    .D1(\u_cpu.IMEM._0134_ ),
    .Y(\u_cpu.IMEM._0474_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1457_  (.A1(\u_cpu.IMEM._0185_ ),
    .A2(\u_cpu.IMEM._0041_ ),
    .A3(\u_cpu.IMEM._0010_ ),
    .B1(\u_cpu.IMEM._0474_ ),
    .C1(\u_cpu.IMEM._0379_ ),
    .X(\u_cpu.IMEM._0475_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1458_  (.A1(\u_cpu.IMEM._0059_ ),
    .A2(\u_cpu.IMEM._0165_ ),
    .B1(\u_cpu.IMEM._0403_ ),
    .C1(\u_cpu.IMEM._0191_ ),
    .Y(\u_cpu.IMEM._0476_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.IMEM._1459_  (.A(\u_cpu.IMEM._0037_ ),
    .B(\u_cpu.IMEM._0003_ ),
    .Y(\u_cpu.IMEM._0478_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.IMEM._1460_  (.A(\u_cpu.IMEM._0218_ ),
    .B(\u_cpu.IMEM._0037_ ),
    .Y(\u_cpu.IMEM._0479_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.IMEM._1461_  (.A1(\u_cpu.IMEM._0096_ ),
    .A2(\u_cpu.IMEM._0217_ ),
    .B1(\u_cpu.IMEM._0180_ ),
    .B2(\u_cpu.IMEM._0214_ ),
    .Y(\u_cpu.IMEM._0480_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.IMEM._1462_  (.A1(\u_cpu.IMEM._0281_ ),
    .A2(\u_cpu.IMEM._0476_ ),
    .A3(\u_cpu.IMEM._0478_ ),
    .B1(\u_cpu.IMEM._0479_ ),
    .B2(\u_cpu.IMEM._0480_ ),
    .X(\u_cpu.IMEM._0481_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.IMEM._1463_  (.A(\u_cpu.IMEM._0424_ ),
    .B(\u_cpu.IMEM._0175_ ),
    .Y(\u_cpu.IMEM._0482_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.IMEM._1464_  (.A(\u_cpu.IMEM._0008_ ),
    .B(\u_cpu.IMEM._0482_ ),
    .C(\u_cpu.IMEM._0086_ ),
    .X(\u_cpu.IMEM._0483_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1465_  (.A1(\u_cpu.IMEM._0615_ ),
    .A2(\u_cpu.IMEM._0179_ ),
    .B1(\u_cpu.IMEM._0483_ ),
    .C1(\u_cpu.IMEM._0699_ ),
    .X(\u_cpu.IMEM._0484_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1466_  (.A1(\u_cpu.IMEM._0028_ ),
    .A2(\u_cpu.IMEM._0441_ ),
    .B1(\u_cpu.IMEM._0333_ ),
    .C1(\u_cpu.IMEM._0484_ ),
    .Y(\u_cpu.IMEM._0485_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1467_  (.A1(\u_cpu.IMEM._0255_ ),
    .A2(\u_cpu.IMEM._0475_ ),
    .A3(\u_cpu.IMEM._0481_ ),
    .B1(\u_cpu.IMEM._0128_ ),
    .C1(\u_cpu.IMEM._0485_ ),
    .X(\u_cpu.IMEM._0486_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1468_  (.A1(\u_cpu.IMEM._0108_ ),
    .A2(\u_cpu.IMEM._0473_ ),
    .B1(\u_cpu.IMEM._0486_ ),
    .Y(\u_cpu.IMEM.rd[12] ));
 sky130_fd_sc_hd__and4bb_2 \u_cpu.IMEM._1469_  (.A_N(\u_cpu.IMEM._0530_ ),
    .B_N(\u_cpu.IMEM._0626_ ),
    .C(\u_cpu.IMEM._0019_ ),
    .D(\u_cpu.IMEM._0509_ ),
    .X(\u_cpu.IMEM._0488_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1470_  (.A1(\u_cpu.IMEM._0363_ ),
    .A2(\u_cpu.IMEM._0080_ ),
    .A3(\u_cpu.IMEM._0498_ ),
    .B1(\u_cpu.IMEM._0488_ ),
    .X(\u_cpu.IMEM._0489_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1471_  (.A1(\u_cpu.IMEM._0910_ ),
    .A2(\u_cpu.IMEM._0153_ ),
    .B1(\u_cpu.IMEM._0131_ ),
    .Y(\u_cpu.IMEM._0490_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1472_  (.A1(\u_cpu.IMEM._0489_ ),
    .A2(\u_cpu.IMEM._0131_ ),
    .B1(\u_cpu.IMEM._0490_ ),
    .Y(\u_cpu.IMEM._0491_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1473_  (.A1(\u_cpu.IMEM._0205_ ),
    .A2(\u_cpu.IMEM._0168_ ),
    .B1(\u_cpu.IMEM._0070_ ),
    .C1(\u_cpu.IMEM._0174_ ),
    .Y(\u_cpu.IMEM._0492_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1474_  (.A1(\u_cpu.IMEM._0229_ ),
    .A2(\u_cpu.IMEM._0132_ ),
    .A3(\u_cpu.IMEM._0048_ ),
    .B1(\u_cpu.IMEM._0667_ ),
    .X(\u_cpu.IMEM._0493_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1475_  (.A1(\u_cpu.IMEM._0492_ ),
    .A2(\u_cpu.IMEM._0454_ ),
    .A3(\u_cpu.IMEM._0493_ ),
    .B1(\u_cpu.IMEM._0333_ ),
    .X(\u_cpu.IMEM._0494_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1476_  (.A1(\u_cpu.IMEM._0491_ ),
    .A2(\u_cpu.IMEM._0710_ ),
    .B1(\u_cpu.IMEM._0494_ ),
    .Y(\u_cpu.IMEM._0495_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1477_  (.A1(\u_cpu.IMEM._0188_ ),
    .A2(\u_cpu.IMEM._0121_ ),
    .A3(\u_cpu.IMEM._0138_ ),
    .B1(\u_cpu.IMEM._0025_ ),
    .C1(\u_cpu.IMEM._0145_ ),
    .X(\u_cpu.IMEM._0496_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1478_  (.A(\u_cpu.IMEM._0037_ ),
    .B(\u_cpu.IMEM.a[8] ),
    .Y(\u_cpu.IMEM._0497_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1479_  (.A1(\u_cpu.IMEM._0139_ ),
    .A2(\u_cpu.IMEM._0124_ ),
    .A3(\u_cpu.IMEM._0143_ ),
    .B1(\u_cpu.IMEM._0497_ ),
    .X(\u_cpu.IMEM._0499_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.IMEM._1480_  (.A1(\u_cpu.IMEM._0351_ ),
    .A2(\u_cpu.IMEM._0141_ ),
    .B1(\u_cpu.IMEM._0496_ ),
    .B2(\u_cpu.IMEM._0499_ ),
    .C1(\u_cpu.IMEM._0316_ ),
    .Y(\u_cpu.IMEM._0500_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.IMEM._1481_  (.A(\u_cpu.IMEM._0096_ ),
    .B(\u_cpu.IMEM._0920_ ),
    .C(\u_cpu.IMEM._0415_ ),
    .D(\u_cpu.IMEM._0038_ ),
    .X(\u_cpu.IMEM._0501_ ));
 sky130_fd_sc_hd__or4b_2 \u_cpu.IMEM._1482_  (.A(\u_cpu.IMEM._0889_ ),
    .B(\u_cpu.IMEM._0075_ ),
    .C(\u_cpu.IMEM._0024_ ),
    .D_N(\u_cpu.IMEM._0184_ ),
    .X(\u_cpu.IMEM._0502_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.IMEM._1483_  (.A(\u_cpu.IMEM._0439_ ),
    .B(\u_cpu.IMEM._0176_ ),
    .C(\u_cpu.IMEM._0187_ ),
    .D(\u_cpu.IMEM._0000_ ),
    .Y(\u_cpu.IMEM._0503_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1484_  (.A1(\u_cpu.IMEM._0502_ ),
    .A2(\u_cpu.IMEM._0503_ ),
    .B1(\u_cpu.IMEM._0058_ ),
    .Y(\u_cpu.IMEM._0504_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.IMEM._1485_  (.A1(\u_cpu.IMEM._0501_ ),
    .A2(\u_cpu.IMEM._0504_ ),
    .B1(\u_cpu.IMEM._0125_ ),
    .X(\u_cpu.IMEM._0505_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.IMEM._1486_  (.A(\u_cpu.IMEM._0466_ ),
    .B(\u_cpu.IMEM._0044_ ),
    .C(\u_cpu.IMEM._0121_ ),
    .X(\u_cpu.IMEM._0506_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.IMEM._1487_  (.A1(\u_cpu.IMEM._0288_ ),
    .A2(\u_cpu.IMEM._0506_ ),
    .B1(\u_cpu.IMEM._0199_ ),
    .C1(\u_cpu.IMEM._0124_ ),
    .X(\u_cpu.IMEM._0507_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.IMEM._1488_  (.A1(\u_cpu.IMEM._0076_ ),
    .A2(\u_cpu.IMEM._0339_ ),
    .B1(\u_cpu.IMEM._0731_ ),
    .X(\u_cpu.IMEM._0508_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1489_  (.A1(\u_cpu.IMEM._0032_ ),
    .A2(\u_cpu.IMEM._0059_ ),
    .A3(\u_cpu.IMEM._0061_ ),
    .B1(\u_cpu.IMEM._0721_ ),
    .X(\u_cpu.IMEM._0510_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.IMEM._1490_  (.A1(\u_cpu.IMEM._0184_ ),
    .A2(\u_cpu.IMEM._0024_ ),
    .B1(\u_cpu.IMEM._0816_ ),
    .C1(\u_cpu.IMEM._0043_ ),
    .D1(\u_cpu.IMEM._0466_ ),
    .X(\u_cpu.IMEM._0511_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1491_  (.A(\u_cpu.IMEM._0046_ ),
    .X(\u_cpu.IMEM._0512_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.IMEM._1492_  (.A1(\u_cpu.IMEM._0082_ ),
    .A2(\u_cpu.IMEM._0138_ ),
    .B1(\u_cpu.IMEM._0152_ ),
    .B2(\u_cpu.IMEM._0636_ ),
    .C1(\u_cpu.IMEM._0120_ ),
    .X(\u_cpu.IMEM._0513_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.IMEM._1493_  (.A1(\u_cpu.IMEM._0510_ ),
    .A2(\u_cpu.IMEM._0511_ ),
    .B1(\u_cpu.IMEM._0512_ ),
    .B2(\u_cpu.IMEM._0513_ ),
    .X(\u_cpu.IMEM._0514_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.IMEM._1494_  (.A1(\u_cpu.IMEM._0182_ ),
    .A2(\u_cpu.IMEM._0497_ ),
    .A3(\u_cpu.IMEM._0508_ ),
    .B1(\u_cpu.IMEM._0514_ ),
    .B2(\u_cpu.IMEM._0351_ ),
    .X(\u_cpu.IMEM._0515_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.IMEM._1495_  (.A1(\u_cpu.IMEM._0306_ ),
    .A2(\u_cpu.IMEM._0505_ ),
    .A3(\u_cpu.IMEM._0507_ ),
    .B1(\u_cpu.IMEM._0515_ ),
    .Y(\u_cpu.IMEM._0516_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu.IMEM._1496_  (.A1_N(\u_cpu.IMEM._0495_ ),
    .A2_N(\u_cpu.IMEM._0500_ ),
    .B1(\u_cpu.IMEM._0128_ ),
    .B2(\u_cpu.IMEM._0516_ ),
    .Y(\u_cpu.IMEM.rd[13] ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.IMEM._1497_  (.A1(\u_cpu.IMEM._0753_ ),
    .A2(\u_cpu.IMEM._0059_ ),
    .A3(\u_cpu.IMEM._0415_ ),
    .B1(\u_cpu.IMEM._0000_ ),
    .B2(\u_cpu.IMEM._0150_ ),
    .X(\u_cpu.IMEM._0517_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.IMEM._1498_  (.A1(\u_cpu.IMEM._0046_ ),
    .A2(\u_cpu.IMEM._0482_ ),
    .A3(\u_cpu.IMEM._0190_ ),
    .B1(\u_cpu.IMEM._0396_ ),
    .B2(\u_cpu.IMEM._0142_ ),
    .X(\u_cpu.IMEM._0518_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.IMEM._1499_  (.A1_N(\u_cpu.IMEM._0268_ ),
    .A2_N(\u_cpu.IMEM._0517_ ),
    .B1(\u_cpu.IMEM._0518_ ),
    .B2(\u_cpu.IMEM._0699_ ),
    .X(\u_cpu.IMEM._0520_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1500_  (.A1(\u_cpu.IMEM._0133_ ),
    .A2(\u_cpu.IMEM._0118_ ),
    .B1(\u_cpu.IMEM._0604_ ),
    .C1(\u_cpu.IMEM._0187_ ),
    .X(\u_cpu.IMEM._0521_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1501_  (.A1(\u_cpu.IMEM._0015_ ),
    .A2(\u_cpu.IMEM._0191_ ),
    .A3(\u_cpu.IMEM._0287_ ),
    .B1(\u_cpu.IMEM._0037_ ),
    .X(\u_cpu.IMEM._0522_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1502_  (.A1(\u_cpu.IMEM._0889_ ),
    .A2(\u_cpu.IMEM._0795_ ),
    .A3(\u_cpu.IMEM._0021_ ),
    .B1(\u_cpu.IMEM._0594_ ),
    .X(\u_cpu.IMEM._0523_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.IMEM._1503_  (.A(\u_cpu.IMEM._0061_ ),
    .B(\u_cpu.IMEM._0086_ ),
    .C(\u_cpu.IMEM._0023_ ),
    .D(\u_cpu.IMEM._0238_ ),
    .Y(\u_cpu.IMEM._0524_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.IMEM._1504_  (.A1(\u_cpu.IMEM._0523_ ),
    .A2(\u_cpu.IMEM._0524_ ),
    .A3(\u_cpu.IMEM._0143_ ),
    .B1(\u_cpu.IMEM._0425_ ),
    .B2(\u_cpu.IMEM._0218_ ),
    .X(\u_cpu.IMEM._0525_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.IMEM._1505_  (.A1(\u_cpu.IMEM._0521_ ),
    .A2(\u_cpu.IMEM._0522_ ),
    .B1(\u_cpu.IMEM._0525_ ),
    .B2(\u_cpu.IMEM._0090_ ),
    .Y(\u_cpu.IMEM._0526_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.IMEM._1506_  (.A1(\u_cpu.IMEM._0425_ ),
    .A2(\u_cpu.IMEM._0094_ ),
    .B1(\u_cpu.IMEM._0090_ ),
    .C1(\u_cpu.IMEM._0465_ ),
    .Y(\u_cpu.IMEM._0527_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.IMEM._1507_  (.A(\u_cpu.IMEM._0424_ ),
    .B(\u_cpu.IMEM._0868_ ),
    .C(\u_cpu.IMEM._0338_ ),
    .X(\u_cpu.IMEM._0528_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1508_  (.A1(\u_cpu.IMEM._0604_ ),
    .A2(\u_cpu.IMEM._0488_ ),
    .A3(\u_cpu.IMEM._0528_ ),
    .B1(\u_cpu.IMEM._0657_ ),
    .X(\u_cpu.IMEM._0529_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1509_  (.A1(\u_cpu.IMEM._0187_ ),
    .A2(\u_cpu.IMEM._0042_ ),
    .A3(\u_cpu.IMEM._0041_ ),
    .B1(\u_cpu.IMEM._0038_ ),
    .X(\u_cpu.IMEM._0531_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.IMEM._1510_  (.A1(\u_cpu.IMEM._0699_ ),
    .A2(\u_cpu.IMEM._0464_ ),
    .B1(\u_cpu.IMEM._0529_ ),
    .B2(\u_cpu.IMEM._0531_ ),
    .X(\u_cpu.IMEM._0532_ ));
 sky130_fd_sc_hd__mux4_2 \u_cpu.IMEM._1511_  (.A0(\u_cpu.IMEM._0520_ ),
    .A1(\u_cpu.IMEM._0526_ ),
    .A2(\u_cpu.IMEM._0527_ ),
    .A3(\u_cpu.IMEM._0532_ ),
    .S0(\u_cpu.IMEM._0302_ ),
    .S1(\u_cpu.IMEM._0055_ ),
    .X(\u_cpu.IMEM._0533_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.IMEM._1512_  (.A(\u_cpu.IMEM._0533_ ),
    .X(\u_cpu.IMEM.rd[14] ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1513_  (.A1(\u_cpu.IMEM._0020_ ),
    .A2(\u_cpu.IMEM._0083_ ),
    .B1(\u_cpu.IMEM._0753_ ),
    .C1(\u_cpu.IMEM._0827_ ),
    .X(\u_cpu.IMEM._0534_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.IMEM._1514_  (.A1(\u_cpu.IMEM._0211_ ),
    .A2(\u_cpu.IMEM._0534_ ),
    .B1(\u_cpu.IMEM._0036_ ),
    .B2(\u_cpu.IMEM._0837_ ),
    .C1(\u_cpu.IMEM._0094_ ),
    .Y(\u_cpu.IMEM._0535_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1515_  (.A1(\u_cpu.IMEM._0059_ ),
    .A2(\u_cpu.IMEM._0152_ ),
    .B1(\u_cpu.IMEM._0063_ ),
    .C1(\u_cpu.IMEM._0753_ ),
    .Y(\u_cpu.IMEM._0536_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1516_  (.A1(\u_cpu.IMEM._0050_ ),
    .A2(\u_cpu.IMEM._0536_ ),
    .B1(\u_cpu.IMEM._0262_ ),
    .X(\u_cpu.IMEM._0537_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.IMEM._1517_  (.A(\u_cpu.IMEM._0774_ ),
    .B(\u_cpu.IMEM._0069_ ),
    .C(\u_cpu.IMEM._0018_ ),
    .D(\u_cpu.IMEM._0082_ ),
    .X(\u_cpu.IMEM._0538_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.IMEM._1518_  (.A1(\u_cpu.IMEM._0191_ ),
    .A2(\u_cpu.IMEM._0323_ ),
    .A3(\u_cpu.IMEM._0161_ ),
    .B1(\u_cpu.IMEM._0214_ ),
    .C1(\u_cpu.IMEM._0093_ ),
    .Y(\u_cpu.IMEM._0539_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1519_  (.A1(\u_cpu.IMEM._0512_ ),
    .A2(\u_cpu.IMEM._0448_ ),
    .A3(\u_cpu.IMEM._0538_ ),
    .B1(\u_cpu.IMEM._0539_ ),
    .C1(\u_cpu.IMEM._0110_ ),
    .X(\u_cpu.IMEM._0541_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1520_  (.A1(\u_cpu.IMEM._0355_ ),
    .A2(\u_cpu.IMEM._0535_ ),
    .A3(\u_cpu.IMEM._0537_ ),
    .B1(\u_cpu.IMEM._0541_ ),
    .X(\u_cpu.IMEM._0542_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1521_  (.A1(\u_cpu.IMEM._0165_ ),
    .A2(\u_cpu.IMEM._0189_ ),
    .B1(\u_cpu.IMEM._0434_ ),
    .Y(\u_cpu.IMEM._0543_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1522_  (.A1(\u_cpu.IMEM._0413_ ),
    .A2(\u_cpu.IMEM._0347_ ),
    .B1(\u_cpu.IMEM._0543_ ),
    .Y(\u_cpu.IMEM._0544_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.IMEM._1523_  (.A1(\u_cpu.IMEM._0189_ ),
    .A2(\u_cpu.IMEM._0315_ ),
    .B1(\u_cpu.IMEM._0225_ ),
    .B2(\u_cpu.IMEM._0544_ ),
    .C1(\u_cpu.IMEM._0699_ ),
    .X(\u_cpu.IMEM._0545_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1524_  (.A1(\u_cpu.IMEM._0134_ ),
    .A2(\u_cpu.IMEM._0162_ ),
    .B1(\u_cpu.IMEM._0236_ ),
    .Y(\u_cpu.IMEM._0546_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1525_  (.A(\u_cpu.IMEM._0806_ ),
    .B(\u_cpu.IMEM._0626_ ),
    .Y(\u_cpu.IMEM._0547_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1526_  (.A1(\u_cpu.IMEM._0231_ ),
    .A2(\u_cpu.IMEM._0547_ ),
    .B1(\u_cpu.IMEM._0002_ ),
    .Y(\u_cpu.IMEM._0548_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.IMEM._1527_  (.A1(\u_cpu.IMEM._0482_ ),
    .A2(\u_cpu.IMEM._0308_ ),
    .B1(\u_cpu.IMEM._0546_ ),
    .B2(\u_cpu.IMEM._0548_ ),
    .C1(\u_cpu.IMEM._0129_ ),
    .X(\u_cpu.IMEM._0549_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.IMEM._1528_  (.A1(\u_cpu.IMEM._0545_ ),
    .A2(\u_cpu.IMEM._0549_ ),
    .B1(\u_cpu.IMEM._0302_ ),
    .X(\u_cpu.IMEM._0550_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.IMEM._1529_  (.A1(\u_cpu.IMEM._0185_ ),
    .A2(\u_cpu.IMEM._0157_ ),
    .B1(\u_cpu.IMEM._0078_ ),
    .C1(\u_cpu.IMEM._0371_ ),
    .D1(\u_cpu.IMEM._0132_ ),
    .Y(\u_cpu.IMEM._0552_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1530_  (.A1(\u_cpu.IMEM._0153_ ),
    .A2(\u_cpu.IMEM._0552_ ),
    .B1(\u_cpu.IMEM._0447_ ),
    .X(\u_cpu.IMEM._0553_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.IMEM._1531_  (.A1(\u_cpu.IMEM._0010_ ),
    .A2(\u_cpu.IMEM._0287_ ),
    .B1(\u_cpu.IMEM._0071_ ),
    .B2(\u_cpu.IMEM._0407_ ),
    .X(\u_cpu.IMEM._0554_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1532_  (.A1(\u_cpu.IMEM._0553_ ),
    .A2(\u_cpu.IMEM._0554_ ),
    .B1(\u_cpu.IMEM._0173_ ),
    .Y(\u_cpu.IMEM._0555_ ));
 sky130_fd_sc_hd__a311o_2 \u_cpu.IMEM._1533_  (.A1(\u_cpu.IMEM._0439_ ),
    .A2(\u_cpu.IMEM._0434_ ),
    .A3(\u_cpu.IMEM._0018_ ),
    .B1(\u_cpu.IMEM._0088_ ),
    .C1(\u_cpu.IMEM._0142_ ),
    .X(\u_cpu.IMEM._0556_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.IMEM._1534_  (.A(\u_cpu.IMEM._0556_ ),
    .B(\u_cpu.IMEM._0447_ ),
    .C(\u_cpu.IMEM._0240_ ),
    .Y(\u_cpu.IMEM._0557_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.IMEM._1535_  (.A(\u_cpu.IMEM._0112_ ),
    .B(\u_cpu.IMEM._0022_ ),
    .C(\u_cpu.IMEM._0795_ ),
    .D(\u_cpu.IMEM._0927_ ),
    .X(\u_cpu.IMEM._0558_ ));
 sky130_fd_sc_hd__a311o_2 \u_cpu.IMEM._1536_  (.A1(\u_cpu.IMEM._0002_ ),
    .A2(\u_cpu.IMEM._0063_ ),
    .A3(\u_cpu.IMEM._0446_ ),
    .B1(\u_cpu.IMEM._0558_ ),
    .C1(\u_cpu.IMEM._0218_ ),
    .X(\u_cpu.IMEM._0559_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1537_  (.A1(\u_cpu.IMEM._0557_ ),
    .A2(\u_cpu.IMEM._0559_ ),
    .A3(\u_cpu.IMEM._0199_ ),
    .B1(\u_cpu.IMEM._0295_ ),
    .X(\u_cpu.IMEM._0560_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.IMEM._1538_  (.A(\u_cpu.IMEM._0230_ ),
    .B(\u_cpu.IMEM._0309_ ),
    .C(\u_cpu.IMEM._0037_ ),
    .X(\u_cpu.IMEM._0561_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1539_  (.A1(\u_cpu.IMEM._0257_ ),
    .A2(\u_cpu.IMEM._0138_ ),
    .A3(\u_cpu.IMEM._0217_ ),
    .B1(\u_cpu.IMEM._0025_ ),
    .C1(\u_cpu.IMEM._0225_ ),
    .X(\u_cpu.IMEM._0563_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1540_  (.A1(\u_cpu.IMEM._0239_ ),
    .A2(\u_cpu.IMEM._0212_ ),
    .A3(\u_cpu.IMEM._0241_ ),
    .B1(\u_cpu.IMEM._0129_ ),
    .X(\u_cpu.IMEM._0564_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.IMEM._1541_  (.A1(\u_cpu.IMEM._0078_ ),
    .A2(\u_cpu.IMEM._0561_ ),
    .B1(\u_cpu.IMEM._0563_ ),
    .B2(\u_cpu.IMEM._0564_ ),
    .C1(\u_cpu.IMEM._0255_ ),
    .Y(\u_cpu.IMEM._0565_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1542_  (.A1(\u_cpu.IMEM._0555_ ),
    .A2(\u_cpu.IMEM._0560_ ),
    .B1(\u_cpu.IMEM._0565_ ),
    .C1(\u_cpu.IMEM._0431_ ),
    .Y(\u_cpu.IMEM._0566_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.IMEM._1543_  (.A1(\u_cpu.IMEM._0431_ ),
    .A2(\u_cpu.IMEM._0542_ ),
    .A3(\u_cpu.IMEM._0550_ ),
    .B1(\u_cpu.IMEM._0566_ ),
    .Y(\u_cpu.IMEM.rd[15] ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.IMEM._1544_  (.A1(\u_cpu.IMEM._0927_ ),
    .A2(\u_cpu.IMEM._0795_ ),
    .B1(\u_cpu.IMEM._0184_ ),
    .C1(\u_cpu.IMEM._0112_ ),
    .X(\u_cpu.IMEM._0567_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1545_  (.A1(\u_cpu.IMEM._0413_ ),
    .A2(\u_cpu.IMEM._0347_ ),
    .B1(\u_cpu.IMEM._0567_ ),
    .Y(\u_cpu.IMEM._0568_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.IMEM._1546_  (.A1(\u_cpu.IMEM._0646_ ),
    .A2(\u_cpu.IMEM._0071_ ),
    .A3(\u_cpu.IMEM._0583_ ),
    .B1(\u_cpu.IMEM._0262_ ),
    .B2(\u_cpu.IMEM._0568_ ),
    .X(\u_cpu.IMEM._0569_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1547_  (.A1(\u_cpu.IMEM._0359_ ),
    .A2(\u_cpu.IMEM._0392_ ),
    .B1(\u_cpu.IMEM._0061_ ),
    .C1(\u_cpu.IMEM._0083_ ),
    .X(\u_cpu.IMEM._0570_ ));
 sky130_fd_sc_hd__o32ai_2 \u_cpu.IMEM._1548_  (.A1(\u_cpu.IMEM._0148_ ),
    .A2(\u_cpu.IMEM._0315_ ),
    .A3(\u_cpu.IMEM._0646_ ),
    .B1(\u_cpu.IMEM._0731_ ),
    .B2(\u_cpu.IMEM._0570_ ),
    .Y(\u_cpu.IMEM._0571_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1549_  (.A1(\u_cpu.IMEM._0571_ ),
    .A2(\u_cpu.IMEM._0090_ ),
    .B1(\u_cpu.IMEM._0295_ ),
    .Y(\u_cpu.IMEM._0573_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.IMEM._1550_  (.A1(\u_cpu.IMEM._0130_ ),
    .A2(\u_cpu.IMEM._0569_ ),
    .B1(\u_cpu.IMEM._0573_ ),
    .X(\u_cpu.IMEM._0574_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.IMEM._1551_  (.A(\u_cpu.IMEM._0165_ ),
    .B(\u_cpu.IMEM._0014_ ),
    .C(\u_cpu.IMEM._0009_ ),
    .D(\u_cpu.IMEM._0636_ ),
    .Y(\u_cpu.IMEM._0575_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1552_  (.A1(\u_cpu.IMEM._0088_ ),
    .A2(\u_cpu.IMEM._0298_ ),
    .A3(\u_cpu.IMEM._0235_ ),
    .B1(\u_cpu.IMEM._0575_ ),
    .C1(\u_cpu.IMEM._0615_ ),
    .X(\u_cpu.IMEM._0576_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1553_  (.A1(\u_cpu.IMEM._0502_ ),
    .A2(\u_cpu.IMEM._0512_ ),
    .A3(\u_cpu.IMEM._0153_ ),
    .B1(\u_cpu.IMEM._0103_ ),
    .X(\u_cpu.IMEM._0577_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1554_  (.A1(\u_cpu.IMEM._0403_ ),
    .A2(\u_cpu.IMEM._0068_ ),
    .B1(\u_cpu.IMEM._0191_ ),
    .X(\u_cpu.IMEM._0578_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1555_  (.A1(\u_cpu.IMEM._0230_ ),
    .A2(\u_cpu.IMEM._0415_ ),
    .A3(\u_cpu.IMEM._0646_ ),
    .B1(\u_cpu.IMEM._0615_ ),
    .C1(\u_cpu.IMEM._0578_ ),
    .X(\u_cpu.IMEM._0579_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.IMEM._1556_  (.A(\u_cpu.IMEM._0001_ ),
    .B(\u_cpu.IMEM._0827_ ),
    .C(\u_cpu.IMEM._0087_ ),
    .X(\u_cpu.IMEM._0580_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1557_  (.A1(\u_cpu.IMEM._0580_ ),
    .A2(\u_cpu.IMEM._0512_ ),
    .A3(\u_cpu.IMEM._0281_ ),
    .B1(\u_cpu.IMEM._0667_ ),
    .X(\u_cpu.IMEM._0581_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.IMEM._1558_  (.A1(\u_cpu.IMEM._0576_ ),
    .A2(\u_cpu.IMEM._0577_ ),
    .B1(\u_cpu.IMEM._0579_ ),
    .B2(\u_cpu.IMEM._0581_ ),
    .C1(\u_cpu.IMEM._0333_ ),
    .X(\u_cpu.IMEM._0582_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.IMEM._1559_  (.A1(\u_cpu.IMEM._0002_ ),
    .A2(\u_cpu.IMEM._0098_ ),
    .B1(\u_cpu.IMEM._0035_ ),
    .B2(\u_cpu.IMEM._0360_ ),
    .C1(\u_cpu.IMEM._0123_ ),
    .X(\u_cpu.IMEM._0584_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1560_  (.A1(\u_cpu.IMEM._0251_ ),
    .A2(\u_cpu.IMEM._0229_ ),
    .A3(\u_cpu.IMEM._0646_ ),
    .B1(\u_cpu.IMEM._0066_ ),
    .X(\u_cpu.IMEM._0585_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1561_  (.A1(\u_cpu.IMEM._0283_ ),
    .A2(\u_cpu.IMEM._0002_ ),
    .A3(\u_cpu.IMEM._0093_ ),
    .B1(\u_cpu.IMEM._0037_ ),
    .X(\u_cpu.IMEM._0586_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1562_  (.A1(\u_cpu.IMEM._0083_ ),
    .A2(\u_cpu.IMEM._0411_ ),
    .A3(\u_cpu.IMEM._0134_ ),
    .B1(\u_cpu.IMEM._0604_ ),
    .X(\u_cpu.IMEM._0587_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1563_  (.A1(\u_cpu.IMEM._0403_ ),
    .A2(\u_cpu.IMEM._0068_ ),
    .B1(\u_cpu.IMEM._0044_ ),
    .X(\u_cpu.IMEM._0588_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.IMEM._1564_  (.A1(\u_cpu.IMEM._0062_ ),
    .A2(\u_cpu.IMEM._0587_ ),
    .B1(\u_cpu.IMEM._0588_ ),
    .B2(\u_cpu.IMEM._0447_ ),
    .Y(\u_cpu.IMEM._0589_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.IMEM._1565_  (.A1(\u_cpu.IMEM._0584_ ),
    .A2(\u_cpu.IMEM._0585_ ),
    .B1(\u_cpu.IMEM._0586_ ),
    .B2(\u_cpu.IMEM._0589_ ),
    .X(\u_cpu.IMEM._0590_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.IMEM._1566_  (.A(\u_cpu.IMEM._0231_ ),
    .B(\u_cpu.IMEM._0657_ ),
    .C(\u_cpu.IMEM._0096_ ),
    .X(\u_cpu.IMEM._0591_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1567_  (.A1(\u_cpu.IMEM._0229_ ),
    .A2(\u_cpu.IMEM._0309_ ),
    .A3(\u_cpu.IMEM._0033_ ),
    .B1(\u_cpu.IMEM._0284_ ),
    .X(\u_cpu.IMEM._0592_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.IMEM._1568_  (.A1(\u_cpu.IMEM._0363_ ),
    .A2(\u_cpu.IMEM._0591_ ),
    .B1(\u_cpu.IMEM._0592_ ),
    .B2(\u_cpu.IMEM._0077_ ),
    .C1(\u_cpu.IMEM._0109_ ),
    .X(\u_cpu.IMEM._0593_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1569_  (.A1(\u_cpu.IMEM._0305_ ),
    .A2(\u_cpu.IMEM._0590_ ),
    .B1(\u_cpu.IMEM._0593_ ),
    .C1(\u_cpu.IMEM._0431_ ),
    .Y(\u_cpu.IMEM._0595_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.IMEM._1570_  (.A1(\u_cpu.IMEM._0431_ ),
    .A2(\u_cpu.IMEM._0574_ ),
    .A3(\u_cpu.IMEM._0582_ ),
    .B1(\u_cpu.IMEM._0595_ ),
    .Y(\u_cpu.IMEM.rd[16] ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1571_  (.A1(\u_cpu.IMEM._0040_ ),
    .A2(\u_cpu.IMEM._0415_ ),
    .B1(\u_cpu.IMEM._0098_ ),
    .Y(\u_cpu.IMEM._0596_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.IMEM._1572_  (.A1(\u_cpu.IMEM._0257_ ),
    .A2(\u_cpu.IMEM._0596_ ),
    .B1(\u_cpu.IMEM._0035_ ),
    .C1(\u_cpu.IMEM._0615_ ),
    .X(\u_cpu.IMEM._0597_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1573_  (.A1(\u_cpu.IMEM._0051_ ),
    .A2(\u_cpu.IMEM._0583_ ),
    .B1(\u_cpu.IMEM._0287_ ),
    .C1(\u_cpu.IMEM._0061_ ),
    .Y(\u_cpu.IMEM._0598_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1574_  (.A1(\u_cpu.IMEM._0598_ ),
    .A2(\u_cpu.IMEM._0512_ ),
    .A3(\u_cpu.IMEM._0167_ ),
    .B1(\u_cpu.IMEM._0103_ ),
    .X(\u_cpu.IMEM._0599_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.IMEM._1575_  (.A1(\u_cpu.IMEM._0403_ ),
    .A2(\u_cpu.IMEM._0065_ ),
    .A3(\u_cpu.IMEM._0080_ ),
    .B1(\u_cpu.IMEM._0567_ ),
    .Y(\u_cpu.IMEM._0600_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.IMEM._1576_  (.A1(\u_cpu.IMEM._0435_ ),
    .A2(\u_cpu.IMEM._0600_ ),
    .B1_N(\u_cpu.IMEM._0667_ ),
    .Y(\u_cpu.IMEM._0601_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1577_  (.A1(\u_cpu.IMEM._0068_ ),
    .A2(\u_cpu.IMEM._0069_ ),
    .B1(\u_cpu.IMEM._0044_ ),
    .X(\u_cpu.IMEM._0602_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1578_  (.A1(\u_cpu.IMEM._0049_ ),
    .A2(\u_cpu.IMEM._0051_ ),
    .B1(\u_cpu.IMEM._0095_ ),
    .X(\u_cpu.IMEM._0603_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1579_  (.A1(\u_cpu.IMEM._0920_ ),
    .A2(\u_cpu.IMEM._0078_ ),
    .A3(\u_cpu.IMEM._0371_ ),
    .B1(\u_cpu.IMEM._0603_ ),
    .X(\u_cpu.IMEM._0605_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1580_  (.A1(\u_cpu.IMEM._0602_ ),
    .A2(\u_cpu.IMEM._0605_ ),
    .B1(\u_cpu.IMEM._0145_ ),
    .Y(\u_cpu.IMEM._0606_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.IMEM._1581_  (.A1(\u_cpu.IMEM._0597_ ),
    .A2(\u_cpu.IMEM._0599_ ),
    .B1(\u_cpu.IMEM._0601_ ),
    .B2(\u_cpu.IMEM._0606_ ),
    .Y(\u_cpu.IMEM._0607_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1582_  (.A1(\u_cpu.IMEM._0404_ ),
    .A2(\u_cpu.IMEM._0448_ ),
    .B1(\u_cpu.IMEM._0447_ ),
    .Y(\u_cpu.IMEM._0608_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.IMEM._1583_  (.A1(\u_cpu.IMEM._0132_ ),
    .A2(\u_cpu.IMEM._0088_ ),
    .A3(\u_cpu.IMEM._0298_ ),
    .B1(\u_cpu.IMEM._0536_ ),
    .C1(\u_cpu.IMEM._0225_ ),
    .Y(\u_cpu.IMEM._0609_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1584_  (.A1(\u_cpu.IMEM._0077_ ),
    .A2(\u_cpu.IMEM._0608_ ),
    .A3(\u_cpu.IMEM._0609_ ),
    .B1(\u_cpu.IMEM._0109_ ),
    .X(\u_cpu.IMEM._0610_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1585_  (.A1(\u_cpu.IMEM._0096_ ),
    .A2(\u_cpu.IMEM._0162_ ),
    .A3(\u_cpu.IMEM._0197_ ),
    .B1(\u_cpu.IMEM._0476_ ),
    .C1(\u_cpu.IMEM._0731_ ),
    .X(\u_cpu.IMEM._0611_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.IMEM._1586_  (.A1(\u_cpu.IMEM._0483_ ),
    .A2(\u_cpu.IMEM._0611_ ),
    .B1(\u_cpu.IMEM._0208_ ),
    .X(\u_cpu.IMEM._0612_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.IMEM._1587_  (.A1_N(\u_cpu.IMEM._0469_ ),
    .A2_N(\u_cpu.IMEM._0607_ ),
    .B1(\u_cpu.IMEM._0610_ ),
    .B2(\u_cpu.IMEM._0612_ ),
    .Y(\u_cpu.IMEM._0613_ ));
 sky130_fd_sc_hd__and4bb_2 \u_cpu.IMEM._1588_  (.A_N(\u_cpu.IMEM._0927_ ),
    .B_N(\u_cpu.IMEM._0034_ ),
    .C(\u_cpu.IMEM._0626_ ),
    .D(\u_cpu.IMEM._0424_ ),
    .X(\u_cpu.IMEM._0614_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.IMEM._1589_  (.A(\u_cpu.IMEM._0093_ ),
    .B(\u_cpu.IMEM._0614_ ),
    .Y(\u_cpu.IMEM._0616_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1590_  (.A1(\u_cpu.IMEM._0583_ ),
    .A2(\u_cpu.IMEM._0858_ ),
    .B1(\u_cpu.IMEM._0307_ ),
    .C1(\u_cpu.IMEM._0403_ ),
    .Y(\u_cpu.IMEM._0617_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1591_  (.A1(\u_cpu.IMEM._0205_ ),
    .A2(\u_cpu.IMEM._0177_ ),
    .A3(\u_cpu.IMEM._0168_ ),
    .B1(\u_cpu.IMEM._0015_ ),
    .X(\u_cpu.IMEM._0618_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.IMEM._1592_  (.A1(\u_cpu.IMEM._0616_ ),
    .A2(\u_cpu.IMEM._0361_ ),
    .A3(\u_cpu.IMEM._0294_ ),
    .B1(\u_cpu.IMEM._0617_ ),
    .B2(\u_cpu.IMEM._0618_ ),
    .X(\u_cpu.IMEM._0619_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.IMEM._1593_  (.A1(\u_cpu.IMEM._0168_ ),
    .A2(\u_cpu.IMEM._0474_ ),
    .B1(\u_cpu.IMEM._0413_ ),
    .B2(\u_cpu.IMEM._0010_ ),
    .Y(\u_cpu.IMEM._0620_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1594_  (.A1(\u_cpu.IMEM._0205_ ),
    .A2(\u_cpu.IMEM._0168_ ),
    .B1(\u_cpu.IMEM._0134_ ),
    .C1(\u_cpu.IMEM._0190_ ),
    .Y(\u_cpu.IMEM._0621_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1595_  (.A1(\u_cpu.IMEM._0292_ ),
    .A2(\u_cpu.IMEM._0621_ ),
    .B1(\u_cpu.IMEM._0058_ ),
    .Y(\u_cpu.IMEM._0622_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1596_  (.A1(\u_cpu.IMEM._0620_ ),
    .A2(\u_cpu.IMEM._0622_ ),
    .B1(\u_cpu.IMEM._0028_ ),
    .Y(\u_cpu.IMEM._0623_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1597_  (.A1(\u_cpu.IMEM._0130_ ),
    .A2(\u_cpu.IMEM._0619_ ),
    .B1(\u_cpu.IMEM._0623_ ),
    .C1(\u_cpu.IMEM._0302_ ),
    .Y(\u_cpu.IMEM._0624_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1598_  (.A1(\u_cpu.IMEM._0064_ ),
    .A2(\u_cpu.IMEM._0176_ ),
    .B1(\u_cpu.IMEM._0178_ ),
    .Y(\u_cpu.IMEM._0625_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.IMEM._1599_  (.A1_N(\u_cpu.IMEM._0058_ ),
    .A2_N(\u_cpu.IMEM._0625_ ),
    .B1(\u_cpu.IMEM._0546_ ),
    .B2(\u_cpu.IMEM._0271_ ),
    .X(\u_cpu.IMEM._0627_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1600_  (.A1(\u_cpu.IMEM._0699_ ),
    .A2(\u_cpu.IMEM._0211_ ),
    .A3(\u_cpu.IMEM._0214_ ),
    .B1(\u_cpu.IMEM.a[8] ),
    .X(\u_cpu.IMEM._0628_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1601_  (.A1(\u_cpu.IMEM._0173_ ),
    .A2(\u_cpu.IMEM._0627_ ),
    .B1(\u_cpu.IMEM._0628_ ),
    .Y(\u_cpu.IMEM._0629_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1602_  (.A1(\u_cpu.IMEM._0624_ ),
    .A2(\u_cpu.IMEM._0629_ ),
    .B1(\u_cpu.IMEM._0128_ ),
    .Y(\u_cpu.IMEM._0630_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1603_  (.A1(\u_cpu.IMEM._0128_ ),
    .A2(\u_cpu.IMEM._0613_ ),
    .B1(\u_cpu.IMEM._0630_ ),
    .Y(\u_cpu.IMEM.rd[17] ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1604_  (.A1(\u_cpu.IMEM._0435_ ),
    .A2(\u_cpu.IMEM._0341_ ),
    .A3(\u_cpu.IMEM._0169_ ),
    .B1(\u_cpu.IMEM._0159_ ),
    .C1(\u_cpu.IMEM._0320_ ),
    .X(\u_cpu.IMEM._0631_ ));
 sky130_fd_sc_hd__or4_2 \u_cpu.IMEM._1605_  (.A(\u_cpu.IMEM._0927_ ),
    .B(\u_cpu.IMEM._0034_ ),
    .C(\u_cpu.IMEM._0795_ ),
    .D(\u_cpu.IMEM._0112_ ),
    .X(\u_cpu.IMEM._0632_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.IMEM._1606_  (.A1(\u_cpu.IMEM._0114_ ),
    .A2(\u_cpu.IMEM._0631_ ),
    .B1(\u_cpu.IMEM._0632_ ),
    .B2(\u_cpu.IMEM._0272_ ),
    .C1(\u_cpu.IMEM._0469_ ),
    .Y(\u_cpu.IMEM._0633_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.IMEM._1607_  (.A1(\u_cpu.IMEM._0570_ ),
    .A2(\u_cpu.IMEM._0374_ ),
    .B1(\u_cpu.IMEM._0588_ ),
    .B2(\u_cpu.IMEM._0312_ ),
    .C1(\u_cpu.IMEM._0028_ ),
    .X(\u_cpu.IMEM._0634_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1608_  (.A1(\u_cpu.IMEM._0710_ ),
    .A2(\u_cpu.IMEM._0621_ ),
    .B1(\u_cpu.IMEM._0305_ ),
    .C1(\u_cpu.IMEM._0634_ ),
    .Y(\u_cpu.IMEM._0635_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.IMEM._1609_  (.A(\u_cpu.IMEM._0163_ ),
    .B(\u_cpu.IMEM._0371_ ),
    .C(\u_cpu.IMEM._0309_ ),
    .X(\u_cpu.IMEM._0637_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.IMEM._1610_  (.A(\u_cpu.IMEM._0447_ ),
    .B(\u_cpu.IMEM._0600_ ),
    .Y(\u_cpu.IMEM._0638_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1611_  (.A1(\u_cpu.IMEM._0637_ ),
    .A2(\u_cpu.IMEM._0638_ ),
    .B1(\u_cpu.IMEM._0710_ ),
    .Y(\u_cpu.IMEM._0639_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1612_  (.A1(\u_cpu.IMEM._0044_ ),
    .A2(\u_cpu.IMEM._0042_ ),
    .A3(\u_cpu.IMEM._0030_ ),
    .B1(\u_cpu.IMEM._0038_ ),
    .X(\u_cpu.IMEM._0640_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.IMEM._1613_  (.A1(\u_cpu.IMEM._0450_ ),
    .A2(\u_cpu.IMEM._0079_ ),
    .B1(\u_cpu.IMEM._0148_ ),
    .B2(\u_cpu.IMEM._0150_ ),
    .C1(\u_cpu.IMEM._0512_ ),
    .Y(\u_cpu.IMEM._0641_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1614_  (.A1(\u_cpu.IMEM._0339_ ),
    .A2(\u_cpu.IMEM._0640_ ),
    .B1(\u_cpu.IMEM._0090_ ),
    .C1(\u_cpu.IMEM._0641_ ),
    .Y(\u_cpu.IMEM._0642_ ));
 sky130_fd_sc_hd__or4_2 \u_cpu.IMEM._1615_  (.A(\u_cpu.IMEM._0657_ ),
    .B(\u_cpu.IMEM._0157_ ),
    .C(\u_cpu.IMEM._0415_ ),
    .D(\u_cpu.IMEM._0315_ ),
    .X(\u_cpu.IMEM._0643_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1616_  (.A1(\u_cpu.IMEM._0642_ ),
    .A2(\u_cpu.IMEM._0643_ ),
    .A3(\u_cpu.IMEM._0333_ ),
    .B1(\u_cpu.IMEM.a[9] ),
    .X(\u_cpu.IMEM._0644_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1617_  (.A1(\u_cpu.IMEM._0573_ ),
    .A2(\u_cpu.IMEM._0639_ ),
    .B1(\u_cpu.IMEM._0644_ ),
    .Y(\u_cpu.IMEM._0645_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1618_  (.A1(\u_cpu.IMEM._0108_ ),
    .A2(\u_cpu.IMEM._0633_ ),
    .A3(\u_cpu.IMEM._0635_ ),
    .B1(\u_cpu.IMEM._0645_ ),
    .X(\u_cpu.IMEM.rd[18] ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1619_  (.A1(\u_cpu.IMEM._0230_ ),
    .A2(\u_cpu.IMEM._0157_ ),
    .A3(\u_cpu.IMEM._0033_ ),
    .B1(\u_cpu.IMEM._0339_ ),
    .X(\u_cpu.IMEM._0647_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.IMEM._1620_  (.A1(\u_cpu.IMEM._0137_ ),
    .A2(\u_cpu.IMEM._0142_ ),
    .A3(\u_cpu.IMEM._0396_ ),
    .B1(\u_cpu.IMEM._0647_ ),
    .B2(\u_cpu.IMEM._0479_ ),
    .X(\u_cpu.IMEM._0648_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1621_  (.A1(\u_cpu.IMEM._0131_ ),
    .A2(\u_cpu.IMEM._0228_ ),
    .A3(\u_cpu.IMEM._0041_ ),
    .B1(\u_cpu.IMEM._0638_ ),
    .X(\u_cpu.IMEM._0649_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.IMEM._1622_  (.A(\u_cpu.IMEM._0255_ ),
    .B(\u_cpu.IMEM._0173_ ),
    .Y(\u_cpu.IMEM._0650_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.IMEM._1623_  (.A1(\u_cpu.IMEM._0117_ ),
    .A2(\u_cpu.IMEM._0648_ ),
    .B1(\u_cpu.IMEM._0649_ ),
    .B2(\u_cpu.IMEM._0650_ ),
    .Y(\u_cpu.IMEM._0651_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.IMEM._1624_  (.A(\u_cpu.IMEM._0103_ ),
    .B(\u_cpu.IMEM._0216_ ),
    .C(\u_cpu.IMEM._0150_ ),
    .X(\u_cpu.IMEM._0652_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.IMEM._1625_  (.A(\u_cpu.IMEM._0411_ ),
    .B(\u_cpu.IMEM._0858_ ),
    .C(\u_cpu.IMEM._0187_ ),
    .D(\u_cpu.IMEM._0000_ ),
    .Y(\u_cpu.IMEM._0653_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1626_  (.A1(\u_cpu.IMEM._0433_ ),
    .A2(\u_cpu.IMEM._0653_ ),
    .B1(\u_cpu.IMEM._0225_ ),
    .Y(\u_cpu.IMEM._0654_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1627_  (.A1(\u_cpu.IMEM._0009_ ),
    .A2(\u_cpu.IMEM._0020_ ),
    .B1(\u_cpu.IMEM._0415_ ),
    .Y(\u_cpu.IMEM._0655_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.IMEM._1628_  (.A(\u_cpu.IMEM._0236_ ),
    .B(\u_cpu.IMEM._0407_ ),
    .C(\u_cpu.IMEM._0297_ ),
    .D(\u_cpu.IMEM._0655_ ),
    .X(\u_cpu.IMEM._0656_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1629_  (.A1(\u_cpu.IMEM._0654_ ),
    .A2(\u_cpu.IMEM._0656_ ),
    .B1(\u_cpu.IMEM._0125_ ),
    .Y(\u_cpu.IMEM._0658_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1630_  (.A1(\u_cpu.IMEM._0652_ ),
    .A2(\u_cpu.IMEM._0658_ ),
    .B1(\u_cpu.IMEM._0302_ ),
    .Y(\u_cpu.IMEM._0659_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1631_  (.A1(\u_cpu.IMEM._0033_ ),
    .A2(\u_cpu.IMEM._0251_ ),
    .B1(\u_cpu.IMEM._0347_ ),
    .Y(\u_cpu.IMEM._0660_ ));
 sky130_fd_sc_hd__a2bb2o_2 \u_cpu.IMEM._1632_  (.A1_N(\u_cpu.IMEM._0212_ ),
    .A2_N(\u_cpu.IMEM._0660_ ),
    .B1(\u_cpu.IMEM._0388_ ),
    .B2(\u_cpu.IMEM._0141_ ),
    .X(\u_cpu.IMEM._0661_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.IMEM._1633_  (.A1(\u_cpu.IMEM._0010_ ),
    .A2(\u_cpu.IMEM._0287_ ),
    .B1(\u_cpu.IMEM._0463_ ),
    .B2(\u_cpu.IMEM._0188_ ),
    .C1(\u_cpu.IMEM._0470_ ),
    .X(\u_cpu.IMEM._0662_ ));
 sky130_fd_sc_hd__a311oi_2 \u_cpu.IMEM._1634_  (.A1(\u_cpu.IMEM._0661_ ),
    .A2(\u_cpu.IMEM._0130_ ),
    .A3(\u_cpu.IMEM._0116_ ),
    .B1(\u_cpu.IMEM._0662_ ),
    .C1(\u_cpu.IMEM._0255_ ),
    .Y(\u_cpu.IMEM._0663_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1635_  (.A1(\u_cpu.IMEM._0659_ ),
    .A2(\u_cpu.IMEM._0663_ ),
    .B1(\u_cpu.IMEM._0246_ ),
    .Y(\u_cpu.IMEM._0664_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1636_  (.A1(\u_cpu.IMEM._0108_ ),
    .A2(\u_cpu.IMEM._0651_ ),
    .B1(\u_cpu.IMEM._0664_ ),
    .Y(\u_cpu.IMEM.rd[19] ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.IMEM._1637_  (.A1(\u_cpu.IMEM._0270_ ),
    .A2(\u_cpu.IMEM._0069_ ),
    .B1(\u_cpu.IMEM._0228_ ),
    .B2(\u_cpu.IMEM._0337_ ),
    .C1(\u_cpu.IMEM._0237_ ),
    .X(\u_cpu.IMEM._0665_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1638_  (.A1(\u_cpu.IMEM._0262_ ),
    .A2(\u_cpu.IMEM._0899_ ),
    .A3(\u_cpu.IMEM._0319_ ),
    .B1(\u_cpu.IMEM._0137_ ),
    .X(\u_cpu.IMEM._0666_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.IMEM._1639_  (.A1(\u_cpu.IMEM._0176_ ),
    .A2(\u_cpu.IMEM._0123_ ),
    .B1(\u_cpu.IMEM._0439_ ),
    .B2(\u_cpu.IMEM._0216_ ),
    .X(\u_cpu.IMEM._0668_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1640_  (.A1(\u_cpu.IMEM._0668_ ),
    .A2(\u_cpu.IMEM._0188_ ),
    .B1(\u_cpu.IMEM._0710_ ),
    .Y(\u_cpu.IMEM._0669_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.IMEM._1641_  (.A1(\u_cpu.IMEM._0665_ ),
    .A2(\u_cpu.IMEM._0666_ ),
    .B1(\u_cpu.IMEM._0669_ ),
    .B2(\u_cpu.IMEM._0412_ ),
    .C1(\u_cpu.IMEM._0117_ ),
    .Y(\u_cpu.IMEM._0670_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1642_  (.A1(\u_cpu.IMEM._0307_ ),
    .A2(\u_cpu.IMEM._0042_ ),
    .B1(\u_cpu.IMEM._0157_ ),
    .Y(\u_cpu.IMEM._0671_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.IMEM._1643_  (.A1(\u_cpu.IMEM._0216_ ),
    .A2(\u_cpu.IMEM._0671_ ),
    .B1(\u_cpu.IMEM._0536_ ),
    .B2(\u_cpu.IMEM._0050_ ),
    .C1(\u_cpu.IMEM._0058_ ),
    .X(\u_cpu.IMEM._0672_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1644_  (.A1(\u_cpu.IMEM._0069_ ),
    .A2(\u_cpu.IMEM._0287_ ),
    .A3(\u_cpu.IMEM._0540_ ),
    .B1(\u_cpu.IMEM._0319_ ),
    .X(\u_cpu.IMEM._0673_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1645_  (.A1(\u_cpu.IMEM._0673_ ),
    .A2(\u_cpu.IMEM._0094_ ),
    .B1(\u_cpu.IMEM._0351_ ),
    .Y(\u_cpu.IMEM._0674_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1646_  (.A1(\u_cpu.IMEM._0134_ ),
    .A2(\u_cpu.IMEM._0879_ ),
    .A3(\u_cpu.IMEM._0168_ ),
    .B1(\u_cpu.IMEM._0236_ ),
    .X(\u_cpu.IMEM._0675_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.IMEM._1647_  (.A1(\u_cpu.IMEM._0203_ ),
    .A2(\u_cpu.IMEM._0212_ ),
    .A3(\u_cpu.IMEM._0910_ ),
    .B1(\u_cpu.IMEM._0524_ ),
    .B2(\u_cpu.IMEM._0675_ ),
    .X(\u_cpu.IMEM._0676_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.IMEM._1648_  (.A1(\u_cpu.IMEM._0672_ ),
    .A2(\u_cpu.IMEM._0674_ ),
    .B1(\u_cpu.IMEM._0676_ ),
    .B2(\u_cpu.IMEM._0355_ ),
    .C1(\u_cpu.IMEM.a[9] ),
    .X(\u_cpu.IMEM._0677_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1649_  (.A1(\u_cpu.IMEM._0230_ ),
    .A2(\u_cpu.IMEM._0101_ ),
    .A3(\u_cpu.IMEM._0088_ ),
    .B1(\u_cpu.IMEM._0632_ ),
    .X(\u_cpu.IMEM._0679_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1650_  (.A1(\u_cpu.IMEM._0646_ ),
    .A2(\u_cpu.IMEM._0415_ ),
    .A3(\u_cpu.IMEM._0010_ ),
    .B1(\u_cpu.IMEM._0103_ ),
    .X(\u_cpu.IMEM._0680_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1651_  (.A1(\u_cpu.IMEM._0131_ ),
    .A2(\u_cpu.IMEM._0679_ ),
    .B1(\u_cpu.IMEM._0680_ ),
    .C1(\u_cpu.IMEM._0521_ ),
    .Y(\u_cpu.IMEM._0681_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1652_  (.A1(\u_cpu.IMEM._0540_ ),
    .A2(\u_cpu.IMEM._0235_ ),
    .B1(\u_cpu.IMEM._0208_ ),
    .Y(\u_cpu.IMEM._0682_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.IMEM._1653_  (.A(\u_cpu.IMEM._0868_ ),
    .B(\u_cpu.IMEM._0112_ ),
    .C(\u_cpu.IMEM._0795_ ),
    .X(\u_cpu.IMEM._0683_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.IMEM._1654_  (.A1(\u_cpu.IMEM._0683_ ),
    .A2(\u_cpu.IMEM._0528_ ),
    .B1(\u_cpu.IMEM._0262_ ),
    .X(\u_cpu.IMEM._0684_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1655_  (.A(\u_cpu.IMEM._0070_ ),
    .B(\u_cpu.IMEM._0238_ ),
    .Y(\u_cpu.IMEM._0685_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1656_  (.A1(\u_cpu.IMEM._0048_ ),
    .A2(\u_cpu.IMEM._0685_ ),
    .B1(\u_cpu.IMEM._0632_ ),
    .Y(\u_cpu.IMEM._0686_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1657_  (.A1(\u_cpu.IMEM._0489_ ),
    .A2(\u_cpu.IMEM._0435_ ),
    .B1(\u_cpu.IMEM._0686_ ),
    .Y(\u_cpu.IMEM._0687_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1658_  (.A1(\u_cpu.IMEM._0684_ ),
    .A2(\u_cpu.IMEM._0687_ ),
    .B1(\u_cpu.IMEM._0710_ ),
    .Y(\u_cpu.IMEM._0688_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1659_  (.A1(\u_cpu.IMEM._0660_ ),
    .A2(\u_cpu.IMEM._0617_ ),
    .B1(\u_cpu.IMEM._0237_ ),
    .Y(\u_cpu.IMEM._0690_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1660_  (.A1(\u_cpu.IMEM._0037_ ),
    .A2(\u_cpu.IMEM._0614_ ),
    .A3(\u_cpu.IMEM._0113_ ),
    .B1(\u_cpu.IMEM._0272_ ),
    .X(\u_cpu.IMEM._0691_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.IMEM._1661_  (.A1(\u_cpu.IMEM._0690_ ),
    .A2(\u_cpu.IMEM._0691_ ),
    .B1(\u_cpu.IMEM._0302_ ),
    .X(\u_cpu.IMEM._0692_ ));
 sky130_fd_sc_hd__a32oi_2 \u_cpu.IMEM._1662_  (.A1(\u_cpu.IMEM._0681_ ),
    .A2(\u_cpu.IMEM._0682_ ),
    .A3(\u_cpu.IMEM._0306_ ),
    .B1(\u_cpu.IMEM._0688_ ),
    .B2(\u_cpu.IMEM._0692_ ),
    .Y(\u_cpu.IMEM._0693_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.IMEM._1663_  (.A1(\u_cpu.IMEM._0670_ ),
    .A2(\u_cpu.IMEM._0677_ ),
    .B1(\u_cpu.IMEM._0128_ ),
    .B2(\u_cpu.IMEM._0693_ ),
    .Y(\u_cpu.IMEM.rd[20] ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1664_  (.A1(\u_cpu.IMEM._0041_ ),
    .A2(\u_cpu.IMEM._0603_ ),
    .B1(\u_cpu.IMEM._0062_ ),
    .Y(\u_cpu.IMEM._0694_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1665_  (.A1(\u_cpu.IMEM._0288_ ),
    .A2(\u_cpu.IMEM._0511_ ),
    .B1(\u_cpu.IMEM._0478_ ),
    .Y(\u_cpu.IMEM._0695_ ));
 sky130_fd_sc_hd__o41a_2 \u_cpu.IMEM._1666_  (.A1(\u_cpu.IMEM._0001_ ),
    .A2(\u_cpu.IMEM._0827_ ),
    .A3(\u_cpu.IMEM._0211_ ),
    .A4(\u_cpu.IMEM._0205_ ),
    .B1(\u_cpu.IMEM._0046_ ),
    .X(\u_cpu.IMEM._0696_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1667_  (.A1(\u_cpu.IMEM._0185_ ),
    .A2(\u_cpu.IMEM._0223_ ),
    .B1(\u_cpu.IMEM._0696_ ),
    .Y(\u_cpu.IMEM._0697_ ));
 sky130_fd_sc_hd__a311o_2 \u_cpu.IMEM._1668_  (.A1(\u_cpu.IMEM._0080_ ),
    .A2(\u_cpu.IMEM._0466_ ),
    .A3(\u_cpu.IMEM._0439_ ),
    .B1(\u_cpu.IMEM._0683_ ),
    .C1(\u_cpu.IMEM._0038_ ),
    .X(\u_cpu.IMEM._0698_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.IMEM._1669_  (.A(\u_cpu.IMEM._0077_ ),
    .B(\u_cpu.IMEM._0697_ ),
    .C(\u_cpu.IMEM._0698_ ),
    .Y(\u_cpu.IMEM._0700_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.IMEM._1670_  (.A1(\u_cpu.IMEM._0268_ ),
    .A2(\u_cpu.IMEM._0694_ ),
    .B1(\u_cpu.IMEM._0695_ ),
    .C1(\u_cpu.IMEM._0333_ ),
    .D1(\u_cpu.IMEM._0700_ ),
    .X(\u_cpu.IMEM._0701_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1671_  (.A1(\u_cpu.IMEM._0636_ ),
    .A2(\u_cpu.IMEM._0583_ ),
    .B1(\u_cpu.IMEM._0065_ ),
    .C1(\u_cpu.IMEM._0011_ ),
    .Y(\u_cpu.IMEM._0702_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1672_  (.A(\u_cpu.IMEM._0064_ ),
    .B(\u_cpu.IMEM._0197_ ),
    .Y(\u_cpu.IMEM._0703_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.IMEM._1673_  (.A1(\u_cpu.IMEM._0230_ ),
    .A2(\u_cpu.IMEM._0547_ ),
    .B1(\u_cpu.IMEM._0218_ ),
    .C1(\u_cpu.IMEM._0703_ ),
    .X(\u_cpu.IMEM._0704_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1674_  (.A1(\u_cpu.IMEM._0523_ ),
    .A2(\u_cpu.IMEM._0702_ ),
    .B1(\u_cpu.IMEM._0704_ ),
    .Y(\u_cpu.IMEM._0705_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1675_  (.A1(\u_cpu.IMEM._0174_ ),
    .A2(\u_cpu.IMEM._0083_ ),
    .B1(\u_cpu.IMEM._0020_ ),
    .Y(\u_cpu.IMEM._0706_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.IMEM._1676_  (.A1(\u_cpu.IMEM._0064_ ),
    .A2(\u_cpu.IMEM._0706_ ),
    .B1(\u_cpu.IMEM._0003_ ),
    .X(\u_cpu.IMEM._0707_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1677_  (.A1(\u_cpu.IMEM._0044_ ),
    .A2(\u_cpu.IMEM._0030_ ),
    .A3(\u_cpu.IMEM._0048_ ),
    .B1(\u_cpu.IMEM._0218_ ),
    .X(\u_cpu.IMEM._0708_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1678_  (.A1(\u_cpu.IMEM._0920_ ),
    .A2(\u_cpu.IMEM._0323_ ),
    .B1(\u_cpu.IMEM._0063_ ),
    .C1(\u_cpu.IMEM._0230_ ),
    .Y(\u_cpu.IMEM._0709_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu.IMEM._1679_  (.A1(\u_cpu.IMEM._0707_ ),
    .A2(\u_cpu.IMEM._0143_ ),
    .B1(\u_cpu.IMEM._0708_ ),
    .B2(\u_cpu.IMEM._0709_ ),
    .C1(\u_cpu.IMEM._0199_ ),
    .Y(\u_cpu.IMEM._0711_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.IMEM._1680_  (.A1(\u_cpu.IMEM._0114_ ),
    .A2(\u_cpu.IMEM._0705_ ),
    .B1(\u_cpu.IMEM._0711_ ),
    .C1(\u_cpu.IMEM._0306_ ),
    .Y(\u_cpu.IMEM._0712_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.IMEM._1681_  (.A1(\u_cpu.IMEM._0858_ ),
    .A2(\u_cpu.IMEM._0165_ ),
    .A3(\u_cpu.IMEM._0371_ ),
    .B1(\u_cpu.IMEM._0080_ ),
    .Y(\u_cpu.IMEM._0713_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1682_  (.A1(\u_cpu.IMEM._0447_ ),
    .A2(\u_cpu.IMEM._0713_ ),
    .A3(\u_cpu.IMEM._0235_ ),
    .B1(\u_cpu.IMEM._0521_ ),
    .X(\u_cpu.IMEM._0714_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.IMEM._1683_  (.A1(\u_cpu.IMEM._0173_ ),
    .A2(\u_cpu.IMEM._0714_ ),
    .B1(\u_cpu.IMEM._0140_ ),
    .X(\u_cpu.IMEM._0715_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.IMEM._1684_  (.A1(\u_cpu.IMEM._0309_ ),
    .A2(\u_cpu.IMEM._0371_ ),
    .A3(\u_cpu.IMEM._0010_ ),
    .B1(\u_cpu.IMEM._0071_ ),
    .B2(\u_cpu.IMEM._0364_ ),
    .X(\u_cpu.IMEM._0716_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1685_  (.A1(\u_cpu.IMEM._0281_ ),
    .A2(\u_cpu.IMEM._0524_ ),
    .B1(\u_cpu.IMEM._0058_ ),
    .X(\u_cpu.IMEM._0717_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1686_  (.A1(\u_cpu.IMEM._0716_ ),
    .A2(\u_cpu.IMEM._0717_ ),
    .B1(\u_cpu.IMEM._0130_ ),
    .Y(\u_cpu.IMEM._0718_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1687_  (.A1(\u_cpu.IMEM._0078_ ),
    .A2(\u_cpu.IMEM._0371_ ),
    .A3(\u_cpu.IMEM._0347_ ),
    .B1(\u_cpu.IMEM._0459_ ),
    .X(\u_cpu.IMEM._0719_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1688_  (.A1(\u_cpu.IMEM._0492_ ),
    .A2(\u_cpu.IMEM._0292_ ),
    .B1(\u_cpu.IMEM._0268_ ),
    .Y(\u_cpu.IMEM._0720_ ));
 sky130_fd_sc_hd__a311o_2 \u_cpu.IMEM._1689_  (.A1(\u_cpu.IMEM._0719_ ),
    .A2(\u_cpu.IMEM._0435_ ),
    .A3(\u_cpu.IMEM._0144_ ),
    .B1(\u_cpu.IMEM._0295_ ),
    .C1(\u_cpu.IMEM._0720_ ),
    .X(\u_cpu.IMEM._0722_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1690_  (.A1(\u_cpu.IMEM._0718_ ),
    .A2(\u_cpu.IMEM._0722_ ),
    .B1(\u_cpu.IMEM._0316_ ),
    .Y(\u_cpu.IMEM._0723_ ));
 sky130_fd_sc_hd__o32ai_2 \u_cpu.IMEM._1691_  (.A1(\u_cpu.IMEM._0431_ ),
    .A2(\u_cpu.IMEM._0701_ ),
    .A3(\u_cpu.IMEM._0712_ ),
    .B1(\u_cpu.IMEM._0715_ ),
    .B2(\u_cpu.IMEM._0723_ ),
    .Y(\u_cpu.IMEM.rd[21] ));
 sky130_fd_sc_hd__and3_2 \u_cpu.IMEM._1692_  (.A(\u_cpu.IMEM._0063_ ),
    .B(\u_cpu.IMEM._0176_ ),
    .C(\u_cpu.IMEM._0043_ ),
    .X(\u_cpu.IMEM._0724_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.IMEM._1693_  (.A1(\u_cpu.IMEM._0065_ ),
    .A2(\u_cpu.IMEM._0899_ ),
    .B1(\u_cpu.IMEM._0363_ ),
    .B2(\u_cpu.IMEM._0324_ ),
    .Y(\u_cpu.IMEM._0725_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.IMEM._1694_  (.A1(\u_cpu.IMEM._0724_ ),
    .A2(\u_cpu.IMEM._0100_ ),
    .B1(\u_cpu.IMEM._0124_ ),
    .B2(\u_cpu.IMEM._0725_ ),
    .C1(\u_cpu.IMEM._0125_ ),
    .X(\u_cpu.IMEM._0726_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1695_  (.A1(\u_cpu.IMEM._0363_ ),
    .A2(\u_cpu.IMEM._0257_ ),
    .A3(\u_cpu.IMEM._0119_ ),
    .B1(\u_cpu.IMEM._0123_ ),
    .X(\u_cpu.IMEM._0727_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.IMEM._1696_  (.A1(\u_cpu.IMEM._0145_ ),
    .A2(\u_cpu.IMEM._0136_ ),
    .B1(\u_cpu.IMEM._0448_ ),
    .B2(\u_cpu.IMEM._0727_ ),
    .C1(\u_cpu.IMEM._0208_ ),
    .X(\u_cpu.IMEM._0728_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1697_  (.A1(\u_cpu.IMEM._0060_ ),
    .A2(\u_cpu.IMEM._0238_ ),
    .B1(\u_cpu.IMEM._0540_ ),
    .C1(\u_cpu.IMEM._0287_ ),
    .Y(\u_cpu.IMEM._0729_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1698_  (.A1(\u_cpu.IMEM._0178_ ),
    .A2(\u_cpu.IMEM._0729_ ),
    .B1(\u_cpu.IMEM._0093_ ),
    .X(\u_cpu.IMEM._0730_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1699_  (.A1(\u_cpu.IMEM._0148_ ),
    .A2(\u_cpu.IMEM._0157_ ),
    .B1(\u_cpu.IMEM._0121_ ),
    .Y(\u_cpu.IMEM._0732_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1700_  (.A1(\u_cpu.IMEM._0920_ ),
    .A2(\u_cpu.IMEM._0323_ ),
    .B1(\u_cpu.IMEM._0132_ ),
    .Y(\u_cpu.IMEM._0733_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1701_  (.A1(\u_cpu.IMEM._0228_ ),
    .A2(\u_cpu.IMEM._0732_ ),
    .B1(\u_cpu.IMEM._0262_ ),
    .C1(\u_cpu.IMEM._0733_ ),
    .Y(\u_cpu.IMEM._0734_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1702_  (.A1(\u_cpu.IMEM._0730_ ),
    .A2(\u_cpu.IMEM._0734_ ),
    .B1(\u_cpu.IMEM._0208_ ),
    .Y(\u_cpu.IMEM._0735_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1703_  (.A1(\u_cpu.IMEM._0591_ ),
    .A2(\u_cpu.IMEM._0735_ ),
    .B1(\u_cpu.IMEM._0055_ ),
    .Y(\u_cpu.IMEM._0736_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.IMEM._1704_  (.A1(\u_cpu.IMEM._0316_ ),
    .A2(\u_cpu.IMEM._0726_ ),
    .A3(\u_cpu.IMEM._0728_ ),
    .B1(\u_cpu.IMEM._0736_ ),
    .Y(\u_cpu.IMEM._0737_ ));
 sky130_fd_sc_hd__a311o_2 \u_cpu.IMEM._1705_  (.A1(\u_cpu.IMEM._0078_ ),
    .A2(\u_cpu.IMEM._0371_ ),
    .A3(\u_cpu.IMEM._0030_ ),
    .B1(\u_cpu.IMEM._0298_ ),
    .C1(\u_cpu.IMEM._0064_ ),
    .X(\u_cpu.IMEM._0738_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1706_  (.A1(\u_cpu.IMEM._0121_ ),
    .A2(\u_cpu.IMEM._0018_ ),
    .B1(\u_cpu.IMEM._0096_ ),
    .X(\u_cpu.IMEM._0739_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1707_  (.A1(\u_cpu.IMEM._0228_ ),
    .A2(\u_cpu.IMEM._0287_ ),
    .B1(\u_cpu.IMEM._0141_ ),
    .Y(\u_cpu.IMEM._0740_ ));
 sky130_fd_sc_hd__a32oi_2 \u_cpu.IMEM._1708_  (.A1(\u_cpu.IMEM._0738_ ),
    .A2(\u_cpu.IMEM._0739_ ),
    .A3(\u_cpu.IMEM._0479_ ),
    .B1(\u_cpu.IMEM._0740_ ),
    .B2(\u_cpu.IMEM._0478_ ),
    .Y(\u_cpu.IMEM._0741_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1709_  (.A1(\u_cpu.IMEM._0434_ ),
    .A2(\u_cpu.IMEM._0411_ ),
    .A3(\u_cpu.IMEM._0041_ ),
    .B1(\u_cpu.IMEM._0236_ ),
    .X(\u_cpu.IMEM._0743_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1710_  (.A1(\u_cpu.IMEM._0060_ ),
    .A2(\u_cpu.IMEM._0049_ ),
    .B1(\u_cpu.IMEM._0001_ ),
    .C1(\u_cpu.IMEM._0018_ ),
    .Y(\u_cpu.IMEM._0744_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1711_  (.A1(\u_cpu.IMEM._0434_ ),
    .A2(\u_cpu.IMEM._0020_ ),
    .A3(\u_cpu.IMEM._0190_ ),
    .B1(\u_cpu.IMEM._0038_ ),
    .C1(\u_cpu.IMEM._0744_ ),
    .X(\u_cpu.IMEM._0745_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1712_  (.A1(\u_cpu.IMEM._0743_ ),
    .A2(\u_cpu.IMEM._0281_ ),
    .B1(\u_cpu.IMEM._0144_ ),
    .C1(\u_cpu.IMEM._0745_ ),
    .X(\u_cpu.IMEM._0746_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1713_  (.A1(\u_cpu.IMEM._0741_ ),
    .A2(\u_cpu.IMEM._0091_ ),
    .A3(\u_cpu.IMEM._0746_ ),
    .B1(\u_cpu.IMEM._0306_ ),
    .X(\u_cpu.IMEM._0747_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1714_  (.A1(\u_cpu.IMEM._0377_ ),
    .A2(\u_cpu.IMEM._0228_ ),
    .A3(\u_cpu.IMEM._0360_ ),
    .B1(\u_cpu.IMEM._0150_ ),
    .X(\u_cpu.IMEM._0748_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1715_  (.A1(\u_cpu.IMEM._0602_ ),
    .A2(\u_cpu.IMEM._0709_ ),
    .B1(\u_cpu.IMEM._0137_ ),
    .C1(\u_cpu.IMEM._0435_ ),
    .X(\u_cpu.IMEM._0749_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.IMEM._1716_  (.A1(\u_cpu.IMEM._0149_ ),
    .A2(\u_cpu.IMEM._0111_ ),
    .B1(\u_cpu.IMEM._0070_ ),
    .X(\u_cpu.IMEM._0750_ ));
 sky130_fd_sc_hd__a311oi_2 \u_cpu.IMEM._1717_  (.A1(\u_cpu.IMEM._0445_ ),
    .A2(\u_cpu.IMEM._0413_ ),
    .A3(\u_cpu.IMEM._0068_ ),
    .B1(\u_cpu.IMEM._0750_ ),
    .C1(\u_cpu.IMEM._0212_ ),
    .Y(\u_cpu.IMEM._0751_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.IMEM._1718_  (.A1(\u_cpu.IMEM._0013_ ),
    .A2(\u_cpu.IMEM._0190_ ),
    .B1(\u_cpu.IMEM._0434_ ),
    .C1(\u_cpu.IMEM._0162_ ),
    .Y(\u_cpu.IMEM._0752_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.IMEM._1719_  (.A1(\u_cpu.IMEM._0752_ ),
    .A2(\u_cpu.IMEM._0724_ ),
    .B1(\u_cpu.IMEM._0212_ ),
    .X(\u_cpu.IMEM._0754_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1720_  (.A1(\u_cpu.IMEM._0751_ ),
    .A2(\u_cpu.IMEM._0754_ ),
    .B1(\u_cpu.IMEM._0710_ ),
    .Y(\u_cpu.IMEM._0755_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.IMEM._1721_  (.A1(\u_cpu.IMEM._0272_ ),
    .A2(\u_cpu.IMEM._0748_ ),
    .B1(\u_cpu.IMEM._0749_ ),
    .C1(\u_cpu.IMEM._0055_ ),
    .D1(\u_cpu.IMEM._0755_ ),
    .X(\u_cpu.IMEM._0756_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu.IMEM._1722_  (.A1_N(\u_cpu.IMEM._0305_ ),
    .A2_N(\u_cpu.IMEM._0737_ ),
    .B1(\u_cpu.IMEM._0747_ ),
    .B2(\u_cpu.IMEM._0756_ ),
    .Y(\u_cpu.IMEM.rd[22] ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1723_  (.A1(\u_cpu.IMEM._0228_ ),
    .A2(\u_cpu.IMEM._0337_ ),
    .B1(\u_cpu.IMEM._0707_ ),
    .Y(\u_cpu.IMEM._0757_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1724_  (.A1(\u_cpu.IMEM._0331_ ),
    .A2(\u_cpu.IMEM._0317_ ),
    .B1(\u_cpu.IMEM._0295_ ),
    .Y(\u_cpu.IMEM._0758_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1725_  (.A1(\u_cpu.IMEM._0104_ ),
    .A2(\u_cpu.IMEM._0757_ ),
    .B1(\u_cpu.IMEM._0758_ ),
    .X(\u_cpu.IMEM._0759_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.IMEM._1726_  (.A1(\u_cpu.IMEM._0133_ ),
    .A2(\u_cpu.IMEM._0324_ ),
    .A3(\u_cpu.IMEM._0119_ ),
    .B1(\u_cpu.IMEM._0752_ ),
    .Y(\u_cpu.IMEM._0760_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.IMEM._1727_  (.A1(\u_cpu.IMEM._0003_ ),
    .A2(\u_cpu.IMEM._0096_ ),
    .A3(\u_cpu.IMEM._0364_ ),
    .B1(\u_cpu.IMEM._0474_ ),
    .B2(\u_cpu.IMEM._0168_ ),
    .X(\u_cpu.IMEM._0761_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.IMEM._1728_  (.A1(\u_cpu.IMEM._0124_ ),
    .A2(\u_cpu.IMEM._0760_ ),
    .B1(\u_cpu.IMEM._0761_ ),
    .X(\u_cpu.IMEM._0762_ ));
 sky130_fd_sc_hd__a2111o_2 \u_cpu.IMEM._1729_  (.A1(\u_cpu.IMEM._0816_ ),
    .A2(\u_cpu.IMEM._0051_ ),
    .B1(\u_cpu.IMEM._0070_ ),
    .C1(\u_cpu.IMEM._0721_ ),
    .D1(\u_cpu.IMEM._0377_ ),
    .X(\u_cpu.IMEM._0764_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.IMEM._1730_  (.A1(\u_cpu.IMEM._0364_ ),
    .A2(\u_cpu.IMEM._0315_ ),
    .B1(\u_cpu.IMEM._0216_ ),
    .B2(\u_cpu.IMEM._0150_ ),
    .C1(\u_cpu.IMEM._0764_ ),
    .Y(\u_cpu.IMEM._0765_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1731_  (.A1(\u_cpu.IMEM._0765_ ),
    .A2(\u_cpu.IMEM._0130_ ),
    .B1(\u_cpu.IMEM._0255_ ),
    .Y(\u_cpu.IMEM._0766_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1732_  (.A1(\u_cpu.IMEM._0114_ ),
    .A2(\u_cpu.IMEM._0762_ ),
    .B1(\u_cpu.IMEM._0766_ ),
    .Y(\u_cpu.IMEM._0767_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.IMEM._1733_  (.A(\u_cpu.IMEM._0013_ ),
    .B(\u_cpu.IMEM._0411_ ),
    .C(\u_cpu.IMEM._0134_ ),
    .X(\u_cpu.IMEM._0768_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.IMEM._1734_  (.A1(\u_cpu.IMEM._0281_ ),
    .A2(\u_cpu.IMEM._0502_ ),
    .A3(\u_cpu.IMEM._0768_ ),
    .B1(\u_cpu.IMEM._0131_ ),
    .Y(\u_cpu.IMEM._0769_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1735_  (.A1(\u_cpu.IMEM._0879_ ),
    .A2(\u_cpu.IMEM._0858_ ),
    .A3(\u_cpu.IMEM._0033_ ),
    .B1(\u_cpu.IMEM._0269_ ),
    .C1(\u_cpu.IMEM._0064_ ),
    .X(\u_cpu.IMEM._0770_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu.IMEM._1736_  (.A1(\u_cpu.IMEM._0435_ ),
    .A2(\u_cpu.IMEM._0770_ ),
    .B1(\u_cpu.IMEM._0768_ ),
    .C1(\u_cpu.IMEM._0502_ ),
    .D1(\u_cpu.IMEM._0281_ ),
    .X(\u_cpu.IMEM._0771_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.IMEM._1737_  (.A(\u_cpu.IMEM._0512_ ),
    .B(\u_cpu.IMEM._0142_ ),
    .C(\u_cpu.IMEM._0763_ ),
    .X(\u_cpu.IMEM._0772_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.IMEM._1738_  (.A1(\u_cpu.IMEM._0157_ ),
    .A2(\u_cpu.IMEM._0148_ ),
    .B1(\u_cpu.IMEM._0217_ ),
    .B2(\u_cpu.IMEM._0033_ ),
    .C1(\u_cpu.IMEM._0132_ ),
    .Y(\u_cpu.IMEM._0773_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1739_  (.A1(\u_cpu.IMEM._0773_ ),
    .A2(\u_cpu.IMEM._0702_ ),
    .B1(\u_cpu.IMEM._0094_ ),
    .Y(\u_cpu.IMEM._0775_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1740_  (.A1(\u_cpu.IMEM._0772_ ),
    .A2(\u_cpu.IMEM._0775_ ),
    .B1(\u_cpu.IMEM._0173_ ),
    .Y(\u_cpu.IMEM._0776_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.IMEM._1741_  (.A1(\u_cpu.IMEM._0114_ ),
    .A2(\u_cpu.IMEM._0769_ ),
    .A3(\u_cpu.IMEM._0771_ ),
    .B1(\u_cpu.IMEM._0776_ ),
    .C1(\u_cpu.IMEM._0469_ ),
    .Y(\u_cpu.IMEM._0777_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1742_  (.A1(\u_cpu.IMEM._0153_ ),
    .A2(\u_cpu.IMEM._0154_ ),
    .B1(\u_cpu.IMEM._0093_ ),
    .Y(\u_cpu.IMEM._0778_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1743_  (.A1(\u_cpu.IMEM._0281_ ),
    .A2(\u_cpu.IMEM._0492_ ),
    .B1(\u_cpu.IMEM._0229_ ),
    .Y(\u_cpu.IMEM._0779_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1744_  (.A1(\u_cpu.IMEM._0778_ ),
    .A2(\u_cpu.IMEM._0779_ ),
    .B1(\u_cpu.IMEM._0137_ ),
    .Y(\u_cpu.IMEM._0780_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1745_  (.A1(\u_cpu.IMEM._0307_ ),
    .A2(\u_cpu.IMEM._0323_ ),
    .A3(\u_cpu.IMEM._0858_ ),
    .B1(\u_cpu.IMEM._0003_ ),
    .C1(\u_cpu.IMEM._0598_ ),
    .X(\u_cpu.IMEM._0781_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.IMEM._1746_  (.A(\u_cpu.IMEM._0359_ ),
    .B(\u_cpu.IMEM._0014_ ),
    .C(\u_cpu.IMEM._0636_ ),
    .X(\u_cpu.IMEM._0782_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.IMEM._1747_  (.A1(\u_cpu.IMEM._0068_ ),
    .A2(\u_cpu.IMEM._0439_ ),
    .A3(\u_cpu.IMEM._0177_ ),
    .B1(\u_cpu.IMEM._0731_ ),
    .Y(\u_cpu.IMEM._0783_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1748_  (.A1(\u_cpu.IMEM._0782_ ),
    .A2(\u_cpu.IMEM._0252_ ),
    .B1(\u_cpu.IMEM._0783_ ),
    .Y(\u_cpu.IMEM._0784_ ));
 sky130_fd_sc_hd__nand3b_2 \u_cpu.IMEM._1749_  (.A_N(\u_cpu.IMEM._0781_ ),
    .B(\u_cpu.IMEM._0208_ ),
    .C(\u_cpu.IMEM._0784_ ),
    .Y(\u_cpu.IMEM._0786_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.IMEM._1750_  (.A1(\u_cpu.IMEM._0780_ ),
    .A2(\u_cpu.IMEM._0786_ ),
    .A3(\u_cpu.IMEM._0306_ ),
    .B1(\u_cpu.IMEM._0316_ ),
    .Y(\u_cpu.IMEM._0787_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.IMEM._1751_  (.A1(\u_cpu.IMEM._0246_ ),
    .A2(\u_cpu.IMEM._0759_ ),
    .A3(\u_cpu.IMEM._0767_ ),
    .B1(\u_cpu.IMEM._0777_ ),
    .B2(\u_cpu.IMEM._0787_ ),
    .X(\u_cpu.IMEM.rd[23] ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1752_  (.A1(\u_cpu.IMEM._0064_ ),
    .A2(\u_cpu.IMEM._0157_ ),
    .A3(\u_cpu.IMEM._0048_ ),
    .B1(\u_cpu.IMEM._0702_ ),
    .X(\u_cpu.IMEM._0788_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.IMEM._1753_  (.A1(\u_cpu.IMEM._0094_ ),
    .A2(\u_cpu.IMEM._0788_ ),
    .B1(\u_cpu.IMEM._0287_ ),
    .B2(\u_cpu.IMEM._0010_ ),
    .C1(\u_cpu.IMEM._0028_ ),
    .Y(\u_cpu.IMEM._0789_ ));
 sky130_fd_sc_hd__a32oi_2 \u_cpu.IMEM._1754_  (.A1(\u_cpu.IMEM._0445_ ),
    .A2(\u_cpu.IMEM._0018_ ),
    .A3(\u_cpu.IMEM._0439_ ),
    .B1(\u_cpu.IMEM._0713_ ),
    .B2(\u_cpu.IMEM._0446_ ),
    .Y(\u_cpu.IMEM._0790_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.IMEM._1755_  (.A1(\u_cpu.IMEM._0319_ ),
    .A2(\u_cpu.IMEM._0567_ ),
    .B1(\u_cpu.IMEM._0003_ ),
    .X(\u_cpu.IMEM._0791_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.IMEM._1756_  (.A(\u_cpu.IMEM._0144_ ),
    .B(\u_cpu.IMEM._0791_ ),
    .Y(\u_cpu.IMEM._0792_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1757_  (.A1(\u_cpu.IMEM._0145_ ),
    .A2(\u_cpu.IMEM._0790_ ),
    .B1(\u_cpu.IMEM._0792_ ),
    .Y(\u_cpu.IMEM._0793_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1758_  (.A1(\u_cpu.IMEM._0789_ ),
    .A2(\u_cpu.IMEM._0793_ ),
    .B1(\u_cpu.IMEM._0306_ ),
    .Y(\u_cpu.IMEM._0794_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1759_  (.A1(\u_cpu.IMEM._0190_ ),
    .A2(\u_cpu.IMEM._0411_ ),
    .A3(\u_cpu.IMEM._0040_ ),
    .B1(\u_cpu.IMEM._0191_ ),
    .X(\u_cpu.IMEM._0796_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1760_  (.A1(\u_cpu.IMEM._0150_ ),
    .A2(\u_cpu.IMEM._0575_ ),
    .B1(\u_cpu.IMEM._0512_ ),
    .Y(\u_cpu.IMEM._0797_ ));
 sky130_fd_sc_hd__a311o_2 \u_cpu.IMEM._1761_  (.A1(\u_cpu.IMEM._0447_ ),
    .A2(\u_cpu.IMEM._0376_ ),
    .A3(\u_cpu.IMEM._0796_ ),
    .B1(\u_cpu.IMEM._0137_ ),
    .C1(\u_cpu.IMEM._0797_ ),
    .X(\u_cpu.IMEM._0798_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1762_  (.A1(\u_cpu.IMEM._0377_ ),
    .A2(\u_cpu.IMEM._0744_ ),
    .B1(\u_cpu.IMEM._0598_ ),
    .Y(\u_cpu.IMEM._0799_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1763_  (.A1(\u_cpu.IMEM._0799_ ),
    .A2(\u_cpu.IMEM._0435_ ),
    .B1(\u_cpu.IMEM._0144_ ),
    .C1(\u_cpu.IMEM._0778_ ),
    .X(\u_cpu.IMEM._0800_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1764_  (.A1(\u_cpu.IMEM._0798_ ),
    .A2(\u_cpu.IMEM._0800_ ),
    .B1(\u_cpu.IMEM._0469_ ),
    .Y(\u_cpu.IMEM._0801_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.IMEM._1765_  (.A1(\u_cpu.IMEM._0323_ ),
    .A2(\u_cpu.IMEM._0309_ ),
    .B1(\u_cpu.IMEM._0212_ ),
    .C1(\u_cpu.IMEM._0119_ ),
    .D1(\u_cpu.IMEM._0324_ ),
    .Y(\u_cpu.IMEM._0802_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1766_  (.A1(\u_cpu.IMEM._0030_ ),
    .A2(\u_cpu.IMEM._0371_ ),
    .B1(\u_cpu.IMEM._0015_ ),
    .C1(\u_cpu.IMEM._0158_ ),
    .X(\u_cpu.IMEM._0803_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.IMEM._1767_  (.A1(\u_cpu.IMEM._0141_ ),
    .A2(\u_cpu.IMEM._0802_ ),
    .A3(\u_cpu.IMEM._0803_ ),
    .B1(\u_cpu.IMEM._0208_ ),
    .Y(\u_cpu.IMEM._0804_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.IMEM._1768_  (.A(\u_cpu.IMEM._0307_ ),
    .B(\u_cpu.IMEM._0287_ ),
    .C(\u_cpu.IMEM._0118_ ),
    .X(\u_cpu.IMEM._0805_ ));
 sky130_fd_sc_hd__a311o_2 \u_cpu.IMEM._1769_  (.A1(\u_cpu.IMEM._0002_ ),
    .A2(\u_cpu.IMEM._0407_ ),
    .A3(\u_cpu.IMEM._0446_ ),
    .B1(\u_cpu.IMEM._0750_ ),
    .C1(\u_cpu.IMEM._0218_ ),
    .X(\u_cpu.IMEM._0807_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1770_  (.A1(\u_cpu.IMEM._0145_ ),
    .A2(\u_cpu.IMEM._0770_ ),
    .A3(\u_cpu.IMEM._0805_ ),
    .B1(\u_cpu.IMEM._0199_ ),
    .C1(\u_cpu.IMEM._0807_ ),
    .X(\u_cpu.IMEM._0808_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1771_  (.A1(\u_cpu.IMEM._0009_ ),
    .A2(\u_cpu.IMEM._0088_ ),
    .A3(\u_cpu.IMEM._0298_ ),
    .B1(\u_cpu.IMEM._0046_ ),
    .X(\u_cpu.IMEM._0809_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1772_  (.A1(\u_cpu.IMEM._0013_ ),
    .A2(\u_cpu.IMEM._0165_ ),
    .A3(\u_cpu.IMEM._0014_ ),
    .B1(\u_cpu.IMEM._0252_ ),
    .X(\u_cpu.IMEM._0810_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu.IMEM._1773_  (.A1(\u_cpu.IMEM._0753_ ),
    .A2(\u_cpu.IMEM._0023_ ),
    .B1(\u_cpu.IMEM._0363_ ),
    .B2(\u_cpu.IMEM._0324_ ),
    .X(\u_cpu.IMEM._0811_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu.IMEM._1774_  (.A1_N(\u_cpu.IMEM._0809_ ),
    .A2_N(\u_cpu.IMEM._0810_ ),
    .B1(\u_cpu.IMEM._0512_ ),
    .B2(\u_cpu.IMEM._0811_ ),
    .X(\u_cpu.IMEM._0812_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.IMEM._1775_  (.A1(\u_cpu.IMEM._0331_ ),
    .A2(\u_cpu.IMEM._0317_ ),
    .B1(\u_cpu.IMEM._0130_ ),
    .B2(\u_cpu.IMEM._0812_ ),
    .C1(\u_cpu.IMEM._0255_ ),
    .Y(\u_cpu.IMEM._0813_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.IMEM._1776_  (.A1(\u_cpu.IMEM._0306_ ),
    .A2(\u_cpu.IMEM._0804_ ),
    .A3(\u_cpu.IMEM._0808_ ),
    .B1(\u_cpu.IMEM._0316_ ),
    .C1(\u_cpu.IMEM._0813_ ),
    .Y(\u_cpu.IMEM._0814_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.IMEM._1777_  (.A1(\u_cpu.IMEM._0431_ ),
    .A2(\u_cpu.IMEM._0794_ ),
    .A3(\u_cpu.IMEM._0801_ ),
    .B1(\u_cpu.IMEM._0814_ ),
    .Y(\u_cpu.IMEM.rd[24] ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1778_  (.A1(\u_cpu.IMEM._0575_ ),
    .A2(\u_cpu.IMEM._0598_ ),
    .B1(\u_cpu.IMEM._0123_ ),
    .Y(\u_cpu.IMEM._0815_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1779_  (.A1(\u_cpu.IMEM._0124_ ),
    .A2(\u_cpu.IMEM._0796_ ),
    .A3(\u_cpu.IMEM._0738_ ),
    .B1(\u_cpu.IMEM._0815_ ),
    .X(\u_cpu.IMEM._0817_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1780_  (.A(\u_cpu.IMEM._0780_ ),
    .B(\u_cpu.IMEM._0194_ ),
    .Y(\u_cpu.IMEM._0818_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1781_  (.A1(\u_cpu.IMEM._0114_ ),
    .A2(\u_cpu.IMEM._0817_ ),
    .B1(\u_cpu.IMEM._0818_ ),
    .Y(\u_cpu.IMEM._0819_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.IMEM._1782_  (.A(\u_cpu.IMEM._0827_ ),
    .B(\u_cpu.IMEM._0095_ ),
    .C(\u_cpu.IMEM._0049_ ),
    .X(\u_cpu.IMEM._0820_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.IMEM._1783_  (.A1(\u_cpu.IMEM._0820_ ),
    .A2(\u_cpu.IMEM._0724_ ),
    .B1(\u_cpu.IMEM._0123_ ),
    .X(\u_cpu.IMEM._0821_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.IMEM._1784_  (.A(\u_cpu.IMEM._0123_ ),
    .B(\u_cpu.IMEM._0161_ ),
    .C(\u_cpu.IMEM._0132_ ),
    .X(\u_cpu.IMEM._0822_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.IMEM._1785_  (.A1(\u_cpu.IMEM._0090_ ),
    .A2(\u_cpu.IMEM._0791_ ),
    .A3(\u_cpu.IMEM._0821_ ),
    .B1(\u_cpu.IMEM._0822_ ),
    .B2(\u_cpu.IMEM._0691_ ),
    .X(\u_cpu.IMEM._0823_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1786_  (.A1(\u_cpu.IMEM._0305_ ),
    .A2(\u_cpu.IMEM._0823_ ),
    .B1(\u_cpu.IMEM._0128_ ),
    .Y(\u_cpu.IMEM._0824_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1787_  (.A1(\u_cpu.IMEM._0440_ ),
    .A2(\u_cpu.IMEM._0621_ ),
    .A3(\u_cpu.IMEM._0764_ ),
    .B1(\u_cpu.IMEM._0699_ ),
    .X(\u_cpu.IMEM._0825_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1788_  (.A1(\u_cpu.IMEM._0141_ ),
    .A2(\u_cpu.IMEM._0143_ ),
    .B1(\u_cpu.IMEM._0129_ ),
    .X(\u_cpu.IMEM._0826_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1789_  (.A1(\u_cpu.IMEM._0141_ ),
    .A2(\u_cpu.IMEM._0503_ ),
    .B1(\u_cpu.IMEM._0129_ ),
    .C1(\u_cpu.IMEM._0058_ ),
    .X(\u_cpu.IMEM._0828_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.IMEM._1790_  (.A1(\u_cpu.IMEM._0825_ ),
    .A2(\u_cpu.IMEM._0826_ ),
    .A3(\u_cpu.IMEM._0828_ ),
    .B1(\u_cpu.IMEM._0194_ ),
    .Y(\u_cpu.IMEM._0829_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1791_  (.A1(\u_cpu.IMEM._0363_ ),
    .A2(\u_cpu.IMEM._0080_ ),
    .A3(\u_cpu.IMEM._0118_ ),
    .B1(\u_cpu.IMEM._0181_ ),
    .X(\u_cpu.IMEM._0830_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1792_  (.A1(\u_cpu.IMEM._0730_ ),
    .A2(\u_cpu.IMEM._0830_ ),
    .B1(\u_cpu.IMEM._0090_ ),
    .X(\u_cpu.IMEM._0831_ ));
 sky130_fd_sc_hd__or4_2 \u_cpu.IMEM._1793_  (.A(\u_cpu.IMEM._0309_ ),
    .B(\u_cpu.IMEM._0323_ ),
    .C(\u_cpu.IMEM._0583_ ),
    .D(\u_cpu.IMEM._0331_ ),
    .X(\u_cpu.IMEM._0832_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1794_  (.A1(\u_cpu.IMEM._0831_ ),
    .A2(\u_cpu.IMEM._0832_ ),
    .B1(\u_cpu.IMEM._0469_ ),
    .Y(\u_cpu.IMEM._0833_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1795_  (.A1(\u_cpu.IMEM._0829_ ),
    .A2(\u_cpu.IMEM._0833_ ),
    .B1(\u_cpu.IMEM._0246_ ),
    .Y(\u_cpu.IMEM._0834_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1796_  (.A1(\u_cpu.IMEM._0819_ ),
    .A2(\u_cpu.IMEM._0824_ ),
    .B1(\u_cpu.IMEM._0834_ ),
    .Y(\u_cpu.IMEM.rd[25] ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu.IMEM._1797_  (.A1(\u_cpu.IMEM._0411_ ),
    .A2(\u_cpu.IMEM._0000_ ),
    .B1(\u_cpu.IMEM._0002_ ),
    .C1(\u_cpu.IMEM._0003_ ),
    .D1(\u_cpu.IMEM._0052_ ),
    .Y(\u_cpu.IMEM._0835_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1798_  (.A1(\u_cpu.IMEM._0621_ ),
    .A2(\u_cpu.IMEM._0764_ ),
    .A3(\u_cpu.IMEM._0835_ ),
    .B1(\u_cpu.IMEM._0137_ ),
    .X(\u_cpu.IMEM._0836_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1799_  (.A1(\u_cpu.IMEM._0302_ ),
    .A2(\u_cpu.IMEM._0826_ ),
    .A3(\u_cpu.IMEM._0836_ ),
    .B1(\u_cpu.IMEM._0091_ ),
    .X(\u_cpu.IMEM._0838_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1800_  (.A1(\u_cpu.IMEM._0024_ ),
    .A2(\u_cpu.IMEM._0023_ ),
    .B1(\u_cpu.IMEM._0043_ ),
    .C1(\u_cpu.IMEM._0547_ ),
    .Y(\u_cpu.IMEM._0839_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1801_  (.A1(\u_cpu.IMEM._0729_ ),
    .A2(\u_cpu.IMEM._0839_ ),
    .B1(\u_cpu.IMEM._0058_ ),
    .X(\u_cpu.IMEM._0840_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1802_  (.A1(\u_cpu.IMEM._0830_ ),
    .A2(\u_cpu.IMEM._0840_ ),
    .B1(\u_cpu.IMEM._0130_ ),
    .Y(\u_cpu.IMEM._0841_ ));
 sky130_fd_sc_hd__a311oi_2 \u_cpu.IMEM._1803_  (.A1(\u_cpu.IMEM._0114_ ),
    .A2(\u_cpu.IMEM._0228_ ),
    .A3(\u_cpu.IMEM._0782_ ),
    .B1(\u_cpu.IMEM._0469_ ),
    .C1(\u_cpu.IMEM._0841_ ),
    .Y(\u_cpu.IMEM._0842_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1804_  (.A1(\u_cpu.IMEM._0307_ ),
    .A2(\u_cpu.IMEM._0231_ ),
    .A3(\u_cpu.IMEM._0042_ ),
    .B1(\u_cpu.IMEM._0614_ ),
    .X(\u_cpu.IMEM._0843_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1805_  (.A1(\u_cpu.IMEM._0435_ ),
    .A2(\u_cpu.IMEM._0843_ ),
    .B1(\u_cpu.IMEM._0815_ ),
    .Y(\u_cpu.IMEM._0844_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1806_  (.A1(\u_cpu.IMEM._0710_ ),
    .A2(\u_cpu.IMEM._0844_ ),
    .B1(\u_cpu.IMEM._0780_ ),
    .Y(\u_cpu.IMEM._0845_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.IMEM._1807_  (.A(\u_cpu.IMEM._0001_ ),
    .B(\u_cpu.IMEM._0032_ ),
    .C(\u_cpu.IMEM._0848_ ),
    .X(\u_cpu.IMEM._0846_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1808_  (.A1(\u_cpu.IMEM._0132_ ),
    .A2(\u_cpu.IMEM._0148_ ),
    .A3(\u_cpu.IMEM._0309_ ),
    .B1(\u_cpu.IMEM._0066_ ),
    .X(\u_cpu.IMEM._0847_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1809_  (.A1(\u_cpu.IMEM._0187_ ),
    .A2(\u_cpu.IMEM._0042_ ),
    .A3(\u_cpu.IMEM._0018_ ),
    .B1(\u_cpu.IMEM._0280_ ),
    .X(\u_cpu.IMEM._0849_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.IMEM._1810_  (.A(\u_cpu.IMEM._0237_ ),
    .B(\u_cpu.IMEM._0849_ ),
    .Y(\u_cpu.IMEM._0850_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.IMEM._1811_  (.A1(\u_cpu.IMEM._0846_ ),
    .A2(\u_cpu.IMEM._0847_ ),
    .B1(\u_cpu.IMEM._0850_ ),
    .B2(\u_cpu.IMEM._0691_ ),
    .C1(\u_cpu.IMEM._0302_ ),
    .X(\u_cpu.IMEM._0851_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1812_  (.A1(\u_cpu.IMEM._0845_ ),
    .A2(\u_cpu.IMEM._0117_ ),
    .B1(\u_cpu.IMEM._0851_ ),
    .Y(\u_cpu.IMEM._0852_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.IMEM._1813_  (.A1(\u_cpu.IMEM._0838_ ),
    .A2(\u_cpu.IMEM._0842_ ),
    .B1(\u_cpu.IMEM._0246_ ),
    .B2(\u_cpu.IMEM._0852_ ),
    .Y(\u_cpu.IMEM.rd[26] ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.IMEM._1814_  (.A1(\u_cpu.IMEM._0307_ ),
    .A2(\u_cpu.IMEM._0180_ ),
    .B1(\u_cpu.IMEM._0298_ ),
    .B2(\u_cpu.IMEM._0099_ ),
    .C1(\u_cpu.IMEM._0093_ ),
    .X(\u_cpu.IMEM._0853_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1815_  (.A1(\u_cpu.IMEM._0853_ ),
    .A2(\u_cpu.IMEM._0815_ ),
    .B1(\u_cpu.IMEM._0199_ ),
    .Y(\u_cpu.IMEM._0854_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1816_  (.A(\u_cpu.IMEM._0780_ ),
    .B(\u_cpu.IMEM._0854_ ),
    .Y(\u_cpu.IMEM._0855_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1817_  (.A1(\u_cpu.IMEM._0596_ ),
    .A2(\u_cpu.IMEM._0763_ ),
    .B1(\u_cpu.IMEM._0724_ ),
    .Y(\u_cpu.IMEM._0856_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1818_  (.A1(\u_cpu.IMEM._0145_ ),
    .A2(\u_cpu.IMEM._0856_ ),
    .B1(\u_cpu.IMEM._0614_ ),
    .C1(\u_cpu.IMEM._0199_ ),
    .Y(\u_cpu.IMEM._0857_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.IMEM._1819_  (.A(\u_cpu.IMEM._0307_ ),
    .B(\u_cpu.IMEM._0231_ ),
    .C(\u_cpu.IMEM._0547_ ),
    .X(\u_cpu.IMEM._0859_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1820_  (.A1(\u_cpu.IMEM._0724_ ),
    .A2(\u_cpu.IMEM._0859_ ),
    .B1(\u_cpu.IMEM._0077_ ),
    .C1(\u_cpu.IMEM._0124_ ),
    .Y(\u_cpu.IMEM._0860_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1821_  (.A1(\u_cpu.IMEM._0857_ ),
    .A2(\u_cpu.IMEM._0860_ ),
    .B1(\u_cpu.IMEM._0194_ ),
    .Y(\u_cpu.IMEM._0861_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1822_  (.A1(\u_cpu.IMEM._0855_ ),
    .A2(\u_cpu.IMEM._0117_ ),
    .B1(\u_cpu.IMEM._0861_ ),
    .Y(\u_cpu.IMEM._0862_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1823_  (.A1(\u_cpu.IMEM._0825_ ),
    .A2(\u_cpu.IMEM._0826_ ),
    .B1(\u_cpu.IMEM._0255_ ),
    .Y(\u_cpu.IMEM._0863_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1824_  (.A1(\u_cpu.IMEM._0178_ ),
    .A2(\u_cpu.IMEM._0536_ ),
    .B1(\u_cpu.IMEM._0212_ ),
    .Y(\u_cpu.IMEM._0864_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1825_  (.A1(\u_cpu.IMEM._0182_ ),
    .A2(\u_cpu.IMEM._0864_ ),
    .B1(\u_cpu.IMEM._0077_ ),
    .Y(\u_cpu.IMEM._0865_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1826_  (.A1(\u_cpu.IMEM._0832_ ),
    .A2(\u_cpu.IMEM._0865_ ),
    .B1(\u_cpu.IMEM._0469_ ),
    .Y(\u_cpu.IMEM._0866_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1827_  (.A1(\u_cpu.IMEM._0863_ ),
    .A2(\u_cpu.IMEM._0866_ ),
    .B1(\u_cpu.IMEM._0246_ ),
    .Y(\u_cpu.IMEM._0867_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1828_  (.A1(\u_cpu.IMEM._0108_ ),
    .A2(\u_cpu.IMEM._0862_ ),
    .B1(\u_cpu.IMEM._0867_ ),
    .Y(\u_cpu.IMEM.rd[27] ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1829_  (.A1(\u_cpu.IMEM._0694_ ),
    .A2(\u_cpu.IMEM._0094_ ),
    .B1(\u_cpu.IMEM._0090_ ),
    .C1(\u_cpu.IMEM._0504_ ),
    .X(\u_cpu.IMEM._0869_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.IMEM._1830_  (.A1(\u_cpu.IMEM._0002_ ),
    .A2(\u_cpu.IMEM._0217_ ),
    .B1(\u_cpu.IMEM._0251_ ),
    .B2(\u_cpu.IMEM._0252_ ),
    .Y(\u_cpu.IMEM._0870_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1831_  (.A1(\u_cpu.IMEM._0870_ ),
    .A2(\u_cpu.IMEM._0435_ ),
    .B1(\u_cpu.IMEM._0137_ ),
    .Y(\u_cpu.IMEM._0871_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1832_  (.A1(\u_cpu.IMEM._0763_ ),
    .A2(\u_cpu.IMEM._0498_ ),
    .A3(\u_cpu.IMEM._0363_ ),
    .B1(\u_cpu.IMEM._0546_ ),
    .X(\u_cpu.IMEM._0872_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1833_  (.A1(\u_cpu.IMEM._0871_ ),
    .A2(\u_cpu.IMEM._0872_ ),
    .B1(\u_cpu.IMEM._0333_ ),
    .Y(\u_cpu.IMEM._0873_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu.IMEM._1834_  (.A1(\u_cpu.IMEM._0869_ ),
    .A2(\u_cpu.IMEM._0873_ ),
    .B1(\u_cpu.IMEM._0845_ ),
    .B2(\u_cpu.IMEM._0117_ ),
    .Y(\u_cpu.IMEM._0874_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1835_  (.A1(\u_cpu.IMEM._0536_ ),
    .A2(\u_cpu.IMEM._0839_ ),
    .B1(\u_cpu.IMEM._0447_ ),
    .Y(\u_cpu.IMEM._0875_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1836_  (.A1(\u_cpu.IMEM._0182_ ),
    .A2(\u_cpu.IMEM._0875_ ),
    .B1(\u_cpu.IMEM._0125_ ),
    .Y(\u_cpu.IMEM._0876_ ));
 sky130_fd_sc_hd__or4_2 \u_cpu.IMEM._1837_  (.A(\u_cpu.IMEM._0216_ ),
    .B(\u_cpu.IMEM._0185_ ),
    .C(\u_cpu.IMEM._0309_ ),
    .D(\u_cpu.IMEM._0331_ ),
    .X(\u_cpu.IMEM._0877_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1838_  (.A1(\u_cpu.IMEM._0876_ ),
    .A2(\u_cpu.IMEM._0877_ ),
    .B1(\u_cpu.IMEM._0469_ ),
    .Y(\u_cpu.IMEM._0878_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1839_  (.A1(\u_cpu.IMEM._0863_ ),
    .A2(\u_cpu.IMEM._0878_ ),
    .B1(\u_cpu.IMEM._0246_ ),
    .Y(\u_cpu.IMEM._0880_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1840_  (.A1(\u_cpu.IMEM._0108_ ),
    .A2(\u_cpu.IMEM._0874_ ),
    .B1(\u_cpu.IMEM._0880_ ),
    .Y(\u_cpu.IMEM.rd[28] ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1841_  (.A1(\u_cpu.IMEM._0753_ ),
    .A2(\u_cpu.IMEM._0879_ ),
    .A3(\u_cpu.IMEM._0377_ ),
    .B1(\u_cpu.IMEM._0685_ ),
    .X(\u_cpu.IMEM._0881_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.IMEM._1842_  (.A1(\u_cpu.IMEM._0225_ ),
    .A2(\u_cpu.IMEM._0881_ ),
    .B1(\u_cpu.IMEM._0546_ ),
    .B2(\u_cpu.IMEM._0081_ ),
    .Y(\u_cpu.IMEM._0882_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.IMEM._1843_  (.A(\u_cpu.IMEM._0882_ ),
    .B(\u_cpu.IMEM._0028_ ),
    .Y(\u_cpu.IMEM._0883_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1844_  (.A1(\u_cpu.IMEM._0148_ ),
    .A2(\u_cpu.IMEM._0411_ ),
    .B1(\u_cpu.IMEM._0353_ ),
    .Y(\u_cpu.IMEM._0884_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu.IMEM._1845_  (.A1(\u_cpu.IMEM._0615_ ),
    .A2(\u_cpu.IMEM._0121_ ),
    .B1(\u_cpu.IMEM._0534_ ),
    .B2(\u_cpu.IMEM._0884_ ),
    .C1(\u_cpu.IMEM._0129_ ),
    .X(\u_cpu.IMEM._0885_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1846_  (.A1(\u_cpu.IMEM._0883_ ),
    .A2(\u_cpu.IMEM._0885_ ),
    .B1(\u_cpu.IMEM._0194_ ),
    .Y(\u_cpu.IMEM._0886_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1847_  (.A1(\u_cpu.IMEM._0855_ ),
    .A2(\u_cpu.IMEM._0117_ ),
    .B1(\u_cpu.IMEM._0886_ ),
    .Y(\u_cpu.IMEM._0887_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1848_  (.A1(\u_cpu.IMEM._0865_ ),
    .A2(\u_cpu.IMEM._0877_ ),
    .B1(\u_cpu.IMEM._0469_ ),
    .Y(\u_cpu.IMEM._0888_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1849_  (.A1(\u_cpu.IMEM._0863_ ),
    .A2(\u_cpu.IMEM._0888_ ),
    .B1(\u_cpu.IMEM._0431_ ),
    .Y(\u_cpu.IMEM._0890_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1850_  (.A1(\u_cpu.IMEM._0108_ ),
    .A2(\u_cpu.IMEM._0887_ ),
    .B1(\u_cpu.IMEM._0890_ ),
    .Y(\u_cpu.IMEM.rd[29] ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.IMEM._1851_  (.A1(\u_cpu.IMEM._0079_ ),
    .A2(\u_cpu.IMEM._0450_ ),
    .B1(\u_cpu.IMEM._0161_ ),
    .B2(\u_cpu.IMEM._0169_ ),
    .C1(\u_cpu.IMEM._0058_ ),
    .X(\u_cpu.IMEM._0891_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1852_  (.A1(\u_cpu.IMEM._0763_ ),
    .A2(\u_cpu.IMEM._0583_ ),
    .A3(\u_cpu.IMEM._0377_ ),
    .B1(\u_cpu.IMEM._0580_ ),
    .C1(\u_cpu.IMEM._0237_ ),
    .X(\u_cpu.IMEM._0892_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1853_  (.A1(\u_cpu.IMEM._0228_ ),
    .A2(\u_cpu.IMEM._0837_ ),
    .B1(\u_cpu.IMEM._0237_ ),
    .Y(\u_cpu.IMEM._0893_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu.IMEM._1854_  (.A1(\u_cpu.IMEM._0089_ ),
    .A2(\u_cpu.IMEM._0810_ ),
    .A3(\u_cpu.IMEM._0058_ ),
    .B1(\u_cpu.IMEM._0497_ ),
    .Y(\u_cpu.IMEM._0894_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1855_  (.A1(\u_cpu.IMEM._0266_ ),
    .A2(\u_cpu.IMEM._0893_ ),
    .B1(\u_cpu.IMEM._0894_ ),
    .Y(\u_cpu.IMEM._0895_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1856_  (.A1(\u_cpu.IMEM._0174_ ),
    .A2(\u_cpu.IMEM._0020_ ),
    .B1(\u_cpu.IMEM._0013_ ),
    .C1(\u_cpu.IMEM._0011_ ),
    .X(\u_cpu.IMEM._0896_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.IMEM._1857_  (.A1(\u_cpu.IMEM._0143_ ),
    .A2(\u_cpu.IMEM._0896_ ),
    .B1(\u_cpu.IMEM._0225_ ),
    .Y(\u_cpu.IMEM._0897_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1858_  (.A1(\u_cpu.IMEM._0161_ ),
    .A2(\u_cpu.IMEM._0229_ ),
    .A3(\u_cpu.IMEM._0230_ ),
    .B1(\u_cpu.IMEM._0066_ ),
    .X(\u_cpu.IMEM._0898_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.IMEM._1859_  (.A(\u_cpu.IMEM._0482_ ),
    .B(\u_cpu.IMEM._0721_ ),
    .C(\u_cpu.IMEM._0060_ ),
    .X(\u_cpu.IMEM._0900_ ));
 sky130_fd_sc_hd__a311o_2 \u_cpu.IMEM._1860_  (.A1(\u_cpu.IMEM._0218_ ),
    .A2(\u_cpu.IMEM._0646_ ),
    .A3(\u_cpu.IMEM._0583_ ),
    .B1(\u_cpu.IMEM._0103_ ),
    .C1(\u_cpu.IMEM._0900_ ),
    .X(\u_cpu.IMEM._0901_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1861_  (.A1(\u_cpu.IMEM._0897_ ),
    .A2(\u_cpu.IMEM._0898_ ),
    .B1(\u_cpu.IMEM._0302_ ),
    .C1(\u_cpu.IMEM._0901_ ),
    .Y(\u_cpu.IMEM._0902_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1862_  (.A1(\u_cpu.IMEM._0351_ ),
    .A2(\u_cpu.IMEM._0891_ ),
    .A3(\u_cpu.IMEM._0892_ ),
    .B1(\u_cpu.IMEM._0895_ ),
    .C1(\u_cpu.IMEM._0902_ ),
    .X(\u_cpu.IMEM._0903_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1863_  (.A1(\u_cpu.IMEM._0033_ ),
    .A2(\u_cpu.IMEM._0217_ ),
    .B1(\u_cpu.IMEM._0257_ ),
    .Y(\u_cpu.IMEM._0904_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1864_  (.A1(\u_cpu.IMEM._0445_ ),
    .A2(\u_cpu.IMEM._0298_ ),
    .A3(\u_cpu.IMEM._0782_ ),
    .B1(\u_cpu.IMEM._0904_ ),
    .C1(\u_cpu.IMEM._0237_ ),
    .X(\u_cpu.IMEM._0905_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu.IMEM._1865_  (.A1(\u_cpu.IMEM._0078_ ),
    .A2(\u_cpu.IMEM._0052_ ),
    .B1(\u_cpu.IMEM._0307_ ),
    .C1(\u_cpu.IMEM._0360_ ),
    .X(\u_cpu.IMEM._0906_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.IMEM._1866_  (.A1(\u_cpu.IMEM._0445_ ),
    .A2(\u_cpu.IMEM._0079_ ),
    .A3(\u_cpu.IMEM._0211_ ),
    .B1(\u_cpu.IMEM._0447_ ),
    .C1(\u_cpu.IMEM._0906_ ),
    .X(\u_cpu.IMEM._0907_ ));
 sky130_fd_sc_hd__o31a_2 \u_cpu.IMEM._1867_  (.A1(\u_cpu.IMEM._0173_ ),
    .A2(\u_cpu.IMEM._0905_ ),
    .A3(\u_cpu.IMEM._0907_ ),
    .B1(\u_cpu.IMEM._0628_ ),
    .X(\u_cpu.IMEM._0908_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.IMEM._1868_  (.A1(\u_cpu.IMEM._0512_ ),
    .A2(\u_cpu.IMEM._0168_ ),
    .A3(\u_cpu.IMEM._0158_ ),
    .B1(\u_cpu.IMEM._0062_ ),
    .C1(\u_cpu.IMEM._0200_ ),
    .Y(\u_cpu.IMEM._0909_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu.IMEM._1869_  (.A1(\u_cpu.IMEM._0348_ ),
    .A2(\u_cpu.IMEM._0234_ ),
    .A3(\u_cpu.IMEM._0586_ ),
    .B1(\u_cpu.IMEM._0028_ ),
    .B2(\u_cpu.IMEM._0909_ ),
    .X(\u_cpu.IMEM._0911_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1870_  (.A1(\u_cpu.IMEM._0117_ ),
    .A2(\u_cpu.IMEM._0911_ ),
    .B1(\u_cpu.IMEM._0431_ ),
    .Y(\u_cpu.IMEM._0912_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.IMEM._1871_  (.A1(\u_cpu.IMEM._0246_ ),
    .A2(\u_cpu.IMEM._0903_ ),
    .B1(\u_cpu.IMEM._0908_ ),
    .B2(\u_cpu.IMEM._0912_ ),
    .Y(\u_cpu.IMEM.rd[30] ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.IMEM._1872_  (.A1(\u_cpu.IMEM._0048_ ),
    .A2(\u_cpu.IMEM._0561_ ),
    .B1(\u_cpu.IMEM._0183_ ),
    .B2(\u_cpu.IMEM._0173_ ),
    .C1(\u_cpu.IMEM._0194_ ),
    .X(\u_cpu.IMEM._0913_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.IMEM._1873_  (.A1(\u_cpu.IMEM._0236_ ),
    .A2(\u_cpu.IMEM._0839_ ),
    .B1(\u_cpu.IMEM._0000_ ),
    .B2(\u_cpu.IMEM._0150_ ),
    .X(\u_cpu.IMEM._0914_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.IMEM._1874_  (.A1(\u_cpu.IMEM._0914_ ),
    .A2(\u_cpu.IMEM._0803_ ),
    .B1(\u_cpu.IMEM._0137_ ),
    .X(\u_cpu.IMEM._0915_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.IMEM._1875_  (.A1(\u_cpu.IMEM._0302_ ),
    .A2(\u_cpu.IMEM._0826_ ),
    .A3(\u_cpu.IMEM._0915_ ),
    .B1(\u_cpu.IMEM._0128_ ),
    .X(\u_cpu.IMEM._0916_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1876_  (.A1(\u_cpu.IMEM._0558_ ),
    .A2(\u_cpu.IMEM._0511_ ),
    .B1(\u_cpu.IMEM._0123_ ),
    .Y(\u_cpu.IMEM._0917_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.IMEM._1877_  (.A1(\u_cpu.IMEM._0262_ ),
    .A2(\u_cpu.IMEM._0425_ ),
    .B1(\u_cpu.IMEM._0917_ ),
    .Y(\u_cpu.IMEM._0918_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.IMEM._1878_  (.A1(\u_cpu.IMEM._0846_ ),
    .A2(\u_cpu.IMEM._0345_ ),
    .B1(\u_cpu.IMEM._0103_ ),
    .C1(\u_cpu.IMEM._0212_ ),
    .Y(\u_cpu.IMEM._0919_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu.IMEM._1879_  (.A1(\u_cpu.IMEM._0918_ ),
    .A2(\u_cpu.IMEM._0028_ ),
    .B1_N(\u_cpu.IMEM._0919_ ),
    .Y(\u_cpu.IMEM._0921_ ));
 sky130_fd_sc_hd__a32o_2 \u_cpu.IMEM._1880_  (.A1(\u_cpu.IMEM._0002_ ),
    .A2(\u_cpu.IMEM._0063_ ),
    .A3(\u_cpu.IMEM._0446_ ),
    .B1(\u_cpu.IMEM._0750_ ),
    .B2(\u_cpu.IMEM._0216_ ),
    .X(\u_cpu.IMEM._0922_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.IMEM._1881_  (.A1(\u_cpu.IMEM._0922_ ),
    .A2(\u_cpu.IMEM._0124_ ),
    .B1(\u_cpu.IMEM._0199_ ),
    .C1(\u_cpu.IMEM._0778_ ),
    .Y(\u_cpu.IMEM._0923_ ));
 sky130_fd_sc_hd__a2111o_2 \u_cpu.IMEM._1882_  (.A1(\u_cpu.IMEM._0013_ ),
    .A2(\u_cpu.IMEM._0411_ ),
    .B1(\u_cpu.IMEM._0434_ ),
    .C1(\u_cpu.IMEM._0046_ ),
    .D1(\u_cpu.IMEM._0052_ ),
    .X(\u_cpu.IMEM._0924_ ));
 sky130_fd_sc_hd__a41o_2 \u_cpu.IMEM._1883_  (.A1(\u_cpu.IMEM._0025_ ),
    .A2(\u_cpu.IMEM._0521_ ),
    .A3(\u_cpu.IMEM._0924_ ),
    .A4(\u_cpu.IMEM._0144_ ),
    .B1(\u_cpu.IMEM._0109_ ),
    .X(\u_cpu.IMEM._0925_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu.IMEM._1884_  (.A1(\u_cpu.IMEM._0194_ ),
    .A2(\u_cpu.IMEM._0921_ ),
    .B1(\u_cpu.IMEM._0923_ ),
    .B2(\u_cpu.IMEM._0925_ ),
    .X(\u_cpu.IMEM._0926_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.IMEM._1885_  (.A1(\u_cpu.IMEM._0913_ ),
    .A2(\u_cpu.IMEM._0916_ ),
    .B1(\u_cpu.IMEM._0246_ ),
    .B2(\u_cpu.IMEM._0926_ ),
    .Y(\u_cpu.IMEM.rd[31] ));
 sky130_fd_sc_hd__conb_1 \u_cpu.IMEM._1886_  (.HI(\u_cpu.IMEM.rd[0] ));
 sky130_fd_sc_hd__conb_1 \u_cpu.IMEM._1887_  (.HI(\u_cpu.IMEM.rd[1] ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05690_  (.A(\u_cpu.M_AXI_WDATA[19] ),
    .X(\u_cpu.REG_FILE._01024_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05691_  (.A(\u_cpu.REG_FILE._01024_ ),
    .X(\u_cpu.REG_FILE._01025_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05692_  (.A(\u_cpu.REG_FILE._01025_ ),
    .X(\u_cpu.REG_FILE._01026_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05693_  (.A(\u_cpu.M_AXI_WDATA[15] ),
    .X(\u_cpu.REG_FILE._01027_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05694_  (.A(\u_cpu.REG_FILE._01027_ ),
    .X(\u_cpu.REG_FILE._01028_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05695_  (.A(\u_cpu.REG_FILE._01028_ ),
    .X(\u_cpu.REG_FILE._01029_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05696_  (.A(\u_cpu.REG_FILE._01029_ ),
    .X(\u_cpu.REG_FILE._01030_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05697_  (.A(\u_cpu.M_AXI_WDATA[16] ),
    .X(\u_cpu.REG_FILE._01031_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05698_  (.A(\u_cpu.REG_FILE._01031_ ),
    .X(\u_cpu.REG_FILE._01032_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05699_  (.A(\u_cpu.REG_FILE._01032_ ),
    .X(\u_cpu.REG_FILE._01033_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05700_  (.A(\u_cpu.REG_FILE._01028_ ),
    .X(\u_cpu.REG_FILE._01034_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._05701_  (.A(\u_cpu.REG_FILE.rf[15][0] ),
    .B_N(\u_cpu.REG_FILE._01034_ ),
    .X(\u_cpu.REG_FILE._01035_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05702_  (.A1(\u_cpu.REG_FILE._01030_ ),
    .A2(\u_cpu.REG_FILE.rf[14][0] ),
    .B1(\u_cpu.REG_FILE._01033_ ),
    .C1(\u_cpu.REG_FILE._01035_ ),
    .Y(\u_cpu.REG_FILE._01036_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._05703_  (.A(\u_cpu.REG_FILE._01027_ ),
    .Y(\u_cpu.REG_FILE._01037_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05704_  (.A(\u_cpu.REG_FILE._01037_ ),
    .X(\u_cpu.REG_FILE._01038_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05705_  (.A(\u_cpu.REG_FILE._01038_ ),
    .X(\u_cpu.REG_FILE._01039_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05706_  (.A(\u_cpu.REG_FILE._01027_ ),
    .X(\u_cpu.REG_FILE._01040_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05707_  (.A(\u_cpu.REG_FILE._01040_ ),
    .X(\u_cpu.REG_FILE._01041_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05708_  (.A(\u_cpu.REG_FILE._01031_ ),
    .X(\u_cpu.REG_FILE._01042_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._05709_  (.A1(\u_cpu.REG_FILE._01041_ ),
    .A2(\u_cpu.REG_FILE.rf[12][0] ),
    .B1_N(\u_cpu.REG_FILE._01042_ ),
    .X(\u_cpu.REG_FILE._01043_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05710_  (.A1(\u_cpu.REG_FILE._01039_ ),
    .A2(\u_cpu.REG_FILE.rf[13][0] ),
    .B1(\u_cpu.REG_FILE._01043_ ),
    .Y(\u_cpu.REG_FILE._01044_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05711_  (.A(\u_cpu.M_AXI_WDATA[17] ),
    .X(\u_cpu.REG_FILE._01045_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05712_  (.A(\u_cpu.REG_FILE._01045_ ),
    .X(\u_cpu.REG_FILE._01046_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05713_  (.A(\u_cpu.REG_FILE._01046_ ),
    .X(\u_cpu.REG_FILE._01047_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._05714_  (.A(\u_cpu.REG_FILE._01036_ ),
    .B(\u_cpu.REG_FILE._01044_ ),
    .C(\u_cpu.REG_FILE._01047_ ),
    .Y(\u_cpu.REG_FILE._01048_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05715_  (.A(\u_cpu.REG_FILE._01027_ ),
    .X(\u_cpu.REG_FILE._01049_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05716_  (.A(\u_cpu.REG_FILE._01049_ ),
    .X(\u_cpu.REG_FILE._01050_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._05717_  (.A_N(\u_cpu.REG_FILE.rf[9][0] ),
    .B(\u_cpu.REG_FILE._01050_ ),
    .X(\u_cpu.REG_FILE._01051_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05718_  (.A(\u_cpu.REG_FILE._01040_ ),
    .X(\u_cpu.REG_FILE._01052_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05719_  (.A(\u_cpu.REG_FILE._01052_ ),
    .X(\u_cpu.REG_FILE._01053_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05720_  (.A(\u_cpu.M_AXI_WDATA[16] ),
    .X(\u_cpu.REG_FILE._01054_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05721_  (.A(\u_cpu.REG_FILE._01054_ ),
    .X(\u_cpu.REG_FILE._01055_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._05722_  (.A1(\u_cpu.REG_FILE._01053_ ),
    .A2(\u_cpu.REG_FILE.rf[8][0] ),
    .B1_N(\u_cpu.REG_FILE._01055_ ),
    .Y(\u_cpu.REG_FILE._01056_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._05723_  (.A(\u_cpu.REG_FILE._01045_ ),
    .Y(\u_cpu.REG_FILE._01057_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05724_  (.A(\u_cpu.REG_FILE._01057_ ),
    .X(\u_cpu.REG_FILE._01058_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05725_  (.A(\u_cpu.REG_FILE._01058_ ),
    .X(\u_cpu.REG_FILE._01059_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05726_  (.A(\u_cpu.REG_FILE._01040_ ),
    .X(\u_cpu.REG_FILE._01060_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05727_  (.A(\u_cpu.REG_FILE._01060_ ),
    .X(\u_cpu.REG_FILE._01061_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05728_  (.A(\u_cpu.REG_FILE._01031_ ),
    .X(\u_cpu.REG_FILE._01062_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05729_  (.A(\u_cpu.REG_FILE._01062_ ),
    .X(\u_cpu.REG_FILE._01063_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05730_  (.A(\u_cpu.REG_FILE._01027_ ),
    .X(\u_cpu.REG_FILE._01064_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05731_  (.A(\u_cpu.REG_FILE._01064_ ),
    .X(\u_cpu.REG_FILE._01065_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._05732_  (.A(\u_cpu.REG_FILE.rf[11][0] ),
    .B_N(\u_cpu.REG_FILE._01065_ ),
    .X(\u_cpu.REG_FILE._01066_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05733_  (.A1(\u_cpu.REG_FILE._01061_ ),
    .A2(\u_cpu.REG_FILE.rf[10][0] ),
    .B1(\u_cpu.REG_FILE._01063_ ),
    .C1(\u_cpu.REG_FILE._01066_ ),
    .Y(\u_cpu.REG_FILE._01067_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05734_  (.A1(\u_cpu.REG_FILE._01051_ ),
    .A2(\u_cpu.REG_FILE._01056_ ),
    .B1(\u_cpu.REG_FILE._01059_ ),
    .C1(\u_cpu.REG_FILE._01067_ ),
    .Y(\u_cpu.REG_FILE._01068_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05735_  (.A(\u_cpu.M_AXI_WDATA[18] ),
    .X(\u_cpu.REG_FILE._01069_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05736_  (.A(\u_cpu.REG_FILE._01069_ ),
    .X(\u_cpu.REG_FILE._01070_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._05737_  (.A(\u_cpu.REG_FILE._01048_ ),
    .B(\u_cpu.REG_FILE._01068_ ),
    .C(\u_cpu.REG_FILE._01070_ ),
    .Y(\u_cpu.REG_FILE._01071_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._05738_  (.A(\u_cpu.REG_FILE.rf[5][0] ),
    .Y(\u_cpu.REG_FILE._01072_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05739_  (.A(\u_cpu.REG_FILE._01027_ ),
    .X(\u_cpu.REG_FILE._01073_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05740_  (.A(\u_cpu.REG_FILE._01073_ ),
    .X(\u_cpu.REG_FILE._01074_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05741_  (.A(\u_cpu.REG_FILE._01074_ ),
    .X(\u_cpu.REG_FILE._01075_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05742_  (.A(\u_cpu.REG_FILE._01027_ ),
    .X(\u_cpu.REG_FILE._01076_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05743_  (.A(\u_cpu.REG_FILE._01076_ ),
    .X(\u_cpu.REG_FILE._01077_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05744_  (.A(\u_cpu.REG_FILE._01054_ ),
    .X(\u_cpu.REG_FILE._01078_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._05745_  (.A1(\u_cpu.REG_FILE._01077_ ),
    .A2(\u_cpu.REG_FILE.rf[4][0] ),
    .B1_N(\u_cpu.REG_FILE._01078_ ),
    .Y(\u_cpu.REG_FILE._01079_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._05746_  (.A1(\u_cpu.REG_FILE._01072_ ),
    .A2(\u_cpu.REG_FILE._01075_ ),
    .B1(\u_cpu.REG_FILE._01079_ ),
    .Y(\u_cpu.REG_FILE._01080_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05747_  (.A(\u_cpu.REG_FILE._01049_ ),
    .X(\u_cpu.REG_FILE._01081_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05748_  (.A(\u_cpu.M_AXI_WDATA[16] ),
    .X(\u_cpu.REG_FILE._01082_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05749_  (.A(\u_cpu.REG_FILE._01082_ ),
    .X(\u_cpu.REG_FILE._01083_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05750_  (.A1(\u_cpu.REG_FILE._01081_ ),
    .A2(\u_cpu.REG_FILE.rf[6][0] ),
    .B1(\u_cpu.REG_FILE._01083_ ),
    .Y(\u_cpu.REG_FILE._01084_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05751_  (.A(\u_cpu.REG_FILE._01073_ ),
    .X(\u_cpu.REG_FILE._01085_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._05752_  (.A_N(\u_cpu.REG_FILE.rf[7][0] ),
    .B(\u_cpu.REG_FILE._01085_ ),
    .X(\u_cpu.REG_FILE._01086_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05753_  (.A(\u_cpu.REG_FILE._01045_ ),
    .X(\u_cpu.REG_FILE._01087_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05754_  (.A1(\u_cpu.REG_FILE._01084_ ),
    .A2(\u_cpu.REG_FILE._01086_ ),
    .B1(\u_cpu.REG_FILE._01087_ ),
    .Y(\u_cpu.REG_FILE._01088_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._05755_  (.A(\u_cpu.M_AXI_WDATA[18] ),
    .Y(\u_cpu.REG_FILE._01089_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05756_  (.A(\u_cpu.REG_FILE._01089_ ),
    .X(\u_cpu.REG_FILE._01090_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05757_  (.A(\u_cpu.REG_FILE._01073_ ),
    .X(\u_cpu.REG_FILE._01091_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._05758_  (.A_N(\u_cpu.REG_FILE.rf[1][0] ),
    .B(\u_cpu.REG_FILE._01091_ ),
    .X(\u_cpu.REG_FILE._01092_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05759_  (.A(\u_cpu.REG_FILE._01052_ ),
    .X(\u_cpu.REG_FILE._01093_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05760_  (.A(\u_cpu.REG_FILE._01054_ ),
    .X(\u_cpu.REG_FILE._01094_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._05761_  (.A1(\u_cpu.REG_FILE.rf[0][0] ),
    .A2(\u_cpu.REG_FILE._01093_ ),
    .B1_N(\u_cpu.REG_FILE._01094_ ),
    .Y(\u_cpu.REG_FILE._01095_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05762_  (.A(\u_cpu.REG_FILE._01057_ ),
    .X(\u_cpu.REG_FILE._01096_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05763_  (.A(\u_cpu.REG_FILE._01052_ ),
    .X(\u_cpu.REG_FILE._01097_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05764_  (.A(\u_cpu.REG_FILE._01031_ ),
    .X(\u_cpu.REG_FILE._01098_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05765_  (.A(\u_cpu.REG_FILE._01098_ ),
    .X(\u_cpu.REG_FILE._01099_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._05766_  (.A(\u_cpu.REG_FILE.rf[3][0] ),
    .B_N(\u_cpu.REG_FILE._01060_ ),
    .X(\u_cpu.REG_FILE._01100_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05767_  (.A1(\u_cpu.REG_FILE._01097_ ),
    .A2(\u_cpu.REG_FILE.rf[2][0] ),
    .B1(\u_cpu.REG_FILE._01099_ ),
    .C1(\u_cpu.REG_FILE._01100_ ),
    .Y(\u_cpu.REG_FILE._01101_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05768_  (.A1(\u_cpu.REG_FILE._01092_ ),
    .A2(\u_cpu.REG_FILE._01095_ ),
    .B1(\u_cpu.REG_FILE._01096_ ),
    .C1(\u_cpu.REG_FILE._01101_ ),
    .Y(\u_cpu.REG_FILE._01102_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05769_  (.A1(\u_cpu.REG_FILE._01080_ ),
    .A2(\u_cpu.REG_FILE._01088_ ),
    .B1(\u_cpu.REG_FILE._01090_ ),
    .C1(\u_cpu.REG_FILE._01102_ ),
    .Y(\u_cpu.REG_FILE._01103_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._05770_  (.A(\u_cpu.REG_FILE._01071_ ),
    .B(\u_cpu.REG_FILE._01103_ ),
    .Y(\u_cpu.REG_FILE._01104_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05771_  (.A(\u_cpu.REG_FILE._01065_ ),
    .X(\u_cpu.REG_FILE._01105_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05772_  (.A(\u_cpu.M_AXI_WDATA[16] ),
    .X(\u_cpu.REG_FILE._01106_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05773_  (.A(\u_cpu.REG_FILE._01106_ ),
    .X(\u_cpu.REG_FILE._01107_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05774_  (.A(\u_cpu.REG_FILE._01064_ ),
    .X(\u_cpu.REG_FILE._01108_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._05775_  (.A(\u_cpu.REG_FILE.rf[27][0] ),
    .B_N(\u_cpu.REG_FILE._01108_ ),
    .X(\u_cpu.REG_FILE._01109_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._05776_  (.A1(\u_cpu.REG_FILE._01105_ ),
    .A2(\u_cpu.REG_FILE.rf[26][0] ),
    .B1(\u_cpu.REG_FILE._01107_ ),
    .C1(\u_cpu.REG_FILE._01109_ ),
    .X(\u_cpu.REG_FILE._01110_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05777_  (.A(\u_cpu.REG_FILE._01028_ ),
    .X(\u_cpu.REG_FILE._01111_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05778_  (.A(\u_cpu.REG_FILE._01031_ ),
    .X(\u_cpu.REG_FILE._01112_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._05779_  (.A1(\u_cpu.REG_FILE._01111_ ),
    .A2(\u_cpu.REG_FILE.rf[24][0] ),
    .B1_N(\u_cpu.REG_FILE._01112_ ),
    .X(\u_cpu.REG_FILE._01113_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._05780_  (.A(\u_cpu.REG_FILE.rf[25][0] ),
    .B_N(\u_cpu.REG_FILE._01029_ ),
    .X(\u_cpu.REG_FILE._01114_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05781_  (.A(\u_cpu.REG_FILE._01045_ ),
    .X(\u_cpu.REG_FILE._01115_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._05782_  (.A1(\u_cpu.REG_FILE._01113_ ),
    .A2(\u_cpu.REG_FILE._01114_ ),
    .B1(\u_cpu.REG_FILE._01115_ ),
    .X(\u_cpu.REG_FILE._01116_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05783_  (.A(\u_cpu.REG_FILE._01069_ ),
    .X(\u_cpu.REG_FILE._01117_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05784_  (.A(\u_cpu.REG_FILE._01065_ ),
    .X(\u_cpu.REG_FILE._01118_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._05785_  (.A(\u_cpu.REG_FILE._01118_ ),
    .B(\u_cpu.REG_FILE.rf[30][0] ),
    .Y(\u_cpu.REG_FILE._01119_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05786_  (.A(\u_cpu.REG_FILE._01037_ ),
    .X(\u_cpu.REG_FILE._01120_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05787_  (.A(\u_cpu.REG_FILE._01112_ ),
    .X(\u_cpu.REG_FILE._01121_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05788_  (.A1(\u_cpu.REG_FILE.rf[31][0] ),
    .A2(\u_cpu.REG_FILE._01120_ ),
    .B1(\u_cpu.REG_FILE._01121_ ),
    .Y(\u_cpu.REG_FILE._01122_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05789_  (.A(\u_cpu.REG_FILE._01037_ ),
    .X(\u_cpu.REG_FILE._01123_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05790_  (.A(\u_cpu.REG_FILE._01123_ ),
    .X(\u_cpu.REG_FILE._01124_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05791_  (.A(\u_cpu.REG_FILE._01028_ ),
    .X(\u_cpu.REG_FILE._01125_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05792_  (.A(\u_cpu.REG_FILE._01031_ ),
    .X(\u_cpu.REG_FILE._01126_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._05793_  (.A1(\u_cpu.REG_FILE._01125_ ),
    .A2(\u_cpu.REG_FILE.rf[28][0] ),
    .B1_N(\u_cpu.REG_FILE._01126_ ),
    .X(\u_cpu.REG_FILE._01127_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05794_  (.A1(\u_cpu.REG_FILE._01124_ ),
    .A2(\u_cpu.REG_FILE.rf[29][0] ),
    .B1(\u_cpu.REG_FILE._01127_ ),
    .Y(\u_cpu.REG_FILE._01128_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05795_  (.A(\u_cpu.REG_FILE._01046_ ),
    .X(\u_cpu.REG_FILE._01129_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05796_  (.A1(\u_cpu.REG_FILE._01119_ ),
    .A2(\u_cpu.REG_FILE._01122_ ),
    .B1(\u_cpu.REG_FILE._01128_ ),
    .C1(\u_cpu.REG_FILE._01129_ ),
    .Y(\u_cpu.REG_FILE._01130_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05797_  (.A1(\u_cpu.REG_FILE._01110_ ),
    .A2(\u_cpu.REG_FILE._01116_ ),
    .B1(\u_cpu.REG_FILE._01117_ ),
    .C1(\u_cpu.REG_FILE._01130_ ),
    .Y(\u_cpu.REG_FILE._01131_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05798_  (.A(\u_cpu.REG_FILE._01089_ ),
    .X(\u_cpu.REG_FILE._01132_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05799_  (.A(\u_cpu.REG_FILE._01076_ ),
    .X(\u_cpu.REG_FILE._01133_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05800_  (.A(\u_cpu.M_AXI_WDATA[16] ),
    .X(\u_cpu.REG_FILE._01134_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05801_  (.A(\u_cpu.REG_FILE._01134_ ),
    .X(\u_cpu.REG_FILE._01135_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05802_  (.A1(\u_cpu.REG_FILE._01133_ ),
    .A2(\u_cpu.REG_FILE.rf[18][0] ),
    .B1(\u_cpu.REG_FILE._01135_ ),
    .Y(\u_cpu.REG_FILE._01136_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05803_  (.A(\u_cpu.REG_FILE._01123_ ),
    .X(\u_cpu.REG_FILE._01137_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._05804_  (.A(\u_cpu.REG_FILE.rf[19][0] ),
    .B(\u_cpu.REG_FILE._01137_ ),
    .Y(\u_cpu.REG_FILE._01138_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05805_  (.A(\u_cpu.REG_FILE._01057_ ),
    .X(\u_cpu.REG_FILE._01139_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05806_  (.A(\u_cpu.REG_FILE._01123_ ),
    .X(\u_cpu.REG_FILE._01140_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05807_  (.A(\u_cpu.REG_FILE._01064_ ),
    .X(\u_cpu.REG_FILE._01141_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05808_  (.A(\u_cpu.M_AXI_WDATA[16] ),
    .X(\u_cpu.REG_FILE._01142_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._05809_  (.A1(\u_cpu.REG_FILE._01141_ ),
    .A2(\u_cpu.REG_FILE.rf[16][0] ),
    .B1_N(\u_cpu.REG_FILE._01142_ ),
    .X(\u_cpu.REG_FILE._01143_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05810_  (.A1(\u_cpu.REG_FILE._01140_ ),
    .A2(\u_cpu.REG_FILE.rf[17][0] ),
    .B1(\u_cpu.REG_FILE._01143_ ),
    .Y(\u_cpu.REG_FILE._01144_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05811_  (.A1(\u_cpu.REG_FILE._01136_ ),
    .A2(\u_cpu.REG_FILE._01138_ ),
    .B1(\u_cpu.REG_FILE._01139_ ),
    .C1(\u_cpu.REG_FILE._01144_ ),
    .Y(\u_cpu.REG_FILE._01145_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05812_  (.A(\u_cpu.REG_FILE._01037_ ),
    .X(\u_cpu.REG_FILE._01146_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05813_  (.A(\u_cpu.REG_FILE._01062_ ),
    .X(\u_cpu.REG_FILE._01147_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05814_  (.A(\u_cpu.REG_FILE._01027_ ),
    .X(\u_cpu.REG_FILE._01148_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._05815_  (.A(\u_cpu.REG_FILE._01148_ ),
    .B(\u_cpu.REG_FILE.rf[22][0] ),
    .X(\u_cpu.REG_FILE._01149_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05816_  (.A1(\u_cpu.REG_FILE._01146_ ),
    .A2(\u_cpu.REG_FILE.rf[23][0] ),
    .B1(\u_cpu.REG_FILE._01147_ ),
    .C1(\u_cpu.REG_FILE._01149_ ),
    .Y(\u_cpu.REG_FILE._01150_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05817_  (.A(\u_cpu.REG_FILE._01037_ ),
    .X(\u_cpu.REG_FILE._01151_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05818_  (.A(\u_cpu.REG_FILE._01064_ ),
    .X(\u_cpu.REG_FILE._01152_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05819_  (.A(\u_cpu.REG_FILE._01031_ ),
    .X(\u_cpu.REG_FILE._01153_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._05820_  (.A1(\u_cpu.REG_FILE._01152_ ),
    .A2(\u_cpu.REG_FILE.rf[20][0] ),
    .B1_N(\u_cpu.REG_FILE._01153_ ),
    .X(\u_cpu.REG_FILE._01154_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05821_  (.A1(\u_cpu.REG_FILE._01151_ ),
    .A2(\u_cpu.REG_FILE.rf[21][0] ),
    .B1(\u_cpu.REG_FILE._01154_ ),
    .Y(\u_cpu.REG_FILE._01155_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05822_  (.A(\u_cpu.REG_FILE._01045_ ),
    .X(\u_cpu.REG_FILE._01156_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._05823_  (.A(\u_cpu.REG_FILE._01150_ ),
    .B(\u_cpu.REG_FILE._01155_ ),
    .C(\u_cpu.REG_FILE._01156_ ),
    .Y(\u_cpu.REG_FILE._01157_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._05824_  (.A(\u_cpu.REG_FILE._01132_ ),
    .B(\u_cpu.REG_FILE._01145_ ),
    .C(\u_cpu.REG_FILE._01157_ ),
    .Y(\u_cpu.REG_FILE._01158_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05825_  (.A(\u_cpu.REG_FILE._01024_ ),
    .X(\u_cpu.REG_FILE._01159_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._05826_  (.A(\u_cpu.REG_FILE._01131_ ),
    .B(\u_cpu.REG_FILE._01158_ ),
    .C(\u_cpu.REG_FILE._01159_ ),
    .Y(\u_cpu.REG_FILE._01160_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05827_  (.A(\u_cpu.REG_FILE._01073_ ),
    .X(\u_cpu.REG_FILE._01161_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.REG_FILE._05828_  (.A(\u_cpu.M_AXI_WDATA[16] ),
    .B(\u_cpu.REG_FILE._01045_ ),
    .C(\u_cpu.M_AXI_WDATA[18] ),
    .X(\u_cpu.REG_FILE._01162_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.REG_FILE._05829_  (.A(\u_cpu.M_AXI_WDATA[19] ),
    .B(\u_cpu.REG_FILE._01161_ ),
    .C(\u_cpu.REG_FILE._01162_ ),
    .X(\u_cpu.REG_FILE._01163_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05830_  (.A(\u_cpu.REG_FILE._01163_ ),
    .X(\u_cpu.REG_FILE._01164_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05831_  (.A(\u_cpu.REG_FILE._01164_ ),
    .X(\u_cpu.REG_FILE._01165_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._05832_  (.A1(\u_cpu.REG_FILE._01026_ ),
    .A2(\u_cpu.REG_FILE._01104_ ),
    .B1(\u_cpu.REG_FILE._01160_ ),
    .C1(\u_cpu.REG_FILE._01165_ ),
    .X(\u_cpu.ALU.SrcA[0] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._05833_  (.A(\u_cpu.REG_FILE.rf[15][1] ),
    .B_N(\u_cpu.REG_FILE._01034_ ),
    .X(\u_cpu.REG_FILE._01166_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05834_  (.A1(\u_cpu.REG_FILE._01030_ ),
    .A2(\u_cpu.REG_FILE.rf[14][1] ),
    .B1(\u_cpu.REG_FILE._01033_ ),
    .C1(\u_cpu.REG_FILE._01166_ ),
    .Y(\u_cpu.REG_FILE._01167_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._05835_  (.A1(\u_cpu.REG_FILE._01041_ ),
    .A2(\u_cpu.REG_FILE.rf[12][1] ),
    .B1_N(\u_cpu.REG_FILE._01042_ ),
    .X(\u_cpu.REG_FILE._01168_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05836_  (.A1(\u_cpu.REG_FILE._01039_ ),
    .A2(\u_cpu.REG_FILE.rf[13][1] ),
    .B1(\u_cpu.REG_FILE._01168_ ),
    .Y(\u_cpu.REG_FILE._01169_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._05837_  (.A(\u_cpu.REG_FILE._01167_ ),
    .B(\u_cpu.REG_FILE._01169_ ),
    .C(\u_cpu.REG_FILE._01047_ ),
    .Y(\u_cpu.REG_FILE._01170_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._05838_  (.A_N(\u_cpu.REG_FILE.rf[9][1] ),
    .B(\u_cpu.REG_FILE._01050_ ),
    .X(\u_cpu.REG_FILE._01171_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._05839_  (.A1(\u_cpu.REG_FILE._01053_ ),
    .A2(\u_cpu.REG_FILE.rf[8][1] ),
    .B1_N(\u_cpu.REG_FILE._01055_ ),
    .Y(\u_cpu.REG_FILE._01172_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._05840_  (.A(\u_cpu.REG_FILE.rf[11][1] ),
    .B_N(\u_cpu.REG_FILE._01065_ ),
    .X(\u_cpu.REG_FILE._01173_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05841_  (.A1(\u_cpu.REG_FILE._01061_ ),
    .A2(\u_cpu.REG_FILE.rf[10][1] ),
    .B1(\u_cpu.REG_FILE._01063_ ),
    .C1(\u_cpu.REG_FILE._01173_ ),
    .Y(\u_cpu.REG_FILE._01174_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05842_  (.A1(\u_cpu.REG_FILE._01171_ ),
    .A2(\u_cpu.REG_FILE._01172_ ),
    .B1(\u_cpu.REG_FILE._01059_ ),
    .C1(\u_cpu.REG_FILE._01174_ ),
    .Y(\u_cpu.REG_FILE._01175_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._05843_  (.A(\u_cpu.REG_FILE._01170_ ),
    .B(\u_cpu.REG_FILE._01175_ ),
    .C(\u_cpu.REG_FILE._01070_ ),
    .Y(\u_cpu.REG_FILE._01176_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._05844_  (.A(\u_cpu.REG_FILE.rf[5][1] ),
    .Y(\u_cpu.REG_FILE._01177_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._05845_  (.A1(\u_cpu.REG_FILE._01077_ ),
    .A2(\u_cpu.REG_FILE.rf[4][1] ),
    .B1_N(\u_cpu.REG_FILE._01078_ ),
    .Y(\u_cpu.REG_FILE._01178_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._05846_  (.A1(\u_cpu.REG_FILE._01177_ ),
    .A2(\u_cpu.REG_FILE._01075_ ),
    .B1(\u_cpu.REG_FILE._01178_ ),
    .Y(\u_cpu.REG_FILE._01179_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05847_  (.A1(\u_cpu.REG_FILE._01081_ ),
    .A2(\u_cpu.REG_FILE.rf[6][1] ),
    .B1(\u_cpu.REG_FILE._01083_ ),
    .Y(\u_cpu.REG_FILE._01180_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._05848_  (.A_N(\u_cpu.REG_FILE.rf[7][1] ),
    .B(\u_cpu.REG_FILE._01085_ ),
    .X(\u_cpu.REG_FILE._01181_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05849_  (.A1(\u_cpu.REG_FILE._01180_ ),
    .A2(\u_cpu.REG_FILE._01181_ ),
    .B1(\u_cpu.REG_FILE._01087_ ),
    .Y(\u_cpu.REG_FILE._01182_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._05850_  (.A_N(\u_cpu.REG_FILE.rf[1][1] ),
    .B(\u_cpu.REG_FILE._01091_ ),
    .X(\u_cpu.REG_FILE._01183_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05851_  (.A(\u_cpu.REG_FILE._01076_ ),
    .X(\u_cpu.REG_FILE._01184_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._05852_  (.A1(\u_cpu.REG_FILE._01184_ ),
    .A2(\u_cpu.REG_FILE.rf[0][1] ),
    .B1_N(\u_cpu.REG_FILE._01094_ ),
    .Y(\u_cpu.REG_FILE._01185_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._05853_  (.A(\u_cpu.REG_FILE.rf[3][1] ),
    .B_N(\u_cpu.REG_FILE._01060_ ),
    .X(\u_cpu.REG_FILE._01186_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05854_  (.A1(\u_cpu.REG_FILE._01097_ ),
    .A2(\u_cpu.REG_FILE.rf[2][1] ),
    .B1(\u_cpu.REG_FILE._01099_ ),
    .C1(\u_cpu.REG_FILE._01186_ ),
    .Y(\u_cpu.REG_FILE._01187_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05855_  (.A1(\u_cpu.REG_FILE._01183_ ),
    .A2(\u_cpu.REG_FILE._01185_ ),
    .B1(\u_cpu.REG_FILE._01096_ ),
    .C1(\u_cpu.REG_FILE._01187_ ),
    .Y(\u_cpu.REG_FILE._01188_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05856_  (.A1(\u_cpu.REG_FILE._01179_ ),
    .A2(\u_cpu.REG_FILE._01182_ ),
    .B1(\u_cpu.REG_FILE._01090_ ),
    .C1(\u_cpu.REG_FILE._01188_ ),
    .Y(\u_cpu.REG_FILE._01189_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._05857_  (.A(\u_cpu.REG_FILE._01176_ ),
    .B(\u_cpu.REG_FILE._01189_ ),
    .Y(\u_cpu.REG_FILE._01190_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._05858_  (.A(\u_cpu.REG_FILE.rf[27][1] ),
    .B_N(\u_cpu.REG_FILE._01108_ ),
    .X(\u_cpu.REG_FILE._01191_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._05859_  (.A1(\u_cpu.REG_FILE._01105_ ),
    .A2(\u_cpu.REG_FILE.rf[26][1] ),
    .B1(\u_cpu.REG_FILE._01107_ ),
    .C1(\u_cpu.REG_FILE._01191_ ),
    .X(\u_cpu.REG_FILE._01192_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._05860_  (.A1(\u_cpu.REG_FILE._01111_ ),
    .A2(\u_cpu.REG_FILE.rf[24][1] ),
    .B1_N(\u_cpu.REG_FILE._01112_ ),
    .X(\u_cpu.REG_FILE._01193_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05861_  (.A(\u_cpu.REG_FILE._01064_ ),
    .X(\u_cpu.REG_FILE._01194_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._05862_  (.A(\u_cpu.REG_FILE.rf[25][1] ),
    .B_N(\u_cpu.REG_FILE._01194_ ),
    .X(\u_cpu.REG_FILE._01195_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05863_  (.A(\u_cpu.REG_FILE._01045_ ),
    .X(\u_cpu.REG_FILE._01196_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._05864_  (.A1(\u_cpu.REG_FILE._01193_ ),
    .A2(\u_cpu.REG_FILE._01195_ ),
    .B1(\u_cpu.REG_FILE._01196_ ),
    .X(\u_cpu.REG_FILE._01197_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05865_  (.A(\u_cpu.REG_FILE._01069_ ),
    .X(\u_cpu.REG_FILE._01198_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._05866_  (.A(\u_cpu.REG_FILE._01118_ ),
    .B(\u_cpu.REG_FILE.rf[30][1] ),
    .Y(\u_cpu.REG_FILE._01199_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05867_  (.A(\u_cpu.REG_FILE._01123_ ),
    .X(\u_cpu.REG_FILE._01200_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05868_  (.A1(\u_cpu.REG_FILE.rf[31][1] ),
    .A2(\u_cpu.REG_FILE._01200_ ),
    .B1(\u_cpu.REG_FILE._01121_ ),
    .Y(\u_cpu.REG_FILE._01201_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._05869_  (.A1(\u_cpu.REG_FILE._01125_ ),
    .A2(\u_cpu.REG_FILE.rf[28][1] ),
    .B1_N(\u_cpu.REG_FILE._01126_ ),
    .X(\u_cpu.REG_FILE._01202_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05870_  (.A1(\u_cpu.REG_FILE._01124_ ),
    .A2(\u_cpu.REG_FILE.rf[29][1] ),
    .B1(\u_cpu.REG_FILE._01202_ ),
    .Y(\u_cpu.REG_FILE._01203_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05871_  (.A1(\u_cpu.REG_FILE._01199_ ),
    .A2(\u_cpu.REG_FILE._01201_ ),
    .B1(\u_cpu.REG_FILE._01203_ ),
    .C1(\u_cpu.REG_FILE._01129_ ),
    .Y(\u_cpu.REG_FILE._01204_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05872_  (.A1(\u_cpu.REG_FILE._01192_ ),
    .A2(\u_cpu.REG_FILE._01197_ ),
    .B1(\u_cpu.REG_FILE._01198_ ),
    .C1(\u_cpu.REG_FILE._01204_ ),
    .Y(\u_cpu.REG_FILE._01205_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05873_  (.A(\u_cpu.REG_FILE._01076_ ),
    .X(\u_cpu.REG_FILE._01206_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05874_  (.A1(\u_cpu.REG_FILE._01206_ ),
    .A2(\u_cpu.REG_FILE.rf[18][1] ),
    .B1(\u_cpu.REG_FILE._01135_ ),
    .Y(\u_cpu.REG_FILE._01207_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._05875_  (.A(\u_cpu.REG_FILE.rf[19][1] ),
    .B(\u_cpu.REG_FILE._01137_ ),
    .Y(\u_cpu.REG_FILE._01208_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._05876_  (.A1(\u_cpu.REG_FILE._01141_ ),
    .A2(\u_cpu.REG_FILE.rf[16][1] ),
    .B1_N(\u_cpu.REG_FILE._01142_ ),
    .X(\u_cpu.REG_FILE._01209_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05877_  (.A1(\u_cpu.REG_FILE._01140_ ),
    .A2(\u_cpu.REG_FILE.rf[17][1] ),
    .B1(\u_cpu.REG_FILE._01209_ ),
    .Y(\u_cpu.REG_FILE._01210_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05878_  (.A1(\u_cpu.REG_FILE._01207_ ),
    .A2(\u_cpu.REG_FILE._01208_ ),
    .B1(\u_cpu.REG_FILE._01139_ ),
    .C1(\u_cpu.REG_FILE._01210_ ),
    .Y(\u_cpu.REG_FILE._01211_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._05879_  (.A(\u_cpu.REG_FILE._01148_ ),
    .B(\u_cpu.REG_FILE.rf[22][1] ),
    .X(\u_cpu.REG_FILE._01212_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05880_  (.A1(\u_cpu.REG_FILE._01146_ ),
    .A2(\u_cpu.REG_FILE.rf[23][1] ),
    .B1(\u_cpu.REG_FILE._01147_ ),
    .C1(\u_cpu.REG_FILE._01212_ ),
    .Y(\u_cpu.REG_FILE._01213_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05881_  (.A(\u_cpu.M_AXI_WDATA[16] ),
    .X(\u_cpu.REG_FILE._01214_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._05882_  (.A1(\u_cpu.REG_FILE._01152_ ),
    .A2(\u_cpu.REG_FILE.rf[20][1] ),
    .B1_N(\u_cpu.REG_FILE._01214_ ),
    .X(\u_cpu.REG_FILE._01215_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05883_  (.A1(\u_cpu.REG_FILE._01151_ ),
    .A2(\u_cpu.REG_FILE.rf[21][1] ),
    .B1(\u_cpu.REG_FILE._01215_ ),
    .Y(\u_cpu.REG_FILE._01216_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._05884_  (.A(\u_cpu.REG_FILE._01213_ ),
    .B(\u_cpu.REG_FILE._01216_ ),
    .C(\u_cpu.REG_FILE._01156_ ),
    .Y(\u_cpu.REG_FILE._01217_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._05885_  (.A(\u_cpu.REG_FILE._01132_ ),
    .B(\u_cpu.REG_FILE._01211_ ),
    .C(\u_cpu.REG_FILE._01217_ ),
    .Y(\u_cpu.REG_FILE._01218_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._05886_  (.A(\u_cpu.REG_FILE._01205_ ),
    .B(\u_cpu.REG_FILE._01218_ ),
    .C(\u_cpu.REG_FILE._01159_ ),
    .Y(\u_cpu.REG_FILE._01219_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._05887_  (.A1(\u_cpu.REG_FILE._01026_ ),
    .A2(\u_cpu.REG_FILE._01190_ ),
    .B1(\u_cpu.REG_FILE._01219_ ),
    .C1(\u_cpu.REG_FILE._01165_ ),
    .X(\u_cpu.ALU.SrcA[1] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._05888_  (.A(\u_cpu.REG_FILE.rf[15][2] ),
    .B_N(\u_cpu.REG_FILE._01034_ ),
    .X(\u_cpu.REG_FILE._01220_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05889_  (.A1(\u_cpu.REG_FILE._01030_ ),
    .A2(\u_cpu.REG_FILE.rf[14][2] ),
    .B1(\u_cpu.REG_FILE._01033_ ),
    .C1(\u_cpu.REG_FILE._01220_ ),
    .Y(\u_cpu.REG_FILE._01221_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._05890_  (.A1(\u_cpu.REG_FILE._01041_ ),
    .A2(\u_cpu.REG_FILE.rf[12][2] ),
    .B1_N(\u_cpu.REG_FILE._01042_ ),
    .X(\u_cpu.REG_FILE._01222_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05891_  (.A1(\u_cpu.REG_FILE._01039_ ),
    .A2(\u_cpu.REG_FILE.rf[13][2] ),
    .B1(\u_cpu.REG_FILE._01222_ ),
    .Y(\u_cpu.REG_FILE._01223_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._05892_  (.A(\u_cpu.REG_FILE._01221_ ),
    .B(\u_cpu.REG_FILE._01223_ ),
    .C(\u_cpu.REG_FILE._01047_ ),
    .Y(\u_cpu.REG_FILE._01224_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._05893_  (.A_N(\u_cpu.REG_FILE.rf[9][2] ),
    .B(\u_cpu.REG_FILE._01050_ ),
    .X(\u_cpu.REG_FILE._01225_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._05894_  (.A1(\u_cpu.REG_FILE._01053_ ),
    .A2(\u_cpu.REG_FILE.rf[8][2] ),
    .B1_N(\u_cpu.REG_FILE._01055_ ),
    .Y(\u_cpu.REG_FILE._01226_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._05895_  (.A(\u_cpu.REG_FILE.rf[11][2] ),
    .B_N(\u_cpu.REG_FILE._01065_ ),
    .X(\u_cpu.REG_FILE._01227_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05896_  (.A1(\u_cpu.REG_FILE._01061_ ),
    .A2(\u_cpu.REG_FILE.rf[10][2] ),
    .B1(\u_cpu.REG_FILE._01063_ ),
    .C1(\u_cpu.REG_FILE._01227_ ),
    .Y(\u_cpu.REG_FILE._01228_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05897_  (.A1(\u_cpu.REG_FILE._01225_ ),
    .A2(\u_cpu.REG_FILE._01226_ ),
    .B1(\u_cpu.REG_FILE._01059_ ),
    .C1(\u_cpu.REG_FILE._01228_ ),
    .Y(\u_cpu.REG_FILE._01229_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._05898_  (.A(\u_cpu.REG_FILE._01224_ ),
    .B(\u_cpu.REG_FILE._01229_ ),
    .C(\u_cpu.REG_FILE._01070_ ),
    .Y(\u_cpu.REG_FILE._01230_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._05899_  (.A(\u_cpu.REG_FILE.rf[5][2] ),
    .Y(\u_cpu.REG_FILE._01231_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._05900_  (.A1(\u_cpu.REG_FILE._01077_ ),
    .A2(\u_cpu.REG_FILE.rf[4][2] ),
    .B1_N(\u_cpu.REG_FILE._01078_ ),
    .Y(\u_cpu.REG_FILE._01232_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._05901_  (.A1(\u_cpu.REG_FILE._01231_ ),
    .A2(\u_cpu.REG_FILE._01075_ ),
    .B1(\u_cpu.REG_FILE._01232_ ),
    .Y(\u_cpu.REG_FILE._01233_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05902_  (.A1(\u_cpu.REG_FILE._01081_ ),
    .A2(\u_cpu.REG_FILE.rf[6][2] ),
    .B1(\u_cpu.REG_FILE._01083_ ),
    .Y(\u_cpu.REG_FILE._01234_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._05903_  (.A_N(\u_cpu.REG_FILE.rf[7][2] ),
    .B(\u_cpu.REG_FILE._01085_ ),
    .X(\u_cpu.REG_FILE._01235_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05904_  (.A1(\u_cpu.REG_FILE._01234_ ),
    .A2(\u_cpu.REG_FILE._01235_ ),
    .B1(\u_cpu.REG_FILE._01087_ ),
    .Y(\u_cpu.REG_FILE._01236_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._05905_  (.A_N(\u_cpu.REG_FILE.rf[1][2] ),
    .B(\u_cpu.REG_FILE._01091_ ),
    .X(\u_cpu.REG_FILE._01237_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._05906_  (.A1(\u_cpu.REG_FILE._01184_ ),
    .A2(\u_cpu.REG_FILE.rf[0][2] ),
    .B1_N(\u_cpu.REG_FILE._01094_ ),
    .Y(\u_cpu.REG_FILE._01238_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05907_  (.A(\u_cpu.REG_FILE._01031_ ),
    .X(\u_cpu.REG_FILE._01239_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05908_  (.A(\u_cpu.REG_FILE._01239_ ),
    .X(\u_cpu.REG_FILE._01240_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05909_  (.A(\u_cpu.REG_FILE._01040_ ),
    .X(\u_cpu.REG_FILE._01241_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._05910_  (.A(\u_cpu.REG_FILE.rf[3][2] ),
    .B_N(\u_cpu.REG_FILE._01241_ ),
    .X(\u_cpu.REG_FILE._01242_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05911_  (.A1(\u_cpu.REG_FILE._01097_ ),
    .A2(\u_cpu.REG_FILE.rf[2][2] ),
    .B1(\u_cpu.REG_FILE._01240_ ),
    .C1(\u_cpu.REG_FILE._01242_ ),
    .Y(\u_cpu.REG_FILE._01243_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05912_  (.A1(\u_cpu.REG_FILE._01237_ ),
    .A2(\u_cpu.REG_FILE._01238_ ),
    .B1(\u_cpu.REG_FILE._01096_ ),
    .C1(\u_cpu.REG_FILE._01243_ ),
    .Y(\u_cpu.REG_FILE._01244_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05913_  (.A1(\u_cpu.REG_FILE._01233_ ),
    .A2(\u_cpu.REG_FILE._01236_ ),
    .B1(\u_cpu.REG_FILE._01090_ ),
    .C1(\u_cpu.REG_FILE._01244_ ),
    .Y(\u_cpu.REG_FILE._01245_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._05914_  (.A(\u_cpu.REG_FILE._01230_ ),
    .B(\u_cpu.REG_FILE._01245_ ),
    .Y(\u_cpu.REG_FILE._01246_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._05915_  (.A(\u_cpu.REG_FILE.rf[27][2] ),
    .B_N(\u_cpu.REG_FILE._01108_ ),
    .X(\u_cpu.REG_FILE._01247_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._05916_  (.A1(\u_cpu.REG_FILE._01105_ ),
    .A2(\u_cpu.REG_FILE.rf[26][2] ),
    .B1(\u_cpu.REG_FILE._01107_ ),
    .C1(\u_cpu.REG_FILE._01247_ ),
    .X(\u_cpu.REG_FILE._01248_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._05917_  (.A1(\u_cpu.REG_FILE._01111_ ),
    .A2(\u_cpu.REG_FILE.rf[24][2] ),
    .B1_N(\u_cpu.REG_FILE._01112_ ),
    .X(\u_cpu.REG_FILE._01249_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._05918_  (.A(\u_cpu.REG_FILE.rf[25][2] ),
    .B_N(\u_cpu.REG_FILE._01194_ ),
    .X(\u_cpu.REG_FILE._01250_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._05919_  (.A1(\u_cpu.REG_FILE._01249_ ),
    .A2(\u_cpu.REG_FILE._01250_ ),
    .B1(\u_cpu.REG_FILE._01196_ ),
    .X(\u_cpu.REG_FILE._01251_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._05920_  (.A(\u_cpu.REG_FILE._01118_ ),
    .B(\u_cpu.REG_FILE.rf[30][2] ),
    .Y(\u_cpu.REG_FILE._01252_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05921_  (.A1(\u_cpu.REG_FILE.rf[31][2] ),
    .A2(\u_cpu.REG_FILE._01200_ ),
    .B1(\u_cpu.REG_FILE._01121_ ),
    .Y(\u_cpu.REG_FILE._01253_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._05922_  (.A1(\u_cpu.REG_FILE._01125_ ),
    .A2(\u_cpu.REG_FILE.rf[28][2] ),
    .B1_N(\u_cpu.REG_FILE._01126_ ),
    .X(\u_cpu.REG_FILE._01254_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05923_  (.A1(\u_cpu.REG_FILE._01124_ ),
    .A2(\u_cpu.REG_FILE.rf[29][2] ),
    .B1(\u_cpu.REG_FILE._01254_ ),
    .Y(\u_cpu.REG_FILE._01255_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05924_  (.A1(\u_cpu.REG_FILE._01252_ ),
    .A2(\u_cpu.REG_FILE._01253_ ),
    .B1(\u_cpu.REG_FILE._01255_ ),
    .C1(\u_cpu.REG_FILE._01129_ ),
    .Y(\u_cpu.REG_FILE._01256_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05925_  (.A1(\u_cpu.REG_FILE._01248_ ),
    .A2(\u_cpu.REG_FILE._01251_ ),
    .B1(\u_cpu.REG_FILE._01198_ ),
    .C1(\u_cpu.REG_FILE._01256_ ),
    .Y(\u_cpu.REG_FILE._01257_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05926_  (.A(\u_cpu.REG_FILE._01054_ ),
    .X(\u_cpu.REG_FILE._01258_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05927_  (.A(\u_cpu.REG_FILE._01258_ ),
    .X(\u_cpu.REG_FILE._01259_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05928_  (.A(\u_cpu.REG_FILE._01076_ ),
    .X(\u_cpu.REG_FILE._01260_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._05929_  (.A(\u_cpu.REG_FILE._01260_ ),
    .B(\u_cpu.REG_FILE.rf[16][2] ),
    .Y(\u_cpu.REG_FILE._01261_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05930_  (.A(\u_cpu.REG_FILE._01028_ ),
    .X(\u_cpu.REG_FILE._01262_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._05931_  (.A_N(\u_cpu.REG_FILE.rf[17][2] ),
    .B(\u_cpu.REG_FILE._01262_ ),
    .X(\u_cpu.REG_FILE._01263_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05932_  (.A(\u_cpu.REG_FILE._01057_ ),
    .X(\u_cpu.REG_FILE._01264_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05933_  (.A(\u_cpu.REG_FILE._01037_ ),
    .X(\u_cpu.REG_FILE._01265_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.REG_FILE._05934_  (.A1(\u_cpu.REG_FILE._01060_ ),
    .A2(\u_cpu.REG_FILE.rf[18][2] ),
    .B1(\u_cpu.REG_FILE._01239_ ),
    .X(\u_cpu.REG_FILE._01266_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05935_  (.A1(\u_cpu.REG_FILE.rf[19][2] ),
    .A2(\u_cpu.REG_FILE._01265_ ),
    .B1(\u_cpu.REG_FILE._01266_ ),
    .Y(\u_cpu.REG_FILE._01267_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._05936_  (.A1(\u_cpu.REG_FILE._01259_ ),
    .A2(\u_cpu.REG_FILE._01261_ ),
    .A3(\u_cpu.REG_FILE._01263_ ),
    .B1(\u_cpu.REG_FILE._01264_ ),
    .C1(\u_cpu.REG_FILE._01267_ ),
    .Y(\u_cpu.REG_FILE._01268_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05937_  (.A(\u_cpu.REG_FILE._01040_ ),
    .X(\u_cpu.REG_FILE._01269_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._05938_  (.A(\u_cpu.REG_FILE._01269_ ),
    .B(\u_cpu.REG_FILE.rf[22][2] ),
    .X(\u_cpu.REG_FILE._01270_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05939_  (.A1(\u_cpu.REG_FILE._01146_ ),
    .A2(\u_cpu.REG_FILE.rf[23][2] ),
    .B1(\u_cpu.REG_FILE._01147_ ),
    .C1(\u_cpu.REG_FILE._01270_ ),
    .Y(\u_cpu.REG_FILE._01271_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._05940_  (.A1(\u_cpu.REG_FILE._01152_ ),
    .A2(\u_cpu.REG_FILE.rf[20][2] ),
    .B1_N(\u_cpu.REG_FILE._01214_ ),
    .X(\u_cpu.REG_FILE._01272_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05941_  (.A1(\u_cpu.REG_FILE._01151_ ),
    .A2(\u_cpu.REG_FILE.rf[21][2] ),
    .B1(\u_cpu.REG_FILE._01272_ ),
    .Y(\u_cpu.REG_FILE._01273_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._05942_  (.A(\u_cpu.REG_FILE._01271_ ),
    .B(\u_cpu.REG_FILE._01273_ ),
    .C(\u_cpu.REG_FILE._01156_ ),
    .Y(\u_cpu.REG_FILE._01274_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._05943_  (.A(\u_cpu.REG_FILE._01132_ ),
    .B(\u_cpu.REG_FILE._01268_ ),
    .C(\u_cpu.REG_FILE._01274_ ),
    .Y(\u_cpu.REG_FILE._01275_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._05944_  (.A(\u_cpu.REG_FILE._01257_ ),
    .B(\u_cpu.REG_FILE._01275_ ),
    .C(\u_cpu.REG_FILE._01159_ ),
    .Y(\u_cpu.REG_FILE._01276_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._05945_  (.A1(\u_cpu.REG_FILE._01026_ ),
    .A2(\u_cpu.REG_FILE._01246_ ),
    .B1(\u_cpu.REG_FILE._01276_ ),
    .C1(\u_cpu.REG_FILE._01165_ ),
    .X(\u_cpu.ALU.SrcA[2] ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05946_  (.A(\u_cpu.REG_FILE._01046_ ),
    .X(\u_cpu.REG_FILE._01277_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._05947_  (.A(\u_cpu.REG_FILE.rf[19][3] ),
    .Y(\u_cpu.REG_FILE._01278_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05948_  (.A(\u_cpu.REG_FILE._01076_ ),
    .X(\u_cpu.REG_FILE._01279_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05949_  (.A(\u_cpu.REG_FILE._01239_ ),
    .X(\u_cpu.REG_FILE._01280_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05950_  (.A1(\u_cpu.REG_FILE._01279_ ),
    .A2(\u_cpu.REG_FILE.rf[18][3] ),
    .B1(\u_cpu.REG_FILE._01280_ ),
    .Y(\u_cpu.REG_FILE._01281_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._05951_  (.A1(\u_cpu.REG_FILE._01278_ ),
    .A2(\u_cpu.REG_FILE._01075_ ),
    .B1(\u_cpu.REG_FILE._01281_ ),
    .Y(\u_cpu.REG_FILE._01282_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._05952_  (.A(\u_cpu.REG_FILE.rf[17][3] ),
    .Y(\u_cpu.REG_FILE._01283_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05953_  (.A(\u_cpu.REG_FILE._01161_ ),
    .X(\u_cpu.REG_FILE._01284_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._05954_  (.A(\u_cpu.REG_FILE._01061_ ),
    .B(\u_cpu.REG_FILE.rf[16][3] ),
    .Y(\u_cpu.REG_FILE._01285_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._05955_  (.A1(\u_cpu.REG_FILE._01283_ ),
    .A2(\u_cpu.REG_FILE._01284_ ),
    .B1(\u_cpu.REG_FILE._01259_ ),
    .C1(\u_cpu.REG_FILE._01285_ ),
    .Y(\u_cpu.REG_FILE._01286_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05956_  (.A(\u_cpu.REG_FILE._01038_ ),
    .X(\u_cpu.REG_FILE._01287_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05957_  (.A(\u_cpu.REG_FILE._01032_ ),
    .X(\u_cpu.REG_FILE._01288_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._05958_  (.A(\u_cpu.REG_FILE._01108_ ),
    .B(\u_cpu.REG_FILE.rf[22][3] ),
    .X(\u_cpu.REG_FILE._01289_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05959_  (.A1(\u_cpu.REG_FILE._01287_ ),
    .A2(\u_cpu.REG_FILE.rf[23][3] ),
    .B1(\u_cpu.REG_FILE._01288_ ),
    .C1(\u_cpu.REG_FILE._01289_ ),
    .Y(\u_cpu.REG_FILE._01290_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._05960_  (.A1(\u_cpu.REG_FILE._01111_ ),
    .A2(\u_cpu.REG_FILE.rf[20][3] ),
    .B1_N(\u_cpu.REG_FILE._01106_ ),
    .X(\u_cpu.REG_FILE._01291_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05961_  (.A1(\u_cpu.REG_FILE._01287_ ),
    .A2(\u_cpu.REG_FILE.rf[21][3] ),
    .B1(\u_cpu.REG_FILE._01291_ ),
    .Y(\u_cpu.REG_FILE._01292_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05962_  (.A(\u_cpu.REG_FILE._01046_ ),
    .X(\u_cpu.REG_FILE._01293_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._05963_  (.A(\u_cpu.REG_FILE._01290_ ),
    .B(\u_cpu.REG_FILE._01292_ ),
    .C(\u_cpu.REG_FILE._01293_ ),
    .Y(\u_cpu.REG_FILE._01294_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.REG_FILE._05964_  (.A1(\u_cpu.REG_FILE._01277_ ),
    .A2(\u_cpu.REG_FILE._01282_ ),
    .A3(\u_cpu.REG_FILE._01286_ ),
    .B1(\u_cpu.REG_FILE._01294_ ),
    .C1(\u_cpu.REG_FILE._01132_ ),
    .X(\u_cpu.REG_FILE._01295_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._05965_  (.A(\u_cpu.REG_FILE.rf[31][3] ),
    .B_N(\u_cpu.REG_FILE._01111_ ),
    .X(\u_cpu.REG_FILE._01296_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05966_  (.A1(\u_cpu.REG_FILE._01030_ ),
    .A2(\u_cpu.REG_FILE.rf[30][3] ),
    .B1(\u_cpu.REG_FILE._01033_ ),
    .C1(\u_cpu.REG_FILE._01296_ ),
    .Y(\u_cpu.REG_FILE._01297_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05967_  (.A(\u_cpu.REG_FILE._01038_ ),
    .X(\u_cpu.REG_FILE._01298_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05968_  (.A(\u_cpu.REG_FILE._01028_ ),
    .X(\u_cpu.REG_FILE._01299_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._05969_  (.A1(\u_cpu.REG_FILE._01299_ ),
    .A2(\u_cpu.REG_FILE.rf[28][3] ),
    .B1_N(\u_cpu.REG_FILE._01106_ ),
    .X(\u_cpu.REG_FILE._01300_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05970_  (.A1(\u_cpu.REG_FILE._01298_ ),
    .A2(\u_cpu.REG_FILE.rf[29][3] ),
    .B1(\u_cpu.REG_FILE._01300_ ),
    .Y(\u_cpu.REG_FILE._01301_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._05971_  (.A(\u_cpu.REG_FILE._01297_ ),
    .B(\u_cpu.REG_FILE._01301_ ),
    .C(\u_cpu.REG_FILE._01293_ ),
    .Y(\u_cpu.REG_FILE._01302_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._05972_  (.A_N(\u_cpu.REG_FILE.rf[25][3] ),
    .B(\u_cpu.REG_FILE._01074_ ),
    .X(\u_cpu.REG_FILE._01303_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05973_  (.A(\u_cpu.M_AXI_WDATA[16] ),
    .X(\u_cpu.REG_FILE._01304_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05974_  (.A(\u_cpu.REG_FILE._01304_ ),
    .X(\u_cpu.REG_FILE._01305_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._05975_  (.A1(\u_cpu.REG_FILE._01093_ ),
    .A2(\u_cpu.REG_FILE.rf[24][3] ),
    .B1_N(\u_cpu.REG_FILE._01305_ ),
    .Y(\u_cpu.REG_FILE._01306_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05976_  (.A(\u_cpu.REG_FILE._01058_ ),
    .X(\u_cpu.REG_FILE._01307_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05977_  (.A(\u_cpu.REG_FILE._01060_ ),
    .X(\u_cpu.REG_FILE._01308_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05978_  (.A(\u_cpu.REG_FILE._01112_ ),
    .X(\u_cpu.REG_FILE._01309_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05979_  (.A(\u_cpu.REG_FILE._01040_ ),
    .X(\u_cpu.REG_FILE._01310_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._05980_  (.A(\u_cpu.REG_FILE.rf[27][3] ),
    .B_N(\u_cpu.REG_FILE._01310_ ),
    .X(\u_cpu.REG_FILE._01311_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05981_  (.A1(\u_cpu.REG_FILE._01308_ ),
    .A2(\u_cpu.REG_FILE.rf[26][3] ),
    .B1(\u_cpu.REG_FILE._01309_ ),
    .C1(\u_cpu.REG_FILE._01311_ ),
    .Y(\u_cpu.REG_FILE._01312_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._05982_  (.A1(\u_cpu.REG_FILE._01303_ ),
    .A2(\u_cpu.REG_FILE._01306_ ),
    .B1(\u_cpu.REG_FILE._01307_ ),
    .C1(\u_cpu.REG_FILE._01312_ ),
    .Y(\u_cpu.REG_FILE._01313_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05983_  (.A(\u_cpu.M_AXI_WDATA[18] ),
    .X(\u_cpu.REG_FILE._01314_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._05984_  (.A(\u_cpu.REG_FILE._01024_ ),
    .Y(\u_cpu.REG_FILE._01315_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._05985_  (.A1(\u_cpu.REG_FILE._01302_ ),
    .A2(\u_cpu.REG_FILE._01313_ ),
    .A3(\u_cpu.REG_FILE._01314_ ),
    .B1(\u_cpu.REG_FILE._01315_ ),
    .X(\u_cpu.REG_FILE._01316_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05986_  (.A(\u_cpu.REG_FILE._01049_ ),
    .X(\u_cpu.REG_FILE._01317_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._05987_  (.A1(\u_cpu.REG_FILE._01317_ ),
    .A2(\u_cpu.REG_FILE.rf[8][3] ),
    .B1_N(\u_cpu.REG_FILE._01032_ ),
    .Y(\u_cpu.REG_FILE._01318_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._05988_  (.A_N(\u_cpu.REG_FILE.rf[9][3] ),
    .B(\u_cpu.REG_FILE._01041_ ),
    .X(\u_cpu.REG_FILE._01319_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05989_  (.A1(\u_cpu.REG_FILE._01318_ ),
    .A2(\u_cpu.REG_FILE._01319_ ),
    .B1(\u_cpu.REG_FILE._01264_ ),
    .Y(\u_cpu.REG_FILE._01320_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05990_  (.A(\u_cpu.REG_FILE._01037_ ),
    .X(\u_cpu.REG_FILE._01321_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._05991_  (.A(\u_cpu.REG_FILE._01148_ ),
    .B(\u_cpu.REG_FILE.rf[10][3] ),
    .X(\u_cpu.REG_FILE._01322_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._05992_  (.A1(\u_cpu.REG_FILE._01321_ ),
    .A2(\u_cpu.REG_FILE.rf[11][3] ),
    .B1(\u_cpu.REG_FILE._01280_ ),
    .C1(\u_cpu.REG_FILE._01322_ ),
    .X(\u_cpu.REG_FILE._01323_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05993_  (.A(\u_cpu.REG_FILE._01040_ ),
    .X(\u_cpu.REG_FILE._01324_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05994_  (.A(\u_cpu.REG_FILE._01324_ ),
    .X(\u_cpu.REG_FILE._01325_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._05995_  (.A(\u_cpu.REG_FILE._01325_ ),
    .B(\u_cpu.REG_FILE.rf[14][3] ),
    .Y(\u_cpu.REG_FILE._01326_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05996_  (.A(\u_cpu.REG_FILE._01037_ ),
    .X(\u_cpu.REG_FILE._01327_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._05997_  (.A1(\u_cpu.REG_FILE.rf[15][3] ),
    .A2(\u_cpu.REG_FILE._01327_ ),
    .B1(\u_cpu.REG_FILE._01099_ ),
    .Y(\u_cpu.REG_FILE._01328_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05998_  (.A(\u_cpu.REG_FILE._01037_ ),
    .X(\u_cpu.REG_FILE._01329_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._05999_  (.A(\u_cpu.REG_FILE._01064_ ),
    .X(\u_cpu.REG_FILE._01330_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06000_  (.A1(\u_cpu.REG_FILE._01330_ ),
    .A2(\u_cpu.REG_FILE.rf[12][3] ),
    .B1_N(\u_cpu.REG_FILE._01082_ ),
    .X(\u_cpu.REG_FILE._01331_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06001_  (.A1(\u_cpu.REG_FILE._01329_ ),
    .A2(\u_cpu.REG_FILE.rf[13][3] ),
    .B1(\u_cpu.REG_FILE._01331_ ),
    .Y(\u_cpu.REG_FILE._01332_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06002_  (.A(\u_cpu.REG_FILE._01046_ ),
    .X(\u_cpu.REG_FILE._01333_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06003_  (.A1(\u_cpu.REG_FILE._01326_ ),
    .A2(\u_cpu.REG_FILE._01328_ ),
    .B1(\u_cpu.REG_FILE._01332_ ),
    .C1(\u_cpu.REG_FILE._01333_ ),
    .Y(\u_cpu.REG_FILE._01334_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06004_  (.A1(\u_cpu.REG_FILE._01320_ ),
    .A2(\u_cpu.REG_FILE._01323_ ),
    .B1(\u_cpu.REG_FILE._01069_ ),
    .C1(\u_cpu.REG_FILE._01334_ ),
    .Y(\u_cpu.REG_FILE._01335_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06005_  (.A1(\u_cpu.REG_FILE._01317_ ),
    .A2(\u_cpu.REG_FILE.rf[0][3] ),
    .B1_N(\u_cpu.REG_FILE._01258_ ),
    .Y(\u_cpu.REG_FILE._01336_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06006_  (.A_N(\u_cpu.REG_FILE.rf[1][3] ),
    .B(\u_cpu.REG_FILE._01041_ ),
    .X(\u_cpu.REG_FILE._01337_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06007_  (.A1(\u_cpu.REG_FILE._01336_ ),
    .A2(\u_cpu.REG_FILE._01337_ ),
    .B1(\u_cpu.REG_FILE._01264_ ),
    .Y(\u_cpu.REG_FILE._01338_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06008_  (.A(\u_cpu.REG_FILE._01062_ ),
    .X(\u_cpu.REG_FILE._01339_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06009_  (.A(\u_cpu.REG_FILE._01040_ ),
    .X(\u_cpu.REG_FILE._01340_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06010_  (.A(\u_cpu.REG_FILE.rf[3][3] ),
    .B_N(\u_cpu.REG_FILE._01340_ ),
    .X(\u_cpu.REG_FILE._01341_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06011_  (.A1(\u_cpu.REG_FILE._01061_ ),
    .A2(\u_cpu.REG_FILE.rf[2][3] ),
    .B1(\u_cpu.REG_FILE._01339_ ),
    .C1(\u_cpu.REG_FILE._01341_ ),
    .X(\u_cpu.REG_FILE._01342_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06012_  (.A(\u_cpu.REG_FILE._01325_ ),
    .B(\u_cpu.REG_FILE.rf[6][3] ),
    .Y(\u_cpu.REG_FILE._01343_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06013_  (.A1(\u_cpu.REG_FILE.rf[7][3] ),
    .A2(\u_cpu.REG_FILE._01329_ ),
    .B1(\u_cpu.REG_FILE._01280_ ),
    .Y(\u_cpu.REG_FILE._01344_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06014_  (.A(\u_cpu.REG_FILE._01064_ ),
    .X(\u_cpu.REG_FILE._01345_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06015_  (.A1(\u_cpu.REG_FILE._01345_ ),
    .A2(\u_cpu.REG_FILE.rf[4][3] ),
    .B1_N(\u_cpu.REG_FILE._01134_ ),
    .X(\u_cpu.REG_FILE._01346_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06016_  (.A1(\u_cpu.REG_FILE._01265_ ),
    .A2(\u_cpu.REG_FILE.rf[5][3] ),
    .B1(\u_cpu.REG_FILE._01346_ ),
    .Y(\u_cpu.REG_FILE._01347_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06017_  (.A1(\u_cpu.REG_FILE._01343_ ),
    .A2(\u_cpu.REG_FILE._01344_ ),
    .B1(\u_cpu.REG_FILE._01347_ ),
    .C1(\u_cpu.REG_FILE._01333_ ),
    .Y(\u_cpu.REG_FILE._01348_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06018_  (.A1(\u_cpu.REG_FILE._01338_ ),
    .A2(\u_cpu.REG_FILE._01342_ ),
    .B1(\u_cpu.REG_FILE._01090_ ),
    .C1(\u_cpu.REG_FILE._01348_ ),
    .Y(\u_cpu.REG_FILE._01349_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06019_  (.A(\u_cpu.REG_FILE._01315_ ),
    .B(\u_cpu.REG_FILE._01335_ ),
    .C(\u_cpu.REG_FILE._01349_ ),
    .Y(\u_cpu.REG_FILE._01350_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06020_  (.A1(\u_cpu.REG_FILE._01295_ ),
    .A2(\u_cpu.REG_FILE._01316_ ),
    .B1(\u_cpu.REG_FILE._01350_ ),
    .C1(\u_cpu.REG_FILE._01165_ ),
    .X(\u_cpu.ALU.SrcA[3] ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06021_  (.A(\u_cpu.REG_FILE._01029_ ),
    .X(\u_cpu.REG_FILE._01351_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06022_  (.A(\u_cpu.REG_FILE._01258_ ),
    .X(\u_cpu.REG_FILE._01352_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06023_  (.A(\u_cpu.REG_FILE.rf[15][4] ),
    .B_N(\u_cpu.REG_FILE._01034_ ),
    .X(\u_cpu.REG_FILE._01353_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06024_  (.A1(\u_cpu.REG_FILE._01351_ ),
    .A2(\u_cpu.REG_FILE.rf[14][4] ),
    .B1(\u_cpu.REG_FILE._01352_ ),
    .C1(\u_cpu.REG_FILE._01353_ ),
    .Y(\u_cpu.REG_FILE._01354_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06025_  (.A1(\u_cpu.REG_FILE._01041_ ),
    .A2(\u_cpu.REG_FILE.rf[12][4] ),
    .B1_N(\u_cpu.REG_FILE._01042_ ),
    .X(\u_cpu.REG_FILE._01355_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06026_  (.A1(\u_cpu.REG_FILE._01039_ ),
    .A2(\u_cpu.REG_FILE.rf[13][4] ),
    .B1(\u_cpu.REG_FILE._01355_ ),
    .Y(\u_cpu.REG_FILE._01356_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06027_  (.A(\u_cpu.REG_FILE._01354_ ),
    .B(\u_cpu.REG_FILE._01356_ ),
    .C(\u_cpu.REG_FILE._01047_ ),
    .Y(\u_cpu.REG_FILE._01357_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06028_  (.A_N(\u_cpu.REG_FILE.rf[9][4] ),
    .B(\u_cpu.REG_FILE._01050_ ),
    .X(\u_cpu.REG_FILE._01358_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06029_  (.A1(\u_cpu.REG_FILE._01053_ ),
    .A2(\u_cpu.REG_FILE.rf[8][4] ),
    .B1_N(\u_cpu.REG_FILE._01055_ ),
    .Y(\u_cpu.REG_FILE._01359_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06030_  (.A(\u_cpu.REG_FILE._01062_ ),
    .X(\u_cpu.REG_FILE._01360_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06031_  (.A(\u_cpu.REG_FILE.rf[11][4] ),
    .B_N(\u_cpu.REG_FILE._01065_ ),
    .X(\u_cpu.REG_FILE._01361_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06032_  (.A1(\u_cpu.REG_FILE._01061_ ),
    .A2(\u_cpu.REG_FILE.rf[10][4] ),
    .B1(\u_cpu.REG_FILE._01360_ ),
    .C1(\u_cpu.REG_FILE._01361_ ),
    .Y(\u_cpu.REG_FILE._01362_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06033_  (.A1(\u_cpu.REG_FILE._01358_ ),
    .A2(\u_cpu.REG_FILE._01359_ ),
    .B1(\u_cpu.REG_FILE._01059_ ),
    .C1(\u_cpu.REG_FILE._01362_ ),
    .Y(\u_cpu.REG_FILE._01363_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06034_  (.A(\u_cpu.REG_FILE._01357_ ),
    .B(\u_cpu.REG_FILE._01363_ ),
    .C(\u_cpu.REG_FILE._01070_ ),
    .Y(\u_cpu.REG_FILE._01364_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06035_  (.A(\u_cpu.REG_FILE.rf[5][4] ),
    .Y(\u_cpu.REG_FILE._01365_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06036_  (.A1(\u_cpu.REG_FILE._01077_ ),
    .A2(\u_cpu.REG_FILE.rf[4][4] ),
    .B1_N(\u_cpu.REG_FILE._01078_ ),
    .Y(\u_cpu.REG_FILE._01366_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._06037_  (.A1(\u_cpu.REG_FILE._01365_ ),
    .A2(\u_cpu.REG_FILE._01075_ ),
    .B1(\u_cpu.REG_FILE._01366_ ),
    .Y(\u_cpu.REG_FILE._01367_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06038_  (.A1(\u_cpu.REG_FILE._01081_ ),
    .A2(\u_cpu.REG_FILE.rf[6][4] ),
    .B1(\u_cpu.REG_FILE._01083_ ),
    .Y(\u_cpu.REG_FILE._01368_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06039_  (.A_N(\u_cpu.REG_FILE.rf[7][4] ),
    .B(\u_cpu.REG_FILE._01085_ ),
    .X(\u_cpu.REG_FILE._01369_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06040_  (.A1(\u_cpu.REG_FILE._01368_ ),
    .A2(\u_cpu.REG_FILE._01369_ ),
    .B1(\u_cpu.REG_FILE._01087_ ),
    .Y(\u_cpu.REG_FILE._01370_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06041_  (.A_N(\u_cpu.REG_FILE.rf[1][4] ),
    .B(\u_cpu.REG_FILE._01091_ ),
    .X(\u_cpu.REG_FILE._01371_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06042_  (.A(\u_cpu.REG_FILE._01076_ ),
    .X(\u_cpu.REG_FILE._01372_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06043_  (.A1(\u_cpu.REG_FILE._01372_ ),
    .A2(\u_cpu.REG_FILE.rf[0][4] ),
    .B1_N(\u_cpu.REG_FILE._01094_ ),
    .Y(\u_cpu.REG_FILE._01373_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06044_  (.A(\u_cpu.REG_FILE.rf[3][4] ),
    .B_N(\u_cpu.REG_FILE._01241_ ),
    .X(\u_cpu.REG_FILE._01374_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06045_  (.A1(\u_cpu.REG_FILE._01097_ ),
    .A2(\u_cpu.REG_FILE.rf[2][4] ),
    .B1(\u_cpu.REG_FILE._01240_ ),
    .C1(\u_cpu.REG_FILE._01374_ ),
    .Y(\u_cpu.REG_FILE._01375_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06046_  (.A1(\u_cpu.REG_FILE._01371_ ),
    .A2(\u_cpu.REG_FILE._01373_ ),
    .B1(\u_cpu.REG_FILE._01096_ ),
    .C1(\u_cpu.REG_FILE._01375_ ),
    .Y(\u_cpu.REG_FILE._01376_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06047_  (.A1(\u_cpu.REG_FILE._01367_ ),
    .A2(\u_cpu.REG_FILE._01370_ ),
    .B1(\u_cpu.REG_FILE._01090_ ),
    .C1(\u_cpu.REG_FILE._01376_ ),
    .Y(\u_cpu.REG_FILE._01377_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._06048_  (.A(\u_cpu.REG_FILE._01364_ ),
    .B(\u_cpu.REG_FILE._01377_ ),
    .Y(\u_cpu.REG_FILE._01378_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06049_  (.A(\u_cpu.REG_FILE._01049_ ),
    .X(\u_cpu.REG_FILE._01379_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06050_  (.A(\u_cpu.REG_FILE._01054_ ),
    .X(\u_cpu.REG_FILE._01380_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06051_  (.A1(\u_cpu.REG_FILE._01379_ ),
    .A2(\u_cpu.REG_FILE.rf[24][4] ),
    .B1_N(\u_cpu.REG_FILE._01380_ ),
    .Y(\u_cpu.REG_FILE._01381_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06052_  (.A(\u_cpu.REG_FILE._01073_ ),
    .X(\u_cpu.REG_FILE._01382_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06053_  (.A_N(\u_cpu.REG_FILE.rf[25][4] ),
    .B(\u_cpu.REG_FILE._01382_ ),
    .X(\u_cpu.REG_FILE._01383_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06054_  (.A(\u_cpu.REG_FILE._01058_ ),
    .X(\u_cpu.REG_FILE._01384_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06055_  (.A1(\u_cpu.REG_FILE._01381_ ),
    .A2(\u_cpu.REG_FILE._01383_ ),
    .B1(\u_cpu.REG_FILE._01384_ ),
    .Y(\u_cpu.REG_FILE._01385_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06056_  (.A(\u_cpu.REG_FILE._01123_ ),
    .X(\u_cpu.REG_FILE._01386_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06057_  (.A(\u_cpu.REG_FILE._01032_ ),
    .X(\u_cpu.REG_FILE._01387_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06058_  (.A(\u_cpu.REG_FILE._01340_ ),
    .B(\u_cpu.REG_FILE.rf[26][4] ),
    .X(\u_cpu.REG_FILE._01388_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06059_  (.A1(\u_cpu.REG_FILE._01386_ ),
    .A2(\u_cpu.REG_FILE.rf[27][4] ),
    .B1(\u_cpu.REG_FILE._01387_ ),
    .C1(\u_cpu.REG_FILE._01388_ ),
    .X(\u_cpu.REG_FILE._01389_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06060_  (.A(\u_cpu.REG_FILE._01345_ ),
    .X(\u_cpu.REG_FILE._01390_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06061_  (.A(\u_cpu.REG_FILE._01390_ ),
    .B(\u_cpu.REG_FILE.rf[30][4] ),
    .Y(\u_cpu.REG_FILE._01391_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06062_  (.A1(\u_cpu.REG_FILE.rf[31][4] ),
    .A2(\u_cpu.REG_FILE._01200_ ),
    .B1(\u_cpu.REG_FILE._01121_ ),
    .Y(\u_cpu.REG_FILE._01392_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06063_  (.A1(\u_cpu.REG_FILE._01125_ ),
    .A2(\u_cpu.REG_FILE.rf[28][4] ),
    .B1_N(\u_cpu.REG_FILE._01126_ ),
    .X(\u_cpu.REG_FILE._01393_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06064_  (.A1(\u_cpu.REG_FILE._01124_ ),
    .A2(\u_cpu.REG_FILE.rf[29][4] ),
    .B1(\u_cpu.REG_FILE._01393_ ),
    .Y(\u_cpu.REG_FILE._01394_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06065_  (.A(\u_cpu.REG_FILE._01046_ ),
    .X(\u_cpu.REG_FILE._01395_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06066_  (.A1(\u_cpu.REG_FILE._01391_ ),
    .A2(\u_cpu.REG_FILE._01392_ ),
    .B1(\u_cpu.REG_FILE._01394_ ),
    .C1(\u_cpu.REG_FILE._01395_ ),
    .Y(\u_cpu.REG_FILE._01396_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06067_  (.A1(\u_cpu.REG_FILE._01385_ ),
    .A2(\u_cpu.REG_FILE._01389_ ),
    .B1(\u_cpu.REG_FILE._01198_ ),
    .C1(\u_cpu.REG_FILE._01396_ ),
    .Y(\u_cpu.REG_FILE._01397_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06068_  (.A(\u_cpu.REG_FILE.rf[19][4] ),
    .Y(\u_cpu.REG_FILE._01398_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06069_  (.A(\u_cpu.REG_FILE._01111_ ),
    .X(\u_cpu.REG_FILE._01399_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06070_  (.A(\u_cpu.REG_FILE._01304_ ),
    .X(\u_cpu.REG_FILE._01400_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06071_  (.A1(\u_cpu.REG_FILE._01317_ ),
    .A2(\u_cpu.REG_FILE.rf[18][4] ),
    .B1(\u_cpu.REG_FILE._01400_ ),
    .Y(\u_cpu.REG_FILE._01401_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._06072_  (.A1(\u_cpu.REG_FILE._01398_ ),
    .A2(\u_cpu.REG_FILE._01399_ ),
    .B1(\u_cpu.REG_FILE._01401_ ),
    .Y(\u_cpu.REG_FILE._01402_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06073_  (.A(\u_cpu.REG_FILE.rf[17][4] ),
    .Y(\u_cpu.REG_FILE._01403_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06074_  (.A(\u_cpu.REG_FILE._01049_ ),
    .X(\u_cpu.REG_FILE._01404_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06075_  (.A1(\u_cpu.REG_FILE._01404_ ),
    .A2(\u_cpu.REG_FILE.rf[16][4] ),
    .B1_N(\u_cpu.REG_FILE._01258_ ),
    .Y(\u_cpu.REG_FILE._01405_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._06076_  (.A1(\u_cpu.REG_FILE._01403_ ),
    .A2(\u_cpu.REG_FILE._01284_ ),
    .B1(\u_cpu.REG_FILE._01405_ ),
    .Y(\u_cpu.REG_FILE._01406_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06077_  (.A(\u_cpu.REG_FILE._01082_ ),
    .X(\u_cpu.REG_FILE._01407_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06078_  (.A(\u_cpu.REG_FILE._01027_ ),
    .X(\u_cpu.REG_FILE._01408_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06079_  (.A(\u_cpu.REG_FILE.rf[23][4] ),
    .B_N(\u_cpu.REG_FILE._01408_ ),
    .X(\u_cpu.REG_FILE._01409_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06080_  (.A1(\u_cpu.REG_FILE._01077_ ),
    .A2(\u_cpu.REG_FILE.rf[22][4] ),
    .B1(\u_cpu.REG_FILE._01407_ ),
    .C1(\u_cpu.REG_FILE._01409_ ),
    .Y(\u_cpu.REG_FILE._01410_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06081_  (.A1(\u_cpu.REG_FILE._01324_ ),
    .A2(\u_cpu.REG_FILE.rf[20][4] ),
    .B1_N(\u_cpu.REG_FILE._01304_ ),
    .X(\u_cpu.REG_FILE._01411_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06082_  (.A1(\u_cpu.REG_FILE._01038_ ),
    .A2(\u_cpu.REG_FILE.rf[21][4] ),
    .B1(\u_cpu.REG_FILE._01411_ ),
    .Y(\u_cpu.REG_FILE._01412_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06083_  (.A(\u_cpu.REG_FILE._01410_ ),
    .B(\u_cpu.REG_FILE._01412_ ),
    .C(\u_cpu.REG_FILE._01115_ ),
    .Y(\u_cpu.REG_FILE._01413_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06084_  (.A(\u_cpu.REG_FILE._01089_ ),
    .X(\u_cpu.REG_FILE._01414_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._06085_  (.A1(\u_cpu.REG_FILE._01277_ ),
    .A2(\u_cpu.REG_FILE._01402_ ),
    .A3(\u_cpu.REG_FILE._01406_ ),
    .B1(\u_cpu.REG_FILE._01413_ ),
    .C1(\u_cpu.REG_FILE._01414_ ),
    .Y(\u_cpu.REG_FILE._01415_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06086_  (.A(\u_cpu.REG_FILE._01397_ ),
    .B(\u_cpu.REG_FILE._01415_ ),
    .C(\u_cpu.REG_FILE._01159_ ),
    .Y(\u_cpu.REG_FILE._01416_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06087_  (.A1(\u_cpu.REG_FILE._01026_ ),
    .A2(\u_cpu.REG_FILE._01378_ ),
    .B1(\u_cpu.REG_FILE._01416_ ),
    .C1(\u_cpu.REG_FILE._01165_ ),
    .X(\u_cpu.ALU.SrcA[4] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06088_  (.A(\u_cpu.REG_FILE.rf[15][5] ),
    .B_N(\u_cpu.REG_FILE._01034_ ),
    .X(\u_cpu.REG_FILE._01417_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06089_  (.A1(\u_cpu.REG_FILE._01351_ ),
    .A2(\u_cpu.REG_FILE.rf[14][5] ),
    .B1(\u_cpu.REG_FILE._01352_ ),
    .C1(\u_cpu.REG_FILE._01417_ ),
    .Y(\u_cpu.REG_FILE._01418_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06090_  (.A1(\u_cpu.REG_FILE._01041_ ),
    .A2(\u_cpu.REG_FILE.rf[12][5] ),
    .B1_N(\u_cpu.REG_FILE._01042_ ),
    .X(\u_cpu.REG_FILE._01419_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06091_  (.A1(\u_cpu.REG_FILE._01039_ ),
    .A2(\u_cpu.REG_FILE.rf[13][5] ),
    .B1(\u_cpu.REG_FILE._01419_ ),
    .Y(\u_cpu.REG_FILE._01420_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06092_  (.A(\u_cpu.REG_FILE._01418_ ),
    .B(\u_cpu.REG_FILE._01420_ ),
    .C(\u_cpu.REG_FILE._01047_ ),
    .Y(\u_cpu.REG_FILE._01421_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06093_  (.A_N(\u_cpu.REG_FILE.rf[9][5] ),
    .B(\u_cpu.REG_FILE._01050_ ),
    .X(\u_cpu.REG_FILE._01422_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06094_  (.A1(\u_cpu.REG_FILE._01053_ ),
    .A2(\u_cpu.REG_FILE.rf[8][5] ),
    .B1_N(\u_cpu.REG_FILE._01055_ ),
    .Y(\u_cpu.REG_FILE._01423_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06095_  (.A(\u_cpu.REG_FILE._01058_ ),
    .X(\u_cpu.REG_FILE._01424_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06096_  (.A(\u_cpu.REG_FILE._01060_ ),
    .X(\u_cpu.REG_FILE._01425_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06097_  (.A(\u_cpu.REG_FILE.rf[11][5] ),
    .B_N(\u_cpu.REG_FILE._01065_ ),
    .X(\u_cpu.REG_FILE._01426_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06098_  (.A1(\u_cpu.REG_FILE._01425_ ),
    .A2(\u_cpu.REG_FILE.rf[10][5] ),
    .B1(\u_cpu.REG_FILE._01360_ ),
    .C1(\u_cpu.REG_FILE._01426_ ),
    .Y(\u_cpu.REG_FILE._01427_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06099_  (.A1(\u_cpu.REG_FILE._01422_ ),
    .A2(\u_cpu.REG_FILE._01423_ ),
    .B1(\u_cpu.REG_FILE._01424_ ),
    .C1(\u_cpu.REG_FILE._01427_ ),
    .Y(\u_cpu.REG_FILE._01428_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06100_  (.A(\u_cpu.REG_FILE._01421_ ),
    .B(\u_cpu.REG_FILE._01428_ ),
    .C(\u_cpu.REG_FILE._01070_ ),
    .Y(\u_cpu.REG_FILE._01429_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06101_  (.A(\u_cpu.REG_FILE.rf[5][5] ),
    .Y(\u_cpu.REG_FILE._01430_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06102_  (.A(\u_cpu.REG_FILE._01076_ ),
    .X(\u_cpu.REG_FILE._01431_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06103_  (.A1(\u_cpu.REG_FILE._01431_ ),
    .A2(\u_cpu.REG_FILE.rf[4][5] ),
    .B1_N(\u_cpu.REG_FILE._01078_ ),
    .Y(\u_cpu.REG_FILE._01432_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._06104_  (.A1(\u_cpu.REG_FILE._01430_ ),
    .A2(\u_cpu.REG_FILE._01075_ ),
    .B1(\u_cpu.REG_FILE._01432_ ),
    .Y(\u_cpu.REG_FILE._01433_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06105_  (.A(\u_cpu.REG_FILE._01049_ ),
    .X(\u_cpu.REG_FILE._01434_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06106_  (.A1(\u_cpu.REG_FILE._01434_ ),
    .A2(\u_cpu.REG_FILE.rf[6][5] ),
    .B1(\u_cpu.REG_FILE._01083_ ),
    .Y(\u_cpu.REG_FILE._01435_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06107_  (.A_N(\u_cpu.REG_FILE.rf[7][5] ),
    .B(\u_cpu.REG_FILE._01085_ ),
    .X(\u_cpu.REG_FILE._01436_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06108_  (.A1(\u_cpu.REG_FILE._01435_ ),
    .A2(\u_cpu.REG_FILE._01436_ ),
    .B1(\u_cpu.REG_FILE._01087_ ),
    .Y(\u_cpu.REG_FILE._01437_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06109_  (.A_N(\u_cpu.REG_FILE.rf[1][5] ),
    .B(\u_cpu.REG_FILE._01091_ ),
    .X(\u_cpu.REG_FILE._01438_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06110_  (.A1(\u_cpu.REG_FILE._01372_ ),
    .A2(\u_cpu.REG_FILE.rf[0][5] ),
    .B1_N(\u_cpu.REG_FILE._01094_ ),
    .Y(\u_cpu.REG_FILE._01439_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06111_  (.A(\u_cpu.REG_FILE.rf[3][5] ),
    .B_N(\u_cpu.REG_FILE._01241_ ),
    .X(\u_cpu.REG_FILE._01440_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06112_  (.A1(\u_cpu.REG_FILE._01097_ ),
    .A2(\u_cpu.REG_FILE.rf[2][5] ),
    .B1(\u_cpu.REG_FILE._01240_ ),
    .C1(\u_cpu.REG_FILE._01440_ ),
    .Y(\u_cpu.REG_FILE._01441_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06113_  (.A1(\u_cpu.REG_FILE._01438_ ),
    .A2(\u_cpu.REG_FILE._01439_ ),
    .B1(\u_cpu.REG_FILE._01096_ ),
    .C1(\u_cpu.REG_FILE._01441_ ),
    .Y(\u_cpu.REG_FILE._01442_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06114_  (.A1(\u_cpu.REG_FILE._01433_ ),
    .A2(\u_cpu.REG_FILE._01437_ ),
    .B1(\u_cpu.REG_FILE._01090_ ),
    .C1(\u_cpu.REG_FILE._01442_ ),
    .Y(\u_cpu.REG_FILE._01443_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._06115_  (.A(\u_cpu.REG_FILE._01429_ ),
    .B(\u_cpu.REG_FILE._01443_ ),
    .Y(\u_cpu.REG_FILE._01444_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06116_  (.A(\u_cpu.REG_FILE.rf[27][5] ),
    .B_N(\u_cpu.REG_FILE._01108_ ),
    .X(\u_cpu.REG_FILE._01445_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06117_  (.A1(\u_cpu.REG_FILE._01105_ ),
    .A2(\u_cpu.REG_FILE.rf[26][5] ),
    .B1(\u_cpu.REG_FILE._01107_ ),
    .C1(\u_cpu.REG_FILE._01445_ ),
    .X(\u_cpu.REG_FILE._01446_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06118_  (.A(\u_cpu.REG_FILE._01028_ ),
    .X(\u_cpu.REG_FILE._01447_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06119_  (.A1(\u_cpu.REG_FILE._01447_ ),
    .A2(\u_cpu.REG_FILE.rf[24][5] ),
    .B1_N(\u_cpu.REG_FILE._01112_ ),
    .X(\u_cpu.REG_FILE._01448_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06120_  (.A(\u_cpu.REG_FILE.rf[25][5] ),
    .B_N(\u_cpu.REG_FILE._01194_ ),
    .X(\u_cpu.REG_FILE._01449_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._06121_  (.A1(\u_cpu.REG_FILE._01448_ ),
    .A2(\u_cpu.REG_FILE._01449_ ),
    .B1(\u_cpu.REG_FILE._01196_ ),
    .X(\u_cpu.REG_FILE._01450_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06122_  (.A(\u_cpu.REG_FILE._01390_ ),
    .B(\u_cpu.REG_FILE.rf[30][5] ),
    .Y(\u_cpu.REG_FILE._01451_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06123_  (.A1(\u_cpu.REG_FILE.rf[31][5] ),
    .A2(\u_cpu.REG_FILE._01200_ ),
    .B1(\u_cpu.REG_FILE._01121_ ),
    .Y(\u_cpu.REG_FILE._01452_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06124_  (.A1(\u_cpu.REG_FILE._01125_ ),
    .A2(\u_cpu.REG_FILE.rf[28][5] ),
    .B1_N(\u_cpu.REG_FILE._01126_ ),
    .X(\u_cpu.REG_FILE._01453_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06125_  (.A1(\u_cpu.REG_FILE._01124_ ),
    .A2(\u_cpu.REG_FILE.rf[29][5] ),
    .B1(\u_cpu.REG_FILE._01453_ ),
    .Y(\u_cpu.REG_FILE._01454_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06126_  (.A1(\u_cpu.REG_FILE._01451_ ),
    .A2(\u_cpu.REG_FILE._01452_ ),
    .B1(\u_cpu.REG_FILE._01454_ ),
    .C1(\u_cpu.REG_FILE._01395_ ),
    .Y(\u_cpu.REG_FILE._01455_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06127_  (.A1(\u_cpu.REG_FILE._01446_ ),
    .A2(\u_cpu.REG_FILE._01450_ ),
    .B1(\u_cpu.REG_FILE._01198_ ),
    .C1(\u_cpu.REG_FILE._01455_ ),
    .Y(\u_cpu.REG_FILE._01456_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06128_  (.A(\u_cpu.REG_FILE._01379_ ),
    .B(\u_cpu.REG_FILE.rf[16][5] ),
    .Y(\u_cpu.REG_FILE._01457_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06129_  (.A_N(\u_cpu.REG_FILE.rf[17][5] ),
    .B(\u_cpu.REG_FILE._01262_ ),
    .X(\u_cpu.REG_FILE._01458_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.REG_FILE._06130_  (.A1(\u_cpu.REG_FILE._01060_ ),
    .A2(\u_cpu.REG_FILE.rf[18][5] ),
    .B1(\u_cpu.REG_FILE._01239_ ),
    .X(\u_cpu.REG_FILE._01459_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06131_  (.A1(\u_cpu.REG_FILE.rf[19][5] ),
    .A2(\u_cpu.REG_FILE._01265_ ),
    .B1(\u_cpu.REG_FILE._01459_ ),
    .Y(\u_cpu.REG_FILE._01460_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._06132_  (.A1(\u_cpu.REG_FILE._01033_ ),
    .A2(\u_cpu.REG_FILE._01457_ ),
    .A3(\u_cpu.REG_FILE._01458_ ),
    .B1(\u_cpu.REG_FILE._01058_ ),
    .C1(\u_cpu.REG_FILE._01460_ ),
    .Y(\u_cpu.REG_FILE._01461_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06133_  (.A(\u_cpu.REG_FILE._01269_ ),
    .B(\u_cpu.REG_FILE.rf[22][5] ),
    .X(\u_cpu.REG_FILE._01462_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06134_  (.A1(\u_cpu.REG_FILE._01146_ ),
    .A2(\u_cpu.REG_FILE.rf[23][5] ),
    .B1(\u_cpu.REG_FILE._01147_ ),
    .C1(\u_cpu.REG_FILE._01462_ ),
    .Y(\u_cpu.REG_FILE._01463_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06135_  (.A1(\u_cpu.REG_FILE._01152_ ),
    .A2(\u_cpu.REG_FILE.rf[20][5] ),
    .B1_N(\u_cpu.REG_FILE._01214_ ),
    .X(\u_cpu.REG_FILE._01464_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06136_  (.A1(\u_cpu.REG_FILE._01151_ ),
    .A2(\u_cpu.REG_FILE.rf[21][5] ),
    .B1(\u_cpu.REG_FILE._01464_ ),
    .Y(\u_cpu.REG_FILE._01465_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06137_  (.A(\u_cpu.REG_FILE._01463_ ),
    .B(\u_cpu.REG_FILE._01465_ ),
    .C(\u_cpu.REG_FILE._01156_ ),
    .Y(\u_cpu.REG_FILE._01466_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06138_  (.A(\u_cpu.REG_FILE._01132_ ),
    .B(\u_cpu.REG_FILE._01461_ ),
    .C(\u_cpu.REG_FILE._01466_ ),
    .Y(\u_cpu.REG_FILE._01467_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06139_  (.A(\u_cpu.REG_FILE._01456_ ),
    .B(\u_cpu.REG_FILE._01467_ ),
    .C(\u_cpu.REG_FILE._01159_ ),
    .Y(\u_cpu.REG_FILE._01468_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06140_  (.A1(\u_cpu.REG_FILE._01026_ ),
    .A2(\u_cpu.REG_FILE._01444_ ),
    .B1(\u_cpu.REG_FILE._01468_ ),
    .C1(\u_cpu.REG_FILE._01165_ ),
    .X(\u_cpu.ALU.SrcA[5] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06141_  (.A(\u_cpu.REG_FILE.rf[15][6] ),
    .B_N(\u_cpu.REG_FILE._01034_ ),
    .X(\u_cpu.REG_FILE._01469_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06142_  (.A1(\u_cpu.REG_FILE._01351_ ),
    .A2(\u_cpu.REG_FILE.rf[14][6] ),
    .B1(\u_cpu.REG_FILE._01352_ ),
    .C1(\u_cpu.REG_FILE._01469_ ),
    .Y(\u_cpu.REG_FILE._01470_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06143_  (.A1(\u_cpu.REG_FILE._01041_ ),
    .A2(\u_cpu.REG_FILE.rf[12][6] ),
    .B1_N(\u_cpu.REG_FILE._01042_ ),
    .X(\u_cpu.REG_FILE._01471_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06144_  (.A1(\u_cpu.REG_FILE._01039_ ),
    .A2(\u_cpu.REG_FILE.rf[13][6] ),
    .B1(\u_cpu.REG_FILE._01471_ ),
    .Y(\u_cpu.REG_FILE._01472_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06145_  (.A(\u_cpu.REG_FILE._01470_ ),
    .B(\u_cpu.REG_FILE._01472_ ),
    .C(\u_cpu.REG_FILE._01047_ ),
    .Y(\u_cpu.REG_FILE._01473_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06146_  (.A_N(\u_cpu.REG_FILE.rf[9][6] ),
    .B(\u_cpu.REG_FILE._01050_ ),
    .X(\u_cpu.REG_FILE._01474_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06147_  (.A(\u_cpu.REG_FILE._01052_ ),
    .X(\u_cpu.REG_FILE._01475_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06148_  (.A1(\u_cpu.REG_FILE._01475_ ),
    .A2(\u_cpu.REG_FILE.rf[8][6] ),
    .B1_N(\u_cpu.REG_FILE._01055_ ),
    .Y(\u_cpu.REG_FILE._01476_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06149_  (.A(\u_cpu.REG_FILE.rf[11][6] ),
    .B_N(\u_cpu.REG_FILE._01065_ ),
    .X(\u_cpu.REG_FILE._01477_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06150_  (.A1(\u_cpu.REG_FILE._01425_ ),
    .A2(\u_cpu.REG_FILE.rf[10][6] ),
    .B1(\u_cpu.REG_FILE._01360_ ),
    .C1(\u_cpu.REG_FILE._01477_ ),
    .Y(\u_cpu.REG_FILE._01478_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06151_  (.A1(\u_cpu.REG_FILE._01474_ ),
    .A2(\u_cpu.REG_FILE._01476_ ),
    .B1(\u_cpu.REG_FILE._01424_ ),
    .C1(\u_cpu.REG_FILE._01478_ ),
    .Y(\u_cpu.REG_FILE._01479_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06152_  (.A(\u_cpu.REG_FILE._01473_ ),
    .B(\u_cpu.REG_FILE._01479_ ),
    .C(\u_cpu.REG_FILE._01070_ ),
    .Y(\u_cpu.REG_FILE._01480_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06153_  (.A(\u_cpu.REG_FILE.rf[5][6] ),
    .Y(\u_cpu.REG_FILE._01481_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06154_  (.A(\u_cpu.REG_FILE._01054_ ),
    .X(\u_cpu.REG_FILE._01482_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06155_  (.A1(\u_cpu.REG_FILE._01431_ ),
    .A2(\u_cpu.REG_FILE.rf[4][6] ),
    .B1_N(\u_cpu.REG_FILE._01482_ ),
    .Y(\u_cpu.REG_FILE._01483_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._06156_  (.A1(\u_cpu.REG_FILE._01481_ ),
    .A2(\u_cpu.REG_FILE._01075_ ),
    .B1(\u_cpu.REG_FILE._01483_ ),
    .Y(\u_cpu.REG_FILE._01484_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06157_  (.A1(\u_cpu.REG_FILE._01434_ ),
    .A2(\u_cpu.REG_FILE.rf[6][6] ),
    .B1(\u_cpu.REG_FILE._01083_ ),
    .Y(\u_cpu.REG_FILE._01485_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06158_  (.A_N(\u_cpu.REG_FILE.rf[7][6] ),
    .B(\u_cpu.REG_FILE._01085_ ),
    .X(\u_cpu.REG_FILE._01486_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06159_  (.A1(\u_cpu.REG_FILE._01485_ ),
    .A2(\u_cpu.REG_FILE._01486_ ),
    .B1(\u_cpu.REG_FILE._01087_ ),
    .Y(\u_cpu.REG_FILE._01487_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06160_  (.A_N(\u_cpu.REG_FILE.rf[1][6] ),
    .B(\u_cpu.REG_FILE._01091_ ),
    .X(\u_cpu.REG_FILE._01488_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06161_  (.A1(\u_cpu.REG_FILE._01372_ ),
    .A2(\u_cpu.REG_FILE.rf[0][6] ),
    .B1_N(\u_cpu.REG_FILE._01094_ ),
    .Y(\u_cpu.REG_FILE._01489_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06162_  (.A(\u_cpu.REG_FILE.rf[3][6] ),
    .B_N(\u_cpu.REG_FILE._01241_ ),
    .X(\u_cpu.REG_FILE._01490_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06163_  (.A1(\u_cpu.REG_FILE._01097_ ),
    .A2(\u_cpu.REG_FILE.rf[2][6] ),
    .B1(\u_cpu.REG_FILE._01240_ ),
    .C1(\u_cpu.REG_FILE._01490_ ),
    .Y(\u_cpu.REG_FILE._01491_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06164_  (.A1(\u_cpu.REG_FILE._01488_ ),
    .A2(\u_cpu.REG_FILE._01489_ ),
    .B1(\u_cpu.REG_FILE._01096_ ),
    .C1(\u_cpu.REG_FILE._01491_ ),
    .Y(\u_cpu.REG_FILE._01492_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06165_  (.A1(\u_cpu.REG_FILE._01484_ ),
    .A2(\u_cpu.REG_FILE._01487_ ),
    .B1(\u_cpu.REG_FILE._01090_ ),
    .C1(\u_cpu.REG_FILE._01492_ ),
    .Y(\u_cpu.REG_FILE._01493_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._06166_  (.A(\u_cpu.REG_FILE._01480_ ),
    .B(\u_cpu.REG_FILE._01493_ ),
    .Y(\u_cpu.REG_FILE._01494_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06167_  (.A(\u_cpu.REG_FILE.rf[27][6] ),
    .B_N(\u_cpu.REG_FILE._01108_ ),
    .X(\u_cpu.REG_FILE._01495_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06168_  (.A1(\u_cpu.REG_FILE._01105_ ),
    .A2(\u_cpu.REG_FILE.rf[26][6] ),
    .B1(\u_cpu.REG_FILE._01107_ ),
    .C1(\u_cpu.REG_FILE._01495_ ),
    .X(\u_cpu.REG_FILE._01496_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06169_  (.A1(\u_cpu.REG_FILE._01447_ ),
    .A2(\u_cpu.REG_FILE.rf[24][6] ),
    .B1_N(\u_cpu.REG_FILE._01112_ ),
    .X(\u_cpu.REG_FILE._01497_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06170_  (.A(\u_cpu.REG_FILE.rf[25][6] ),
    .B_N(\u_cpu.REG_FILE._01194_ ),
    .X(\u_cpu.REG_FILE._01498_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._06171_  (.A1(\u_cpu.REG_FILE._01497_ ),
    .A2(\u_cpu.REG_FILE._01498_ ),
    .B1(\u_cpu.REG_FILE._01196_ ),
    .X(\u_cpu.REG_FILE._01499_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06172_  (.A(\u_cpu.REG_FILE._01390_ ),
    .B(\u_cpu.REG_FILE.rf[30][6] ),
    .Y(\u_cpu.REG_FILE._01500_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06173_  (.A(\u_cpu.REG_FILE._01112_ ),
    .X(\u_cpu.REG_FILE._01501_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06174_  (.A1(\u_cpu.REG_FILE.rf[31][6] ),
    .A2(\u_cpu.REG_FILE._01200_ ),
    .B1(\u_cpu.REG_FILE._01501_ ),
    .Y(\u_cpu.REG_FILE._01502_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06175_  (.A(\u_cpu.REG_FILE._01028_ ),
    .X(\u_cpu.REG_FILE._01503_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06176_  (.A1(\u_cpu.REG_FILE._01503_ ),
    .A2(\u_cpu.REG_FILE.rf[28][6] ),
    .B1_N(\u_cpu.REG_FILE._01126_ ),
    .X(\u_cpu.REG_FILE._01504_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06177_  (.A1(\u_cpu.REG_FILE._01124_ ),
    .A2(\u_cpu.REG_FILE.rf[29][6] ),
    .B1(\u_cpu.REG_FILE._01504_ ),
    .Y(\u_cpu.REG_FILE._01505_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06178_  (.A1(\u_cpu.REG_FILE._01500_ ),
    .A2(\u_cpu.REG_FILE._01502_ ),
    .B1(\u_cpu.REG_FILE._01505_ ),
    .C1(\u_cpu.REG_FILE._01395_ ),
    .Y(\u_cpu.REG_FILE._01506_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06179_  (.A1(\u_cpu.REG_FILE._01496_ ),
    .A2(\u_cpu.REG_FILE._01499_ ),
    .B1(\u_cpu.REG_FILE._01198_ ),
    .C1(\u_cpu.REG_FILE._01506_ ),
    .Y(\u_cpu.REG_FILE._01507_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06180_  (.A1(\u_cpu.REG_FILE._01206_ ),
    .A2(\u_cpu.REG_FILE.rf[18][6] ),
    .B1(\u_cpu.REG_FILE._01135_ ),
    .Y(\u_cpu.REG_FILE._01508_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06181_  (.A(\u_cpu.REG_FILE._01123_ ),
    .X(\u_cpu.REG_FILE._01509_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06182_  (.A(\u_cpu.REG_FILE.rf[19][6] ),
    .B(\u_cpu.REG_FILE._01509_ ),
    .Y(\u_cpu.REG_FILE._01510_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06183_  (.A1(\u_cpu.REG_FILE._01141_ ),
    .A2(\u_cpu.REG_FILE.rf[16][6] ),
    .B1_N(\u_cpu.REG_FILE._01142_ ),
    .X(\u_cpu.REG_FILE._01511_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06184_  (.A1(\u_cpu.REG_FILE._01140_ ),
    .A2(\u_cpu.REG_FILE.rf[17][6] ),
    .B1(\u_cpu.REG_FILE._01511_ ),
    .Y(\u_cpu.REG_FILE._01512_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06185_  (.A1(\u_cpu.REG_FILE._01508_ ),
    .A2(\u_cpu.REG_FILE._01510_ ),
    .B1(\u_cpu.REG_FILE._01139_ ),
    .C1(\u_cpu.REG_FILE._01512_ ),
    .Y(\u_cpu.REG_FILE._01513_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06186_  (.A(\u_cpu.REG_FILE._01269_ ),
    .B(\u_cpu.REG_FILE.rf[22][6] ),
    .X(\u_cpu.REG_FILE._01514_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06187_  (.A1(\u_cpu.REG_FILE._01146_ ),
    .A2(\u_cpu.REG_FILE.rf[23][6] ),
    .B1(\u_cpu.REG_FILE._01147_ ),
    .C1(\u_cpu.REG_FILE._01514_ ),
    .Y(\u_cpu.REG_FILE._01515_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06188_  (.A1(\u_cpu.REG_FILE._01152_ ),
    .A2(\u_cpu.REG_FILE.rf[20][6] ),
    .B1_N(\u_cpu.REG_FILE._01214_ ),
    .X(\u_cpu.REG_FILE._01516_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06189_  (.A1(\u_cpu.REG_FILE._01151_ ),
    .A2(\u_cpu.REG_FILE.rf[21][6] ),
    .B1(\u_cpu.REG_FILE._01516_ ),
    .Y(\u_cpu.REG_FILE._01517_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06190_  (.A(\u_cpu.REG_FILE._01515_ ),
    .B(\u_cpu.REG_FILE._01517_ ),
    .C(\u_cpu.REG_FILE._01156_ ),
    .Y(\u_cpu.REG_FILE._01518_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06191_  (.A(\u_cpu.REG_FILE._01132_ ),
    .B(\u_cpu.REG_FILE._01513_ ),
    .C(\u_cpu.REG_FILE._01518_ ),
    .Y(\u_cpu.REG_FILE._01519_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06192_  (.A(\u_cpu.REG_FILE._01507_ ),
    .B(\u_cpu.REG_FILE._01519_ ),
    .C(\u_cpu.REG_FILE._01159_ ),
    .Y(\u_cpu.REG_FILE._01520_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06193_  (.A1(\u_cpu.REG_FILE._01026_ ),
    .A2(\u_cpu.REG_FILE._01494_ ),
    .B1(\u_cpu.REG_FILE._01520_ ),
    .C1(\u_cpu.REG_FILE._01165_ ),
    .X(\u_cpu.ALU.SrcA[6] ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06194_  (.A(\u_cpu.REG_FILE._01054_ ),
    .X(\u_cpu.REG_FILE._01521_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06195_  (.A1(\u_cpu.REG_FILE._01279_ ),
    .A2(\u_cpu.REG_FILE.rf[8][7] ),
    .B1_N(\u_cpu.REG_FILE._01521_ ),
    .Y(\u_cpu.REG_FILE._01522_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06196_  (.A(\u_cpu.REG_FILE._01049_ ),
    .X(\u_cpu.REG_FILE._01523_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06197_  (.A_N(\u_cpu.REG_FILE.rf[9][7] ),
    .B(\u_cpu.REG_FILE._01523_ ),
    .X(\u_cpu.REG_FILE._01524_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06198_  (.A(\u_cpu.REG_FILE._01058_ ),
    .X(\u_cpu.REG_FILE._01525_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06199_  (.A1(\u_cpu.REG_FILE._01522_ ),
    .A2(\u_cpu.REG_FILE._01524_ ),
    .B1(\u_cpu.REG_FILE._01525_ ),
    .Y(\u_cpu.REG_FILE._01526_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06200_  (.A(\u_cpu.REG_FILE._01032_ ),
    .X(\u_cpu.REG_FILE._01527_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06201_  (.A(\u_cpu.REG_FILE._01064_ ),
    .X(\u_cpu.REG_FILE._01528_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06202_  (.A(\u_cpu.REG_FILE._01528_ ),
    .B(\u_cpu.REG_FILE.rf[10][7] ),
    .X(\u_cpu.REG_FILE._01529_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06203_  (.A1(\u_cpu.REG_FILE._01137_ ),
    .A2(\u_cpu.REG_FILE.rf[11][7] ),
    .B1(\u_cpu.REG_FILE._01527_ ),
    .C1(\u_cpu.REG_FILE._01529_ ),
    .X(\u_cpu.REG_FILE._01530_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06204_  (.A(\u_cpu.REG_FILE._01125_ ),
    .X(\u_cpu.REG_FILE._01531_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06205_  (.A(\u_cpu.REG_FILE._01531_ ),
    .B(\u_cpu.REG_FILE.rf[12][7] ),
    .Y(\u_cpu.REG_FILE._01532_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06206_  (.A(\u_cpu.REG_FILE._01304_ ),
    .X(\u_cpu.REG_FILE._01533_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06207_  (.A1(\u_cpu.REG_FILE.rf[13][7] ),
    .A2(\u_cpu.REG_FILE._01287_ ),
    .B1_N(\u_cpu.REG_FILE._01533_ ),
    .Y(\u_cpu.REG_FILE._01534_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06208_  (.A(\u_cpu.REG_FILE._01123_ ),
    .X(\u_cpu.REG_FILE._01535_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06209_  (.A(\u_cpu.REG_FILE._01064_ ),
    .X(\u_cpu.REG_FILE._01536_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06210_  (.A(\u_cpu.REG_FILE._01536_ ),
    .B(\u_cpu.REG_FILE.rf[14][7] ),
    .X(\u_cpu.REG_FILE._01537_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06211_  (.A1(\u_cpu.REG_FILE._01535_ ),
    .A2(\u_cpu.REG_FILE.rf[15][7] ),
    .B1(\u_cpu.REG_FILE._01527_ ),
    .C1(\u_cpu.REG_FILE._01537_ ),
    .Y(\u_cpu.REG_FILE._01538_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06212_  (.A1(\u_cpu.REG_FILE._01532_ ),
    .A2(\u_cpu.REG_FILE._01534_ ),
    .B1(\u_cpu.REG_FILE._01129_ ),
    .C1(\u_cpu.REG_FILE._01538_ ),
    .Y(\u_cpu.REG_FILE._01539_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06213_  (.A1(\u_cpu.REG_FILE._01526_ ),
    .A2(\u_cpu.REG_FILE._01530_ ),
    .B1(\u_cpu.REG_FILE._01117_ ),
    .C1(\u_cpu.REG_FILE._01539_ ),
    .X(\u_cpu.REG_FILE._01540_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06214_  (.A(\u_cpu.REG_FILE._01089_ ),
    .X(\u_cpu.REG_FILE._01541_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06215_  (.A_N(\u_cpu.REG_FILE.rf[1][7] ),
    .B(\u_cpu.REG_FILE._01074_ ),
    .X(\u_cpu.REG_FILE._01542_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06216_  (.A1(\u_cpu.REG_FILE._01093_ ),
    .A2(\u_cpu.REG_FILE.rf[0][7] ),
    .B1_N(\u_cpu.REG_FILE._01305_ ),
    .Y(\u_cpu.REG_FILE._01543_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06217_  (.A(\u_cpu.REG_FILE.rf[3][7] ),
    .B_N(\u_cpu.REG_FILE._01310_ ),
    .X(\u_cpu.REG_FILE._01544_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06218_  (.A1(\u_cpu.REG_FILE._01308_ ),
    .A2(\u_cpu.REG_FILE.rf[2][7] ),
    .B1(\u_cpu.REG_FILE._01309_ ),
    .C1(\u_cpu.REG_FILE._01544_ ),
    .Y(\u_cpu.REG_FILE._01545_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06219_  (.A1(\u_cpu.REG_FILE._01542_ ),
    .A2(\u_cpu.REG_FILE._01543_ ),
    .B1(\u_cpu.REG_FILE._01307_ ),
    .C1(\u_cpu.REG_FILE._01545_ ),
    .Y(\u_cpu.REG_FILE._01546_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06220_  (.A(\u_cpu.REG_FILE._01049_ ),
    .X(\u_cpu.REG_FILE._01547_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06221_  (.A_N(\u_cpu.REG_FILE.rf[5][7] ),
    .B(\u_cpu.REG_FILE._01547_ ),
    .X(\u_cpu.REG_FILE._01548_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06222_  (.A(\u_cpu.REG_FILE._01052_ ),
    .X(\u_cpu.REG_FILE._01549_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06223_  (.A(\u_cpu.REG_FILE._01304_ ),
    .X(\u_cpu.REG_FILE._01550_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06224_  (.A1(\u_cpu.REG_FILE._01549_ ),
    .A2(\u_cpu.REG_FILE.rf[4][7] ),
    .B1_N(\u_cpu.REG_FILE._01550_ ),
    .Y(\u_cpu.REG_FILE._01551_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06225_  (.A(\u_cpu.REG_FILE._01045_ ),
    .X(\u_cpu.REG_FILE._01552_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06226_  (.A(\u_cpu.REG_FILE._01054_ ),
    .X(\u_cpu.REG_FILE._01553_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.REG_FILE._06227_  (.A1(\u_cpu.REG_FILE._01262_ ),
    .A2(\u_cpu.REG_FILE.rf[6][7] ),
    .B1(\u_cpu.REG_FILE._01553_ ),
    .X(\u_cpu.REG_FILE._01554_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06228_  (.A1(\u_cpu.REG_FILE.rf[7][7] ),
    .A2(\u_cpu.REG_FILE._01298_ ),
    .B1(\u_cpu.REG_FILE._01554_ ),
    .Y(\u_cpu.REG_FILE._01555_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06229_  (.A1(\u_cpu.REG_FILE._01548_ ),
    .A2(\u_cpu.REG_FILE._01551_ ),
    .B1(\u_cpu.REG_FILE._01552_ ),
    .C1(\u_cpu.REG_FILE._01555_ ),
    .Y(\u_cpu.REG_FILE._01556_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._06230_  (.A1(\u_cpu.REG_FILE._01541_ ),
    .A2(\u_cpu.REG_FILE._01546_ ),
    .A3(\u_cpu.REG_FILE._01556_ ),
    .B1(\u_cpu.REG_FILE._01024_ ),
    .X(\u_cpu.REG_FILE._01557_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06231_  (.A(\u_cpu.REG_FILE.rf[27][7] ),
    .B_N(\u_cpu.REG_FILE._01108_ ),
    .X(\u_cpu.REG_FILE._01558_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06232_  (.A1(\u_cpu.REG_FILE._01105_ ),
    .A2(\u_cpu.REG_FILE.rf[26][7] ),
    .B1(\u_cpu.REG_FILE._01107_ ),
    .C1(\u_cpu.REG_FILE._01558_ ),
    .X(\u_cpu.REG_FILE._01559_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06233_  (.A1(\u_cpu.REG_FILE._01447_ ),
    .A2(\u_cpu.REG_FILE.rf[24][7] ),
    .B1_N(\u_cpu.REG_FILE._01112_ ),
    .X(\u_cpu.REG_FILE._01560_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06234_  (.A(\u_cpu.REG_FILE.rf[25][7] ),
    .B_N(\u_cpu.REG_FILE._01194_ ),
    .X(\u_cpu.REG_FILE._01561_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._06235_  (.A1(\u_cpu.REG_FILE._01560_ ),
    .A2(\u_cpu.REG_FILE._01561_ ),
    .B1(\u_cpu.REG_FILE._01196_ ),
    .X(\u_cpu.REG_FILE._01562_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06236_  (.A(\u_cpu.REG_FILE._01390_ ),
    .B(\u_cpu.REG_FILE.rf[30][7] ),
    .Y(\u_cpu.REG_FILE._01563_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06237_  (.A1(\u_cpu.REG_FILE.rf[31][7] ),
    .A2(\u_cpu.REG_FILE._01200_ ),
    .B1(\u_cpu.REG_FILE._01501_ ),
    .Y(\u_cpu.REG_FILE._01564_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06238_  (.A1(\u_cpu.REG_FILE._01503_ ),
    .A2(\u_cpu.REG_FILE.rf[28][7] ),
    .B1_N(\u_cpu.REG_FILE._01126_ ),
    .X(\u_cpu.REG_FILE._01565_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06239_  (.A1(\u_cpu.REG_FILE._01124_ ),
    .A2(\u_cpu.REG_FILE.rf[29][7] ),
    .B1(\u_cpu.REG_FILE._01565_ ),
    .Y(\u_cpu.REG_FILE._01566_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06240_  (.A1(\u_cpu.REG_FILE._01563_ ),
    .A2(\u_cpu.REG_FILE._01564_ ),
    .B1(\u_cpu.REG_FILE._01566_ ),
    .C1(\u_cpu.REG_FILE._01395_ ),
    .Y(\u_cpu.REG_FILE._01567_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06241_  (.A1(\u_cpu.REG_FILE._01559_ ),
    .A2(\u_cpu.REG_FILE._01562_ ),
    .B1(\u_cpu.REG_FILE._01198_ ),
    .C1(\u_cpu.REG_FILE._01567_ ),
    .Y(\u_cpu.REG_FILE._01568_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06242_  (.A(\u_cpu.REG_FILE._01089_ ),
    .X(\u_cpu.REG_FILE._01569_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06243_  (.A1(\u_cpu.REG_FILE._01206_ ),
    .A2(\u_cpu.REG_FILE.rf[18][7] ),
    .B1(\u_cpu.REG_FILE._01135_ ),
    .Y(\u_cpu.REG_FILE._01570_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06244_  (.A(\u_cpu.REG_FILE.rf[19][7] ),
    .B(\u_cpu.REG_FILE._01509_ ),
    .Y(\u_cpu.REG_FILE._01571_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06245_  (.A1(\u_cpu.REG_FILE._01141_ ),
    .A2(\u_cpu.REG_FILE.rf[16][7] ),
    .B1_N(\u_cpu.REG_FILE._01142_ ),
    .X(\u_cpu.REG_FILE._01572_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06246_  (.A1(\u_cpu.REG_FILE._01140_ ),
    .A2(\u_cpu.REG_FILE.rf[17][7] ),
    .B1(\u_cpu.REG_FILE._01572_ ),
    .Y(\u_cpu.REG_FILE._01573_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06247_  (.A1(\u_cpu.REG_FILE._01570_ ),
    .A2(\u_cpu.REG_FILE._01571_ ),
    .B1(\u_cpu.REG_FILE._01139_ ),
    .C1(\u_cpu.REG_FILE._01573_ ),
    .Y(\u_cpu.REG_FILE._01574_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06248_  (.A(\u_cpu.REG_FILE._01260_ ),
    .B(\u_cpu.REG_FILE.rf[20][7] ),
    .Y(\u_cpu.REG_FILE._01575_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06249_  (.A_N(\u_cpu.REG_FILE.rf[21][7] ),
    .B(\u_cpu.REG_FILE._01262_ ),
    .X(\u_cpu.REG_FILE._01576_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06250_  (.A(\u_cpu.REG_FILE.rf[23][7] ),
    .B_N(\u_cpu.REG_FILE._01408_ ),
    .X(\u_cpu.REG_FILE._01577_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06251_  (.A1(\u_cpu.REG_FILE._01260_ ),
    .A2(\u_cpu.REG_FILE.rf[22][7] ),
    .B1(\u_cpu.REG_FILE._01400_ ),
    .C1(\u_cpu.REG_FILE._01577_ ),
    .Y(\u_cpu.REG_FILE._01578_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._06252_  (.A1(\u_cpu.REG_FILE._01259_ ),
    .A2(\u_cpu.REG_FILE._01575_ ),
    .A3(\u_cpu.REG_FILE._01576_ ),
    .B1(\u_cpu.REG_FILE._01115_ ),
    .C1(\u_cpu.REG_FILE._01578_ ),
    .Y(\u_cpu.REG_FILE._01579_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06253_  (.A(\u_cpu.REG_FILE._01569_ ),
    .B(\u_cpu.REG_FILE._01574_ ),
    .C(\u_cpu.REG_FILE._01579_ ),
    .Y(\u_cpu.REG_FILE._01580_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06254_  (.A(\u_cpu.REG_FILE._01568_ ),
    .B(\u_cpu.REG_FILE._01580_ ),
    .C(\u_cpu.REG_FILE._01159_ ),
    .Y(\u_cpu.REG_FILE._01581_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06255_  (.A1(\u_cpu.REG_FILE._01540_ ),
    .A2(\u_cpu.REG_FILE._01557_ ),
    .B1(\u_cpu.REG_FILE._01581_ ),
    .C1(\u_cpu.REG_FILE._01165_ ),
    .X(\u_cpu.ALU.SrcA[7] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06256_  (.A(\u_cpu.REG_FILE.rf[15][8] ),
    .B_N(\u_cpu.REG_FILE._01034_ ),
    .X(\u_cpu.REG_FILE._01582_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06257_  (.A1(\u_cpu.REG_FILE._01351_ ),
    .A2(\u_cpu.REG_FILE.rf[14][8] ),
    .B1(\u_cpu.REG_FILE._01352_ ),
    .C1(\u_cpu.REG_FILE._01582_ ),
    .Y(\u_cpu.REG_FILE._01583_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06258_  (.A(\u_cpu.REG_FILE._01073_ ),
    .X(\u_cpu.REG_FILE._01584_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06259_  (.A1(\u_cpu.REG_FILE._01584_ ),
    .A2(\u_cpu.REG_FILE.rf[12][8] ),
    .B1_N(\u_cpu.REG_FILE._01042_ ),
    .X(\u_cpu.REG_FILE._01585_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06260_  (.A1(\u_cpu.REG_FILE._01039_ ),
    .A2(\u_cpu.REG_FILE.rf[13][8] ),
    .B1(\u_cpu.REG_FILE._01585_ ),
    .Y(\u_cpu.REG_FILE._01586_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06261_  (.A(\u_cpu.REG_FILE._01583_ ),
    .B(\u_cpu.REG_FILE._01586_ ),
    .C(\u_cpu.REG_FILE._01047_ ),
    .Y(\u_cpu.REG_FILE._01587_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06262_  (.A_N(\u_cpu.REG_FILE.rf[9][8] ),
    .B(\u_cpu.REG_FILE._01050_ ),
    .X(\u_cpu.REG_FILE._01588_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06263_  (.A1(\u_cpu.REG_FILE._01475_ ),
    .A2(\u_cpu.REG_FILE.rf[8][8] ),
    .B1_N(\u_cpu.REG_FILE._01055_ ),
    .Y(\u_cpu.REG_FILE._01589_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06264_  (.A(\u_cpu.REG_FILE._01040_ ),
    .X(\u_cpu.REG_FILE._01590_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06265_  (.A(\u_cpu.REG_FILE.rf[11][8] ),
    .B_N(\u_cpu.REG_FILE._01590_ ),
    .X(\u_cpu.REG_FILE._01591_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06266_  (.A1(\u_cpu.REG_FILE._01425_ ),
    .A2(\u_cpu.REG_FILE.rf[10][8] ),
    .B1(\u_cpu.REG_FILE._01360_ ),
    .C1(\u_cpu.REG_FILE._01591_ ),
    .Y(\u_cpu.REG_FILE._01592_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06267_  (.A1(\u_cpu.REG_FILE._01588_ ),
    .A2(\u_cpu.REG_FILE._01589_ ),
    .B1(\u_cpu.REG_FILE._01424_ ),
    .C1(\u_cpu.REG_FILE._01592_ ),
    .Y(\u_cpu.REG_FILE._01593_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06268_  (.A(\u_cpu.REG_FILE._01587_ ),
    .B(\u_cpu.REG_FILE._01593_ ),
    .C(\u_cpu.REG_FILE._01070_ ),
    .Y(\u_cpu.REG_FILE._01594_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06269_  (.A(\u_cpu.REG_FILE.rf[5][8] ),
    .Y(\u_cpu.REG_FILE._01595_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06270_  (.A1(\u_cpu.REG_FILE._01431_ ),
    .A2(\u_cpu.REG_FILE.rf[4][8] ),
    .B1_N(\u_cpu.REG_FILE._01482_ ),
    .Y(\u_cpu.REG_FILE._01596_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._06271_  (.A1(\u_cpu.REG_FILE._01595_ ),
    .A2(\u_cpu.REG_FILE._01075_ ),
    .B1(\u_cpu.REG_FILE._01596_ ),
    .Y(\u_cpu.REG_FILE._01597_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06272_  (.A(\u_cpu.REG_FILE._01082_ ),
    .X(\u_cpu.REG_FILE._01598_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06273_  (.A1(\u_cpu.REG_FILE._01434_ ),
    .A2(\u_cpu.REG_FILE.rf[6][8] ),
    .B1(\u_cpu.REG_FILE._01598_ ),
    .Y(\u_cpu.REG_FILE._01599_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06274_  (.A_N(\u_cpu.REG_FILE.rf[7][8] ),
    .B(\u_cpu.REG_FILE._01085_ ),
    .X(\u_cpu.REG_FILE._01600_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06275_  (.A(\u_cpu.REG_FILE._01045_ ),
    .X(\u_cpu.REG_FILE._01601_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06276_  (.A1(\u_cpu.REG_FILE._01599_ ),
    .A2(\u_cpu.REG_FILE._01600_ ),
    .B1(\u_cpu.REG_FILE._01601_ ),
    .Y(\u_cpu.REG_FILE._01602_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06277_  (.A(\u_cpu.REG_FILE._01089_ ),
    .X(\u_cpu.REG_FILE._01603_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06278_  (.A_N(\u_cpu.REG_FILE.rf[1][8] ),
    .B(\u_cpu.REG_FILE._01091_ ),
    .X(\u_cpu.REG_FILE._01604_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06279_  (.A1(\u_cpu.REG_FILE._01372_ ),
    .A2(\u_cpu.REG_FILE.rf[0][8] ),
    .B1_N(\u_cpu.REG_FILE._01094_ ),
    .Y(\u_cpu.REG_FILE._01605_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06280_  (.A(\u_cpu.REG_FILE.rf[3][8] ),
    .B_N(\u_cpu.REG_FILE._01241_ ),
    .X(\u_cpu.REG_FILE._01606_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06281_  (.A1(\u_cpu.REG_FILE._01097_ ),
    .A2(\u_cpu.REG_FILE.rf[2][8] ),
    .B1(\u_cpu.REG_FILE._01240_ ),
    .C1(\u_cpu.REG_FILE._01606_ ),
    .Y(\u_cpu.REG_FILE._01607_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06282_  (.A1(\u_cpu.REG_FILE._01604_ ),
    .A2(\u_cpu.REG_FILE._01605_ ),
    .B1(\u_cpu.REG_FILE._01096_ ),
    .C1(\u_cpu.REG_FILE._01607_ ),
    .Y(\u_cpu.REG_FILE._01608_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06283_  (.A1(\u_cpu.REG_FILE._01597_ ),
    .A2(\u_cpu.REG_FILE._01602_ ),
    .B1(\u_cpu.REG_FILE._01603_ ),
    .C1(\u_cpu.REG_FILE._01608_ ),
    .Y(\u_cpu.REG_FILE._01609_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._06284_  (.A(\u_cpu.REG_FILE._01594_ ),
    .B(\u_cpu.REG_FILE._01609_ ),
    .Y(\u_cpu.REG_FILE._01610_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06285_  (.A(\u_cpu.REG_FILE._01031_ ),
    .X(\u_cpu.REG_FILE._01611_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06286_  (.A1(\u_cpu.REG_FILE._01379_ ),
    .A2(\u_cpu.REG_FILE.rf[24][8] ),
    .B1_N(\u_cpu.REG_FILE._01611_ ),
    .Y(\u_cpu.REG_FILE._01612_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06287_  (.A_N(\u_cpu.REG_FILE.rf[25][8] ),
    .B(\u_cpu.REG_FILE._01382_ ),
    .X(\u_cpu.REG_FILE._01613_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06288_  (.A1(\u_cpu.REG_FILE._01612_ ),
    .A2(\u_cpu.REG_FILE._01613_ ),
    .B1(\u_cpu.REG_FILE._01384_ ),
    .Y(\u_cpu.REG_FILE._01614_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06289_  (.A(\u_cpu.REG_FILE._01340_ ),
    .B(\u_cpu.REG_FILE.rf[26][8] ),
    .X(\u_cpu.REG_FILE._01615_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06290_  (.A1(\u_cpu.REG_FILE._01386_ ),
    .A2(\u_cpu.REG_FILE.rf[27][8] ),
    .B1(\u_cpu.REG_FILE._01387_ ),
    .C1(\u_cpu.REG_FILE._01615_ ),
    .X(\u_cpu.REG_FILE._01616_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06291_  (.A(\u_cpu.REG_FILE._01549_ ),
    .B(\u_cpu.REG_FILE.rf[30][8] ),
    .Y(\u_cpu.REG_FILE._01617_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06292_  (.A(\u_cpu.REG_FILE._01142_ ),
    .X(\u_cpu.REG_FILE._01618_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06293_  (.A1(\u_cpu.REG_FILE.rf[31][8] ),
    .A2(\u_cpu.REG_FILE._01327_ ),
    .B1(\u_cpu.REG_FILE._01618_ ),
    .Y(\u_cpu.REG_FILE._01619_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06294_  (.A(\u_cpu.REG_FILE._01148_ ),
    .X(\u_cpu.REG_FILE._01620_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06295_  (.A(\u_cpu.REG_FILE._01620_ ),
    .B(\u_cpu.REG_FILE.rf[28][8] ),
    .Y(\u_cpu.REG_FILE._01621_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06296_  (.A1(\u_cpu.REG_FILE.rf[29][8] ),
    .A2(\u_cpu.REG_FILE._01321_ ),
    .B1_N(\u_cpu.REG_FILE._01521_ ),
    .Y(\u_cpu.REG_FILE._01622_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._06297_  (.A1(\u_cpu.REG_FILE._01617_ ),
    .A2(\u_cpu.REG_FILE._01619_ ),
    .B1(\u_cpu.REG_FILE._01621_ ),
    .B2(\u_cpu.REG_FILE._01622_ ),
    .C1(\u_cpu.REG_FILE._01333_ ),
    .Y(\u_cpu.REG_FILE._01623_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06298_  (.A1(\u_cpu.REG_FILE._01614_ ),
    .A2(\u_cpu.REG_FILE._01616_ ),
    .B1(\u_cpu.REG_FILE._01198_ ),
    .C1(\u_cpu.REG_FILE._01623_ ),
    .Y(\u_cpu.REG_FILE._01624_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06299_  (.A1(\u_cpu.REG_FILE._01206_ ),
    .A2(\u_cpu.REG_FILE.rf[18][8] ),
    .B1(\u_cpu.REG_FILE._01135_ ),
    .Y(\u_cpu.REG_FILE._01625_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06300_  (.A(\u_cpu.REG_FILE.rf[19][8] ),
    .B(\u_cpu.REG_FILE._01509_ ),
    .Y(\u_cpu.REG_FILE._01626_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06301_  (.A1(\u_cpu.REG_FILE._01141_ ),
    .A2(\u_cpu.REG_FILE.rf[16][8] ),
    .B1_N(\u_cpu.REG_FILE._01142_ ),
    .X(\u_cpu.REG_FILE._01627_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06302_  (.A1(\u_cpu.REG_FILE._01140_ ),
    .A2(\u_cpu.REG_FILE.rf[17][8] ),
    .B1(\u_cpu.REG_FILE._01627_ ),
    .Y(\u_cpu.REG_FILE._01628_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06303_  (.A1(\u_cpu.REG_FILE._01625_ ),
    .A2(\u_cpu.REG_FILE._01626_ ),
    .B1(\u_cpu.REG_FILE._01139_ ),
    .C1(\u_cpu.REG_FILE._01628_ ),
    .Y(\u_cpu.REG_FILE._01629_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06304_  (.A(\u_cpu.REG_FILE._01269_ ),
    .B(\u_cpu.REG_FILE.rf[22][8] ),
    .X(\u_cpu.REG_FILE._01630_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06305_  (.A1(\u_cpu.REG_FILE._01146_ ),
    .A2(\u_cpu.REG_FILE.rf[23][8] ),
    .B1(\u_cpu.REG_FILE._01147_ ),
    .C1(\u_cpu.REG_FILE._01630_ ),
    .Y(\u_cpu.REG_FILE._01631_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06306_  (.A(\u_cpu.REG_FILE._01064_ ),
    .X(\u_cpu.REG_FILE._01632_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06307_  (.A1(\u_cpu.REG_FILE._01632_ ),
    .A2(\u_cpu.REG_FILE.rf[20][8] ),
    .B1_N(\u_cpu.REG_FILE._01214_ ),
    .X(\u_cpu.REG_FILE._01633_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06308_  (.A1(\u_cpu.REG_FILE._01151_ ),
    .A2(\u_cpu.REG_FILE.rf[21][8] ),
    .B1(\u_cpu.REG_FILE._01633_ ),
    .Y(\u_cpu.REG_FILE._01634_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06309_  (.A(\u_cpu.REG_FILE._01631_ ),
    .B(\u_cpu.REG_FILE._01634_ ),
    .C(\u_cpu.REG_FILE._01156_ ),
    .Y(\u_cpu.REG_FILE._01635_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06310_  (.A(\u_cpu.REG_FILE._01569_ ),
    .B(\u_cpu.REG_FILE._01629_ ),
    .C(\u_cpu.REG_FILE._01635_ ),
    .Y(\u_cpu.REG_FILE._01636_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06311_  (.A(\u_cpu.REG_FILE._01624_ ),
    .B(\u_cpu.REG_FILE._01636_ ),
    .C(\u_cpu.REG_FILE._01159_ ),
    .Y(\u_cpu.REG_FILE._01637_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06312_  (.A1(\u_cpu.REG_FILE._01026_ ),
    .A2(\u_cpu.REG_FILE._01610_ ),
    .B1(\u_cpu.REG_FILE._01637_ ),
    .C1(\u_cpu.REG_FILE._01165_ ),
    .X(\u_cpu.ALU.SrcA[8] ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06313_  (.A1(\u_cpu.REG_FILE._01279_ ),
    .A2(\u_cpu.REG_FILE.rf[8][9] ),
    .B1_N(\u_cpu.REG_FILE._01521_ ),
    .Y(\u_cpu.REG_FILE._01638_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06314_  (.A_N(\u_cpu.REG_FILE.rf[9][9] ),
    .B(\u_cpu.REG_FILE._01523_ ),
    .X(\u_cpu.REG_FILE._01639_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06315_  (.A1(\u_cpu.REG_FILE._01638_ ),
    .A2(\u_cpu.REG_FILE._01639_ ),
    .B1(\u_cpu.REG_FILE._01525_ ),
    .Y(\u_cpu.REG_FILE._01640_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06316_  (.A(\u_cpu.REG_FILE._01528_ ),
    .B(\u_cpu.REG_FILE.rf[10][9] ),
    .X(\u_cpu.REG_FILE._01641_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06317_  (.A1(\u_cpu.REG_FILE._01137_ ),
    .A2(\u_cpu.REG_FILE.rf[11][9] ),
    .B1(\u_cpu.REG_FILE._01527_ ),
    .C1(\u_cpu.REG_FILE._01641_ ),
    .X(\u_cpu.REG_FILE._01642_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06318_  (.A(\u_cpu.REG_FILE._01118_ ),
    .B(\u_cpu.REG_FILE.rf[12][9] ),
    .Y(\u_cpu.REG_FILE._01643_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06319_  (.A1(\u_cpu.REG_FILE.rf[13][9] ),
    .A2(\u_cpu.REG_FILE._01287_ ),
    .B1_N(\u_cpu.REG_FILE._01305_ ),
    .Y(\u_cpu.REG_FILE._01644_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06320_  (.A(\u_cpu.REG_FILE._01536_ ),
    .B(\u_cpu.REG_FILE.rf[14][9] ),
    .X(\u_cpu.REG_FILE._01645_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06321_  (.A1(\u_cpu.REG_FILE._01535_ ),
    .A2(\u_cpu.REG_FILE.rf[15][9] ),
    .B1(\u_cpu.REG_FILE._01527_ ),
    .C1(\u_cpu.REG_FILE._01645_ ),
    .Y(\u_cpu.REG_FILE._01646_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06322_  (.A1(\u_cpu.REG_FILE._01643_ ),
    .A2(\u_cpu.REG_FILE._01644_ ),
    .B1(\u_cpu.REG_FILE._01129_ ),
    .C1(\u_cpu.REG_FILE._01646_ ),
    .Y(\u_cpu.REG_FILE._01647_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06323_  (.A1(\u_cpu.REG_FILE._01640_ ),
    .A2(\u_cpu.REG_FILE._01642_ ),
    .B1(\u_cpu.REG_FILE._01117_ ),
    .C1(\u_cpu.REG_FILE._01647_ ),
    .X(\u_cpu.REG_FILE._01648_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06324_  (.A_N(\u_cpu.REG_FILE.rf[1][9] ),
    .B(\u_cpu.REG_FILE._01074_ ),
    .X(\u_cpu.REG_FILE._01649_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06325_  (.A1(\u_cpu.REG_FILE._01093_ ),
    .A2(\u_cpu.REG_FILE.rf[0][9] ),
    .B1_N(\u_cpu.REG_FILE._01305_ ),
    .Y(\u_cpu.REG_FILE._01650_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06326_  (.A(\u_cpu.REG_FILE.rf[3][9] ),
    .B_N(\u_cpu.REG_FILE._01310_ ),
    .X(\u_cpu.REG_FILE._01651_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06327_  (.A1(\u_cpu.REG_FILE._01308_ ),
    .A2(\u_cpu.REG_FILE.rf[2][9] ),
    .B1(\u_cpu.REG_FILE._01309_ ),
    .C1(\u_cpu.REG_FILE._01651_ ),
    .Y(\u_cpu.REG_FILE._01652_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06328_  (.A1(\u_cpu.REG_FILE._01649_ ),
    .A2(\u_cpu.REG_FILE._01650_ ),
    .B1(\u_cpu.REG_FILE._01307_ ),
    .C1(\u_cpu.REG_FILE._01652_ ),
    .Y(\u_cpu.REG_FILE._01653_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06329_  (.A_N(\u_cpu.REG_FILE.rf[5][9] ),
    .B(\u_cpu.REG_FILE._01547_ ),
    .X(\u_cpu.REG_FILE._01654_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06330_  (.A1(\u_cpu.REG_FILE._01549_ ),
    .A2(\u_cpu.REG_FILE.rf[4][9] ),
    .B1_N(\u_cpu.REG_FILE._01550_ ),
    .Y(\u_cpu.REG_FILE._01655_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.REG_FILE._06331_  (.A1(\u_cpu.REG_FILE._01262_ ),
    .A2(\u_cpu.REG_FILE.rf[6][9] ),
    .B1(\u_cpu.REG_FILE._01553_ ),
    .X(\u_cpu.REG_FILE._01656_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06332_  (.A1(\u_cpu.REG_FILE.rf[7][9] ),
    .A2(\u_cpu.REG_FILE._01287_ ),
    .B1(\u_cpu.REG_FILE._01656_ ),
    .Y(\u_cpu.REG_FILE._01657_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06333_  (.A1(\u_cpu.REG_FILE._01654_ ),
    .A2(\u_cpu.REG_FILE._01655_ ),
    .B1(\u_cpu.REG_FILE._01552_ ),
    .C1(\u_cpu.REG_FILE._01657_ ),
    .Y(\u_cpu.REG_FILE._01658_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._06334_  (.A1(\u_cpu.REG_FILE._01541_ ),
    .A2(\u_cpu.REG_FILE._01653_ ),
    .A3(\u_cpu.REG_FILE._01658_ ),
    .B1(\u_cpu.REG_FILE._01024_ ),
    .X(\u_cpu.REG_FILE._01659_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06335_  (.A(\u_cpu.REG_FILE._01106_ ),
    .X(\u_cpu.REG_FILE._01660_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06336_  (.A(\u_cpu.REG_FILE.rf[27][9] ),
    .B_N(\u_cpu.REG_FILE._01108_ ),
    .X(\u_cpu.REG_FILE._01661_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06337_  (.A1(\u_cpu.REG_FILE._01105_ ),
    .A2(\u_cpu.REG_FILE.rf[26][9] ),
    .B1(\u_cpu.REG_FILE._01660_ ),
    .C1(\u_cpu.REG_FILE._01661_ ),
    .X(\u_cpu.REG_FILE._01662_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06338_  (.A1(\u_cpu.REG_FILE._01447_ ),
    .A2(\u_cpu.REG_FILE.rf[24][9] ),
    .B1_N(\u_cpu.REG_FILE._01112_ ),
    .X(\u_cpu.REG_FILE._01663_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06339_  (.A(\u_cpu.REG_FILE.rf[25][9] ),
    .B_N(\u_cpu.REG_FILE._01194_ ),
    .X(\u_cpu.REG_FILE._01664_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._06340_  (.A1(\u_cpu.REG_FILE._01663_ ),
    .A2(\u_cpu.REG_FILE._01664_ ),
    .B1(\u_cpu.REG_FILE._01196_ ),
    .X(\u_cpu.REG_FILE._01665_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06341_  (.A(\u_cpu.REG_FILE._01390_ ),
    .B(\u_cpu.REG_FILE.rf[30][9] ),
    .Y(\u_cpu.REG_FILE._01666_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06342_  (.A1(\u_cpu.REG_FILE.rf[31][9] ),
    .A2(\u_cpu.REG_FILE._01200_ ),
    .B1(\u_cpu.REG_FILE._01501_ ),
    .Y(\u_cpu.REG_FILE._01667_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06343_  (.A(\u_cpu.REG_FILE._01123_ ),
    .X(\u_cpu.REG_FILE._01668_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06344_  (.A1(\u_cpu.REG_FILE._01503_ ),
    .A2(\u_cpu.REG_FILE.rf[28][9] ),
    .B1_N(\u_cpu.REG_FILE._01126_ ),
    .X(\u_cpu.REG_FILE._01669_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06345_  (.A1(\u_cpu.REG_FILE._01668_ ),
    .A2(\u_cpu.REG_FILE.rf[29][9] ),
    .B1(\u_cpu.REG_FILE._01669_ ),
    .Y(\u_cpu.REG_FILE._01670_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06346_  (.A1(\u_cpu.REG_FILE._01666_ ),
    .A2(\u_cpu.REG_FILE._01667_ ),
    .B1(\u_cpu.REG_FILE._01670_ ),
    .C1(\u_cpu.REG_FILE._01395_ ),
    .Y(\u_cpu.REG_FILE._01671_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06347_  (.A1(\u_cpu.REG_FILE._01662_ ),
    .A2(\u_cpu.REG_FILE._01665_ ),
    .B1(\u_cpu.REG_FILE._01198_ ),
    .C1(\u_cpu.REG_FILE._01671_ ),
    .Y(\u_cpu.REG_FILE._01672_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06348_  (.A(\u_cpu.REG_FILE._01379_ ),
    .B(\u_cpu.REG_FILE.rf[16][9] ),
    .Y(\u_cpu.REG_FILE._01673_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06349_  (.A_N(\u_cpu.REG_FILE.rf[17][9] ),
    .B(\u_cpu.REG_FILE._01029_ ),
    .X(\u_cpu.REG_FILE._01674_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.REG_FILE._06350_  (.A1(\u_cpu.REG_FILE._01060_ ),
    .A2(\u_cpu.REG_FILE.rf[18][9] ),
    .B1(\u_cpu.REG_FILE._01239_ ),
    .X(\u_cpu.REG_FILE._01675_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06351_  (.A1(\u_cpu.REG_FILE.rf[19][9] ),
    .A2(\u_cpu.REG_FILE._01265_ ),
    .B1(\u_cpu.REG_FILE._01675_ ),
    .Y(\u_cpu.REG_FILE._01676_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._06352_  (.A1(\u_cpu.REG_FILE._01033_ ),
    .A2(\u_cpu.REG_FILE._01673_ ),
    .A3(\u_cpu.REG_FILE._01674_ ),
    .B1(\u_cpu.REG_FILE._01058_ ),
    .C1(\u_cpu.REG_FILE._01676_ ),
    .Y(\u_cpu.REG_FILE._01677_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06353_  (.A(\u_cpu.REG_FILE._01269_ ),
    .B(\u_cpu.REG_FILE.rf[22][9] ),
    .X(\u_cpu.REG_FILE._01678_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06354_  (.A1(\u_cpu.REG_FILE._01146_ ),
    .A2(\u_cpu.REG_FILE.rf[23][9] ),
    .B1(\u_cpu.REG_FILE._01147_ ),
    .C1(\u_cpu.REG_FILE._01678_ ),
    .Y(\u_cpu.REG_FILE._01679_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06355_  (.A1(\u_cpu.REG_FILE._01632_ ),
    .A2(\u_cpu.REG_FILE.rf[20][9] ),
    .B1_N(\u_cpu.REG_FILE._01214_ ),
    .X(\u_cpu.REG_FILE._01680_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06356_  (.A1(\u_cpu.REG_FILE._01151_ ),
    .A2(\u_cpu.REG_FILE.rf[21][9] ),
    .B1(\u_cpu.REG_FILE._01680_ ),
    .Y(\u_cpu.REG_FILE._01681_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06357_  (.A(\u_cpu.REG_FILE._01679_ ),
    .B(\u_cpu.REG_FILE._01681_ ),
    .C(\u_cpu.REG_FILE._01156_ ),
    .Y(\u_cpu.REG_FILE._01682_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06358_  (.A(\u_cpu.REG_FILE._01569_ ),
    .B(\u_cpu.REG_FILE._01677_ ),
    .C(\u_cpu.REG_FILE._01682_ ),
    .Y(\u_cpu.REG_FILE._01683_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06359_  (.A(\u_cpu.REG_FILE._01024_ ),
    .X(\u_cpu.REG_FILE._01684_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06360_  (.A(\u_cpu.REG_FILE._01672_ ),
    .B(\u_cpu.REG_FILE._01683_ ),
    .C(\u_cpu.REG_FILE._01684_ ),
    .Y(\u_cpu.REG_FILE._01685_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06361_  (.A1(\u_cpu.REG_FILE._01648_ ),
    .A2(\u_cpu.REG_FILE._01659_ ),
    .B1(\u_cpu.REG_FILE._01685_ ),
    .C1(\u_cpu.REG_FILE._01165_ ),
    .X(\u_cpu.ALU.SrcA[9] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06362_  (.A(\u_cpu.REG_FILE.rf[15][10] ),
    .B_N(\u_cpu.REG_FILE._01034_ ),
    .X(\u_cpu.REG_FILE._01686_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06363_  (.A1(\u_cpu.REG_FILE._01351_ ),
    .A2(\u_cpu.REG_FILE.rf[14][10] ),
    .B1(\u_cpu.REG_FILE._01352_ ),
    .C1(\u_cpu.REG_FILE._01686_ ),
    .Y(\u_cpu.REG_FILE._01687_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06364_  (.A1(\u_cpu.REG_FILE._01584_ ),
    .A2(\u_cpu.REG_FILE.rf[12][10] ),
    .B1_N(\u_cpu.REG_FILE._01042_ ),
    .X(\u_cpu.REG_FILE._01688_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06365_  (.A1(\u_cpu.REG_FILE._01039_ ),
    .A2(\u_cpu.REG_FILE.rf[13][10] ),
    .B1(\u_cpu.REG_FILE._01688_ ),
    .Y(\u_cpu.REG_FILE._01689_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06366_  (.A(\u_cpu.REG_FILE._01046_ ),
    .X(\u_cpu.REG_FILE._01690_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06367_  (.A(\u_cpu.REG_FILE._01687_ ),
    .B(\u_cpu.REG_FILE._01689_ ),
    .C(\u_cpu.REG_FILE._01690_ ),
    .Y(\u_cpu.REG_FILE._01691_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06368_  (.A_N(\u_cpu.REG_FILE.rf[9][10] ),
    .B(\u_cpu.REG_FILE._01050_ ),
    .X(\u_cpu.REG_FILE._01692_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06369_  (.A1(\u_cpu.REG_FILE._01475_ ),
    .A2(\u_cpu.REG_FILE.rf[8][10] ),
    .B1_N(\u_cpu.REG_FILE._01055_ ),
    .Y(\u_cpu.REG_FILE._01693_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06370_  (.A(\u_cpu.REG_FILE.rf[11][10] ),
    .B_N(\u_cpu.REG_FILE._01590_ ),
    .X(\u_cpu.REG_FILE._01694_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06371_  (.A1(\u_cpu.REG_FILE._01425_ ),
    .A2(\u_cpu.REG_FILE.rf[10][10] ),
    .B1(\u_cpu.REG_FILE._01360_ ),
    .C1(\u_cpu.REG_FILE._01694_ ),
    .Y(\u_cpu.REG_FILE._01695_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06372_  (.A1(\u_cpu.REG_FILE._01692_ ),
    .A2(\u_cpu.REG_FILE._01693_ ),
    .B1(\u_cpu.REG_FILE._01424_ ),
    .C1(\u_cpu.REG_FILE._01695_ ),
    .Y(\u_cpu.REG_FILE._01696_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06373_  (.A(\u_cpu.REG_FILE._01691_ ),
    .B(\u_cpu.REG_FILE._01696_ ),
    .C(\u_cpu.REG_FILE._01070_ ),
    .Y(\u_cpu.REG_FILE._01697_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06374_  (.A(\u_cpu.REG_FILE.rf[5][10] ),
    .Y(\u_cpu.REG_FILE._01698_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06375_  (.A1(\u_cpu.REG_FILE._01431_ ),
    .A2(\u_cpu.REG_FILE.rf[4][10] ),
    .B1_N(\u_cpu.REG_FILE._01482_ ),
    .Y(\u_cpu.REG_FILE._01699_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._06376_  (.A1(\u_cpu.REG_FILE._01698_ ),
    .A2(\u_cpu.REG_FILE._01075_ ),
    .B1(\u_cpu.REG_FILE._01699_ ),
    .Y(\u_cpu.REG_FILE._01700_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06377_  (.A1(\u_cpu.REG_FILE._01434_ ),
    .A2(\u_cpu.REG_FILE.rf[6][10] ),
    .B1(\u_cpu.REG_FILE._01598_ ),
    .Y(\u_cpu.REG_FILE._01701_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06378_  (.A_N(\u_cpu.REG_FILE.rf[7][10] ),
    .B(\u_cpu.REG_FILE._01085_ ),
    .X(\u_cpu.REG_FILE._01702_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06379_  (.A1(\u_cpu.REG_FILE._01701_ ),
    .A2(\u_cpu.REG_FILE._01702_ ),
    .B1(\u_cpu.REG_FILE._01601_ ),
    .Y(\u_cpu.REG_FILE._01703_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06380_  (.A_N(\u_cpu.REG_FILE.rf[1][10] ),
    .B(\u_cpu.REG_FILE._01091_ ),
    .X(\u_cpu.REG_FILE._01704_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06381_  (.A(\u_cpu.REG_FILE._01054_ ),
    .X(\u_cpu.REG_FILE._01705_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06382_  (.A1(\u_cpu.REG_FILE._01372_ ),
    .A2(\u_cpu.REG_FILE.rf[0][10] ),
    .B1_N(\u_cpu.REG_FILE._01705_ ),
    .Y(\u_cpu.REG_FILE._01706_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06383_  (.A(\u_cpu.REG_FILE._01052_ ),
    .X(\u_cpu.REG_FILE._01707_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06384_  (.A(\u_cpu.REG_FILE.rf[3][10] ),
    .B_N(\u_cpu.REG_FILE._01241_ ),
    .X(\u_cpu.REG_FILE._01708_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06385_  (.A1(\u_cpu.REG_FILE._01707_ ),
    .A2(\u_cpu.REG_FILE.rf[2][10] ),
    .B1(\u_cpu.REG_FILE._01240_ ),
    .C1(\u_cpu.REG_FILE._01708_ ),
    .Y(\u_cpu.REG_FILE._01709_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06386_  (.A1(\u_cpu.REG_FILE._01704_ ),
    .A2(\u_cpu.REG_FILE._01706_ ),
    .B1(\u_cpu.REG_FILE._01096_ ),
    .C1(\u_cpu.REG_FILE._01709_ ),
    .Y(\u_cpu.REG_FILE._01710_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06387_  (.A1(\u_cpu.REG_FILE._01700_ ),
    .A2(\u_cpu.REG_FILE._01703_ ),
    .B1(\u_cpu.REG_FILE._01603_ ),
    .C1(\u_cpu.REG_FILE._01710_ ),
    .Y(\u_cpu.REG_FILE._01711_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._06388_  (.A(\u_cpu.REG_FILE._01697_ ),
    .B(\u_cpu.REG_FILE._01711_ ),
    .Y(\u_cpu.REG_FILE._01712_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06389_  (.A(\u_cpu.REG_FILE.rf[27][10] ),
    .B_N(\u_cpu.REG_FILE._01108_ ),
    .X(\u_cpu.REG_FILE._01713_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06390_  (.A1(\u_cpu.REG_FILE._01105_ ),
    .A2(\u_cpu.REG_FILE.rf[26][10] ),
    .B1(\u_cpu.REG_FILE._01660_ ),
    .C1(\u_cpu.REG_FILE._01713_ ),
    .X(\u_cpu.REG_FILE._01714_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06391_  (.A1(\u_cpu.REG_FILE._01447_ ),
    .A2(\u_cpu.REG_FILE.rf[24][10] ),
    .B1_N(\u_cpu.REG_FILE._01062_ ),
    .X(\u_cpu.REG_FILE._01715_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06392_  (.A(\u_cpu.REG_FILE.rf[25][10] ),
    .B_N(\u_cpu.REG_FILE._01194_ ),
    .X(\u_cpu.REG_FILE._01716_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._06393_  (.A1(\u_cpu.REG_FILE._01715_ ),
    .A2(\u_cpu.REG_FILE._01716_ ),
    .B1(\u_cpu.REG_FILE._01196_ ),
    .X(\u_cpu.REG_FILE._01717_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06394_  (.A(\u_cpu.REG_FILE._01390_ ),
    .B(\u_cpu.REG_FILE.rf[30][10] ),
    .Y(\u_cpu.REG_FILE._01718_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06395_  (.A1(\u_cpu.REG_FILE.rf[31][10] ),
    .A2(\u_cpu.REG_FILE._01200_ ),
    .B1(\u_cpu.REG_FILE._01501_ ),
    .Y(\u_cpu.REG_FILE._01719_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06396_  (.A1(\u_cpu.REG_FILE._01503_ ),
    .A2(\u_cpu.REG_FILE.rf[28][10] ),
    .B1_N(\u_cpu.REG_FILE._01126_ ),
    .X(\u_cpu.REG_FILE._01720_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06397_  (.A1(\u_cpu.REG_FILE._01668_ ),
    .A2(\u_cpu.REG_FILE.rf[29][10] ),
    .B1(\u_cpu.REG_FILE._01720_ ),
    .Y(\u_cpu.REG_FILE._01721_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06398_  (.A1(\u_cpu.REG_FILE._01718_ ),
    .A2(\u_cpu.REG_FILE._01719_ ),
    .B1(\u_cpu.REG_FILE._01721_ ),
    .C1(\u_cpu.REG_FILE._01395_ ),
    .Y(\u_cpu.REG_FILE._01722_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06399_  (.A1(\u_cpu.REG_FILE._01714_ ),
    .A2(\u_cpu.REG_FILE._01717_ ),
    .B1(\u_cpu.REG_FILE._01198_ ),
    .C1(\u_cpu.REG_FILE._01722_ ),
    .Y(\u_cpu.REG_FILE._01723_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06400_  (.A1(\u_cpu.REG_FILE._01206_ ),
    .A2(\u_cpu.REG_FILE.rf[18][10] ),
    .B1(\u_cpu.REG_FILE._01135_ ),
    .Y(\u_cpu.REG_FILE._01724_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06401_  (.A(\u_cpu.REG_FILE.rf[19][10] ),
    .B(\u_cpu.REG_FILE._01509_ ),
    .Y(\u_cpu.REG_FILE._01725_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06402_  (.A(\u_cpu.REG_FILE._01123_ ),
    .X(\u_cpu.REG_FILE._01726_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06403_  (.A1(\u_cpu.REG_FILE._01141_ ),
    .A2(\u_cpu.REG_FILE.rf[16][10] ),
    .B1_N(\u_cpu.REG_FILE._01142_ ),
    .X(\u_cpu.REG_FILE._01727_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06404_  (.A1(\u_cpu.REG_FILE._01726_ ),
    .A2(\u_cpu.REG_FILE.rf[17][10] ),
    .B1(\u_cpu.REG_FILE._01727_ ),
    .Y(\u_cpu.REG_FILE._01728_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06405_  (.A1(\u_cpu.REG_FILE._01724_ ),
    .A2(\u_cpu.REG_FILE._01725_ ),
    .B1(\u_cpu.REG_FILE._01139_ ),
    .C1(\u_cpu.REG_FILE._01728_ ),
    .Y(\u_cpu.REG_FILE._01729_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06406_  (.A(\u_cpu.REG_FILE._01269_ ),
    .B(\u_cpu.REG_FILE.rf[22][10] ),
    .X(\u_cpu.REG_FILE._01730_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06407_  (.A1(\u_cpu.REG_FILE._01146_ ),
    .A2(\u_cpu.REG_FILE.rf[23][10] ),
    .B1(\u_cpu.REG_FILE._01147_ ),
    .C1(\u_cpu.REG_FILE._01730_ ),
    .Y(\u_cpu.REG_FILE._01731_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06408_  (.A1(\u_cpu.REG_FILE._01632_ ),
    .A2(\u_cpu.REG_FILE.rf[20][10] ),
    .B1_N(\u_cpu.REG_FILE._01214_ ),
    .X(\u_cpu.REG_FILE._01732_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06409_  (.A1(\u_cpu.REG_FILE._01151_ ),
    .A2(\u_cpu.REG_FILE.rf[21][10] ),
    .B1(\u_cpu.REG_FILE._01732_ ),
    .Y(\u_cpu.REG_FILE._01733_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06410_  (.A(\u_cpu.REG_FILE._01731_ ),
    .B(\u_cpu.REG_FILE._01733_ ),
    .C(\u_cpu.REG_FILE._01552_ ),
    .Y(\u_cpu.REG_FILE._01734_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06411_  (.A(\u_cpu.REG_FILE._01569_ ),
    .B(\u_cpu.REG_FILE._01729_ ),
    .C(\u_cpu.REG_FILE._01734_ ),
    .Y(\u_cpu.REG_FILE._01735_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06412_  (.A(\u_cpu.REG_FILE._01723_ ),
    .B(\u_cpu.REG_FILE._01735_ ),
    .C(\u_cpu.REG_FILE._01684_ ),
    .Y(\u_cpu.REG_FILE._01736_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06413_  (.A(\u_cpu.REG_FILE._01164_ ),
    .X(\u_cpu.REG_FILE._01737_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06414_  (.A1(\u_cpu.REG_FILE._01026_ ),
    .A2(\u_cpu.REG_FILE._01712_ ),
    .B1(\u_cpu.REG_FILE._01736_ ),
    .C1(\u_cpu.REG_FILE._01737_ ),
    .X(\u_cpu.ALU.SrcA[10] ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06415_  (.A1(\u_cpu.REG_FILE._01523_ ),
    .A2(\u_cpu.REG_FILE.rf[16][11] ),
    .B1_N(\u_cpu.REG_FILE._01032_ ),
    .Y(\u_cpu.REG_FILE._01738_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06416_  (.A_N(\u_cpu.REG_FILE.rf[17][11] ),
    .B(\u_cpu.REG_FILE._01111_ ),
    .X(\u_cpu.REG_FILE._01739_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06417_  (.A1(\u_cpu.REG_FILE._01260_ ),
    .A2(\u_cpu.REG_FILE.rf[18][11] ),
    .B1(\u_cpu.REG_FILE._01407_ ),
    .Y(\u_cpu.REG_FILE._01740_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06418_  (.A_N(\u_cpu.REG_FILE.rf[19][11] ),
    .B(\u_cpu.REG_FILE._01074_ ),
    .X(\u_cpu.REG_FILE._01741_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.REG_FILE._06419_  (.A1(\u_cpu.REG_FILE._01738_ ),
    .A2(\u_cpu.REG_FILE._01739_ ),
    .B1(\u_cpu.REG_FILE._01740_ ),
    .B2(\u_cpu.REG_FILE._01741_ ),
    .Y(\u_cpu.REG_FILE._01742_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06420_  (.A(\u_cpu.REG_FILE.rf[23][11] ),
    .B_N(\u_cpu.REG_FILE._01125_ ),
    .X(\u_cpu.REG_FILE._01743_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06421_  (.A1(\u_cpu.REG_FILE._01118_ ),
    .A2(\u_cpu.REG_FILE.rf[22][11] ),
    .B1(\u_cpu.REG_FILE._01121_ ),
    .C1(\u_cpu.REG_FILE._01743_ ),
    .X(\u_cpu.REG_FILE._01744_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06422_  (.A(\u_cpu.REG_FILE._01184_ ),
    .B(\u_cpu.REG_FILE.rf[20][11] ),
    .Y(\u_cpu.REG_FILE._01745_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06423_  (.A_N(\u_cpu.REG_FILE.rf[21][11] ),
    .B(\u_cpu.REG_FILE._01161_ ),
    .X(\u_cpu.REG_FILE._01746_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.REG_FILE._06424_  (.A1(\u_cpu.REG_FILE._01259_ ),
    .A2(\u_cpu.REG_FILE._01745_ ),
    .A3(\u_cpu.REG_FILE._01746_ ),
    .B1(\u_cpu.REG_FILE._01087_ ),
    .Y(\u_cpu.REG_FILE._01747_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.REG_FILE._06425_  (.A1(\u_cpu.REG_FILE._01277_ ),
    .A2(\u_cpu.REG_FILE._01742_ ),
    .B1(\u_cpu.REG_FILE._01744_ ),
    .B2(\u_cpu.REG_FILE._01747_ ),
    .C1(\u_cpu.REG_FILE._01132_ ),
    .X(\u_cpu.REG_FILE._01748_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06426_  (.A(\u_cpu.REG_FILE._01549_ ),
    .B(\u_cpu.REG_FILE.rf[28][11] ),
    .Y(\u_cpu.REG_FILE._01749_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06427_  (.A(\u_cpu.REG_FILE._01073_ ),
    .X(\u_cpu.REG_FILE._01750_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06428_  (.A_N(\u_cpu.REG_FILE.rf[29][11] ),
    .B(\u_cpu.REG_FILE._01750_ ),
    .X(\u_cpu.REG_FILE._01751_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06429_  (.A(\u_cpu.REG_FILE.rf[31][11] ),
    .B_N(\u_cpu.REG_FILE._01060_ ),
    .X(\u_cpu.REG_FILE._01752_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06430_  (.A1(\u_cpu.REG_FILE._01325_ ),
    .A2(\u_cpu.REG_FILE.rf[30][11] ),
    .B1(\u_cpu.REG_FILE._01280_ ),
    .C1(\u_cpu.REG_FILE._01752_ ),
    .Y(\u_cpu.REG_FILE._01753_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._06431_  (.A1(\u_cpu.REG_FILE._01259_ ),
    .A2(\u_cpu.REG_FILE._01749_ ),
    .A3(\u_cpu.REG_FILE._01751_ ),
    .B1(\u_cpu.REG_FILE._01087_ ),
    .C1(\u_cpu.REG_FILE._01753_ ),
    .Y(\u_cpu.REG_FILE._01754_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06432_  (.A_N(\u_cpu.REG_FILE.rf[25][11] ),
    .B(\u_cpu.REG_FILE._01074_ ),
    .X(\u_cpu.REG_FILE._01755_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06433_  (.A1(\u_cpu.REG_FILE._01093_ ),
    .A2(\u_cpu.REG_FILE.rf[24][11] ),
    .B1_N(\u_cpu.REG_FILE._01550_ ),
    .Y(\u_cpu.REG_FILE._01756_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06434_  (.A(\u_cpu.REG_FILE.rf[27][11] ),
    .B_N(\u_cpu.REG_FILE._01310_ ),
    .X(\u_cpu.REG_FILE._01757_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06435_  (.A1(\u_cpu.REG_FILE._01308_ ),
    .A2(\u_cpu.REG_FILE.rf[26][11] ),
    .B1(\u_cpu.REG_FILE._01309_ ),
    .C1(\u_cpu.REG_FILE._01757_ ),
    .Y(\u_cpu.REG_FILE._01758_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06436_  (.A1(\u_cpu.REG_FILE._01755_ ),
    .A2(\u_cpu.REG_FILE._01756_ ),
    .B1(\u_cpu.REG_FILE._01307_ ),
    .C1(\u_cpu.REG_FILE._01758_ ),
    .Y(\u_cpu.REG_FILE._01759_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._06437_  (.A1(\u_cpu.REG_FILE._01754_ ),
    .A2(\u_cpu.REG_FILE._01759_ ),
    .A3(\u_cpu.REG_FILE._01314_ ),
    .B1(\u_cpu.REG_FILE._01315_ ),
    .X(\u_cpu.REG_FILE._01760_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06438_  (.A1(\u_cpu.REG_FILE._01317_ ),
    .A2(\u_cpu.REG_FILE.rf[8][11] ),
    .B1_N(\u_cpu.REG_FILE._01032_ ),
    .Y(\u_cpu.REG_FILE._01761_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06439_  (.A_N(\u_cpu.REG_FILE.rf[9][11] ),
    .B(\u_cpu.REG_FILE._01041_ ),
    .X(\u_cpu.REG_FILE._01762_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06440_  (.A1(\u_cpu.REG_FILE._01761_ ),
    .A2(\u_cpu.REG_FILE._01762_ ),
    .B1(\u_cpu.REG_FILE._01264_ ),
    .Y(\u_cpu.REG_FILE._01763_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06441_  (.A(\u_cpu.REG_FILE._01148_ ),
    .B(\u_cpu.REG_FILE.rf[10][11] ),
    .X(\u_cpu.REG_FILE._01764_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06442_  (.A1(\u_cpu.REG_FILE._01321_ ),
    .A2(\u_cpu.REG_FILE.rf[11][11] ),
    .B1(\u_cpu.REG_FILE._01280_ ),
    .C1(\u_cpu.REG_FILE._01764_ ),
    .X(\u_cpu.REG_FILE._01765_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06443_  (.A(\u_cpu.REG_FILE._01325_ ),
    .B(\u_cpu.REG_FILE.rf[14][11] ),
    .Y(\u_cpu.REG_FILE._01766_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06444_  (.A1(\u_cpu.REG_FILE.rf[15][11] ),
    .A2(\u_cpu.REG_FILE._01327_ ),
    .B1(\u_cpu.REG_FILE._01099_ ),
    .Y(\u_cpu.REG_FILE._01767_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06445_  (.A1(\u_cpu.REG_FILE._01330_ ),
    .A2(\u_cpu.REG_FILE.rf[12][11] ),
    .B1_N(\u_cpu.REG_FILE._01082_ ),
    .X(\u_cpu.REG_FILE._01768_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06446_  (.A1(\u_cpu.REG_FILE._01329_ ),
    .A2(\u_cpu.REG_FILE.rf[13][11] ),
    .B1(\u_cpu.REG_FILE._01768_ ),
    .Y(\u_cpu.REG_FILE._01769_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06447_  (.A1(\u_cpu.REG_FILE._01766_ ),
    .A2(\u_cpu.REG_FILE._01767_ ),
    .B1(\u_cpu.REG_FILE._01769_ ),
    .C1(\u_cpu.REG_FILE._01333_ ),
    .Y(\u_cpu.REG_FILE._01770_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06448_  (.A1(\u_cpu.REG_FILE._01763_ ),
    .A2(\u_cpu.REG_FILE._01765_ ),
    .B1(\u_cpu.REG_FILE._01069_ ),
    .C1(\u_cpu.REG_FILE._01770_ ),
    .Y(\u_cpu.REG_FILE._01771_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06449_  (.A1(\u_cpu.REG_FILE._01523_ ),
    .A2(\u_cpu.REG_FILE.rf[6][11] ),
    .B1(\u_cpu.REG_FILE._01533_ ),
    .Y(\u_cpu.REG_FILE._01772_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06450_  (.A_N(\u_cpu.REG_FILE.rf[7][11] ),
    .B(\u_cpu.REG_FILE._01029_ ),
    .X(\u_cpu.REG_FILE._01773_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06451_  (.A(\u_cpu.REG_FILE._01049_ ),
    .X(\u_cpu.REG_FILE._01774_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06452_  (.A1(\u_cpu.REG_FILE._01774_ ),
    .A2(\u_cpu.REG_FILE.rf[4][11] ),
    .B1_N(\u_cpu.REG_FILE._01553_ ),
    .Y(\u_cpu.REG_FILE._01775_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06453_  (.A_N(\u_cpu.REG_FILE.rf[5][11] ),
    .B(\u_cpu.REG_FILE._01382_ ),
    .X(\u_cpu.REG_FILE._01776_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.REG_FILE._06454_  (.A1(\u_cpu.REG_FILE._01772_ ),
    .A2(\u_cpu.REG_FILE._01773_ ),
    .B1(\u_cpu.REG_FILE._01775_ ),
    .B2(\u_cpu.REG_FILE._01776_ ),
    .Y(\u_cpu.REG_FILE._01777_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06455_  (.A(\u_cpu.REG_FILE._01317_ ),
    .B(\u_cpu.REG_FILE.rf[0][11] ),
    .Y(\u_cpu.REG_FILE._01778_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06456_  (.A_N(\u_cpu.REG_FILE.rf[1][11] ),
    .B(\u_cpu.REG_FILE._01125_ ),
    .X(\u_cpu.REG_FILE._01779_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06457_  (.A(\u_cpu.REG_FILE.rf[3][11] ),
    .B_N(\u_cpu.REG_FILE._01076_ ),
    .X(\u_cpu.REG_FILE._01780_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06458_  (.A1(\u_cpu.REG_FILE._01404_ ),
    .A2(\u_cpu.REG_FILE.rf[2][11] ),
    .B1(\u_cpu.REG_FILE._01533_ ),
    .C1(\u_cpu.REG_FILE._01780_ ),
    .Y(\u_cpu.REG_FILE._01781_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._06459_  (.A1(\u_cpu.REG_FILE._01527_ ),
    .A2(\u_cpu.REG_FILE._01778_ ),
    .A3(\u_cpu.REG_FILE._01779_ ),
    .B1(\u_cpu.REG_FILE._01058_ ),
    .C1(\u_cpu.REG_FILE._01781_ ),
    .Y(\u_cpu.REG_FILE._01782_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06460_  (.A1(\u_cpu.REG_FILE._01525_ ),
    .A2(\u_cpu.REG_FILE._01777_ ),
    .B1(\u_cpu.REG_FILE._01782_ ),
    .C1(\u_cpu.REG_FILE._01541_ ),
    .Y(\u_cpu.REG_FILE._01783_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06461_  (.A(\u_cpu.REG_FILE._01315_ ),
    .B(\u_cpu.REG_FILE._01771_ ),
    .C(\u_cpu.REG_FILE._01783_ ),
    .Y(\u_cpu.REG_FILE._01784_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06462_  (.A1(\u_cpu.REG_FILE._01748_ ),
    .A2(\u_cpu.REG_FILE._01760_ ),
    .B1(\u_cpu.REG_FILE._01784_ ),
    .C1(\u_cpu.REG_FILE._01737_ ),
    .X(\u_cpu.ALU.SrcA[11] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06463_  (.A(\u_cpu.REG_FILE.rf[15][12] ),
    .B_N(\u_cpu.REG_FILE._01034_ ),
    .X(\u_cpu.REG_FILE._01785_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06464_  (.A1(\u_cpu.REG_FILE._01351_ ),
    .A2(\u_cpu.REG_FILE.rf[14][12] ),
    .B1(\u_cpu.REG_FILE._01352_ ),
    .C1(\u_cpu.REG_FILE._01785_ ),
    .Y(\u_cpu.REG_FILE._01786_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06465_  (.A(\u_cpu.REG_FILE._01038_ ),
    .X(\u_cpu.REG_FILE._01787_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06466_  (.A1(\u_cpu.REG_FILE._01584_ ),
    .A2(\u_cpu.REG_FILE.rf[12][12] ),
    .B1_N(\u_cpu.REG_FILE._01042_ ),
    .X(\u_cpu.REG_FILE._01788_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06467_  (.A1(\u_cpu.REG_FILE._01787_ ),
    .A2(\u_cpu.REG_FILE.rf[13][12] ),
    .B1(\u_cpu.REG_FILE._01788_ ),
    .Y(\u_cpu.REG_FILE._01789_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06468_  (.A(\u_cpu.REG_FILE._01786_ ),
    .B(\u_cpu.REG_FILE._01789_ ),
    .C(\u_cpu.REG_FILE._01690_ ),
    .Y(\u_cpu.REG_FILE._01790_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06469_  (.A_N(\u_cpu.REG_FILE.rf[9][12] ),
    .B(\u_cpu.REG_FILE._01050_ ),
    .X(\u_cpu.REG_FILE._01791_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06470_  (.A1(\u_cpu.REG_FILE._01475_ ),
    .A2(\u_cpu.REG_FILE.rf[8][12] ),
    .B1_N(\u_cpu.REG_FILE._01055_ ),
    .Y(\u_cpu.REG_FILE._01792_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06471_  (.A(\u_cpu.REG_FILE.rf[11][12] ),
    .B_N(\u_cpu.REG_FILE._01590_ ),
    .X(\u_cpu.REG_FILE._01793_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06472_  (.A1(\u_cpu.REG_FILE._01425_ ),
    .A2(\u_cpu.REG_FILE.rf[10][12] ),
    .B1(\u_cpu.REG_FILE._01360_ ),
    .C1(\u_cpu.REG_FILE._01793_ ),
    .Y(\u_cpu.REG_FILE._01794_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06473_  (.A1(\u_cpu.REG_FILE._01791_ ),
    .A2(\u_cpu.REG_FILE._01792_ ),
    .B1(\u_cpu.REG_FILE._01424_ ),
    .C1(\u_cpu.REG_FILE._01794_ ),
    .Y(\u_cpu.REG_FILE._01795_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06474_  (.A(\u_cpu.REG_FILE._01069_ ),
    .X(\u_cpu.REG_FILE._01796_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06475_  (.A(\u_cpu.REG_FILE._01790_ ),
    .B(\u_cpu.REG_FILE._01795_ ),
    .C(\u_cpu.REG_FILE._01796_ ),
    .Y(\u_cpu.REG_FILE._01797_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06476_  (.A(\u_cpu.REG_FILE.rf[5][12] ),
    .Y(\u_cpu.REG_FILE._01798_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06477_  (.A1(\u_cpu.REG_FILE._01431_ ),
    .A2(\u_cpu.REG_FILE.rf[4][12] ),
    .B1_N(\u_cpu.REG_FILE._01482_ ),
    .Y(\u_cpu.REG_FILE._01799_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._06478_  (.A1(\u_cpu.REG_FILE._01798_ ),
    .A2(\u_cpu.REG_FILE._01075_ ),
    .B1(\u_cpu.REG_FILE._01799_ ),
    .Y(\u_cpu.REG_FILE._01800_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06479_  (.A1(\u_cpu.REG_FILE._01434_ ),
    .A2(\u_cpu.REG_FILE.rf[6][12] ),
    .B1(\u_cpu.REG_FILE._01598_ ),
    .Y(\u_cpu.REG_FILE._01801_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06480_  (.A_N(\u_cpu.REG_FILE.rf[7][12] ),
    .B(\u_cpu.REG_FILE._01085_ ),
    .X(\u_cpu.REG_FILE._01802_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06481_  (.A1(\u_cpu.REG_FILE._01801_ ),
    .A2(\u_cpu.REG_FILE._01802_ ),
    .B1(\u_cpu.REG_FILE._01601_ ),
    .Y(\u_cpu.REG_FILE._01803_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06482_  (.A(\u_cpu.REG_FILE._01073_ ),
    .X(\u_cpu.REG_FILE._01804_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06483_  (.A_N(\u_cpu.REG_FILE.rf[1][12] ),
    .B(\u_cpu.REG_FILE._01804_ ),
    .X(\u_cpu.REG_FILE._01805_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06484_  (.A1(\u_cpu.REG_FILE._01372_ ),
    .A2(\u_cpu.REG_FILE.rf[0][12] ),
    .B1_N(\u_cpu.REG_FILE._01705_ ),
    .Y(\u_cpu.REG_FILE._01806_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06485_  (.A(\u_cpu.REG_FILE.rf[3][12] ),
    .B_N(\u_cpu.REG_FILE._01241_ ),
    .X(\u_cpu.REG_FILE._01807_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06486_  (.A1(\u_cpu.REG_FILE._01707_ ),
    .A2(\u_cpu.REG_FILE.rf[2][12] ),
    .B1(\u_cpu.REG_FILE._01240_ ),
    .C1(\u_cpu.REG_FILE._01807_ ),
    .Y(\u_cpu.REG_FILE._01808_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06487_  (.A1(\u_cpu.REG_FILE._01805_ ),
    .A2(\u_cpu.REG_FILE._01806_ ),
    .B1(\u_cpu.REG_FILE._01096_ ),
    .C1(\u_cpu.REG_FILE._01808_ ),
    .Y(\u_cpu.REG_FILE._01809_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06488_  (.A1(\u_cpu.REG_FILE._01800_ ),
    .A2(\u_cpu.REG_FILE._01803_ ),
    .B1(\u_cpu.REG_FILE._01603_ ),
    .C1(\u_cpu.REG_FILE._01809_ ),
    .Y(\u_cpu.REG_FILE._01810_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._06489_  (.A(\u_cpu.REG_FILE._01797_ ),
    .B(\u_cpu.REG_FILE._01810_ ),
    .Y(\u_cpu.REG_FILE._01811_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06490_  (.A1(\u_cpu.REG_FILE._01379_ ),
    .A2(\u_cpu.REG_FILE.rf[24][12] ),
    .B1_N(\u_cpu.REG_FILE._01611_ ),
    .Y(\u_cpu.REG_FILE._01812_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06491_  (.A_N(\u_cpu.REG_FILE.rf[25][12] ),
    .B(\u_cpu.REG_FILE._01382_ ),
    .X(\u_cpu.REG_FILE._01813_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06492_  (.A(\u_cpu.REG_FILE._01058_ ),
    .X(\u_cpu.REG_FILE._01814_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06493_  (.A1(\u_cpu.REG_FILE._01812_ ),
    .A2(\u_cpu.REG_FILE._01813_ ),
    .B1(\u_cpu.REG_FILE._01814_ ),
    .Y(\u_cpu.REG_FILE._01815_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06494_  (.A(\u_cpu.REG_FILE._01340_ ),
    .B(\u_cpu.REG_FILE.rf[26][12] ),
    .X(\u_cpu.REG_FILE._01816_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06495_  (.A1(\u_cpu.REG_FILE._01386_ ),
    .A2(\u_cpu.REG_FILE.rf[27][12] ),
    .B1(\u_cpu.REG_FILE._01387_ ),
    .C1(\u_cpu.REG_FILE._01816_ ),
    .X(\u_cpu.REG_FILE._01817_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06496_  (.A(\u_cpu.REG_FILE._01097_ ),
    .B(\u_cpu.REG_FILE.rf[30][12] ),
    .Y(\u_cpu.REG_FILE._01818_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06497_  (.A1(\u_cpu.REG_FILE.rf[31][12] ),
    .A2(\u_cpu.REG_FILE._01327_ ),
    .B1(\u_cpu.REG_FILE._01618_ ),
    .Y(\u_cpu.REG_FILE._01819_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06498_  (.A(\u_cpu.REG_FILE._01325_ ),
    .B(\u_cpu.REG_FILE.rf[28][12] ),
    .Y(\u_cpu.REG_FILE._01820_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06499_  (.A1(\u_cpu.REG_FILE.rf[29][12] ),
    .A2(\u_cpu.REG_FILE._01265_ ),
    .B1_N(\u_cpu.REG_FILE._01521_ ),
    .Y(\u_cpu.REG_FILE._01821_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._06500_  (.A1(\u_cpu.REG_FILE._01818_ ),
    .A2(\u_cpu.REG_FILE._01819_ ),
    .B1(\u_cpu.REG_FILE._01820_ ),
    .B2(\u_cpu.REG_FILE._01821_ ),
    .C1(\u_cpu.REG_FILE._01333_ ),
    .Y(\u_cpu.REG_FILE._01822_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06501_  (.A1(\u_cpu.REG_FILE._01815_ ),
    .A2(\u_cpu.REG_FILE._01817_ ),
    .B1(\u_cpu.REG_FILE._01198_ ),
    .C1(\u_cpu.REG_FILE._01822_ ),
    .Y(\u_cpu.REG_FILE._01823_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06502_  (.A1(\u_cpu.REG_FILE._01206_ ),
    .A2(\u_cpu.REG_FILE.rf[18][12] ),
    .B1(\u_cpu.REG_FILE._01135_ ),
    .Y(\u_cpu.REG_FILE._01824_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06503_  (.A(\u_cpu.REG_FILE.rf[19][12] ),
    .B(\u_cpu.REG_FILE._01509_ ),
    .Y(\u_cpu.REG_FILE._01825_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06504_  (.A1(\u_cpu.REG_FILE._01141_ ),
    .A2(\u_cpu.REG_FILE.rf[16][12] ),
    .B1_N(\u_cpu.REG_FILE._01153_ ),
    .X(\u_cpu.REG_FILE._01826_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06505_  (.A1(\u_cpu.REG_FILE._01726_ ),
    .A2(\u_cpu.REG_FILE.rf[17][12] ),
    .B1(\u_cpu.REG_FILE._01826_ ),
    .Y(\u_cpu.REG_FILE._01827_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06506_  (.A1(\u_cpu.REG_FILE._01824_ ),
    .A2(\u_cpu.REG_FILE._01825_ ),
    .B1(\u_cpu.REG_FILE._01139_ ),
    .C1(\u_cpu.REG_FILE._01827_ ),
    .Y(\u_cpu.REG_FILE._01828_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06507_  (.A(\u_cpu.REG_FILE._01269_ ),
    .B(\u_cpu.REG_FILE.rf[22][12] ),
    .X(\u_cpu.REG_FILE._01829_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06508_  (.A1(\u_cpu.REG_FILE._01321_ ),
    .A2(\u_cpu.REG_FILE.rf[23][12] ),
    .B1(\u_cpu.REG_FILE._01063_ ),
    .C1(\u_cpu.REG_FILE._01829_ ),
    .Y(\u_cpu.REG_FILE._01830_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06509_  (.A1(\u_cpu.REG_FILE._01632_ ),
    .A2(\u_cpu.REG_FILE.rf[20][12] ),
    .B1_N(\u_cpu.REG_FILE._01214_ ),
    .X(\u_cpu.REG_FILE._01831_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06510_  (.A1(\u_cpu.REG_FILE._01151_ ),
    .A2(\u_cpu.REG_FILE.rf[21][12] ),
    .B1(\u_cpu.REG_FILE._01831_ ),
    .Y(\u_cpu.REG_FILE._01832_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06511_  (.A(\u_cpu.REG_FILE._01830_ ),
    .B(\u_cpu.REG_FILE._01832_ ),
    .C(\u_cpu.REG_FILE._01552_ ),
    .Y(\u_cpu.REG_FILE._01833_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06512_  (.A(\u_cpu.REG_FILE._01569_ ),
    .B(\u_cpu.REG_FILE._01828_ ),
    .C(\u_cpu.REG_FILE._01833_ ),
    .Y(\u_cpu.REG_FILE._01834_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06513_  (.A(\u_cpu.REG_FILE._01823_ ),
    .B(\u_cpu.REG_FILE._01834_ ),
    .C(\u_cpu.REG_FILE._01684_ ),
    .Y(\u_cpu.REG_FILE._01835_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06514_  (.A1(\u_cpu.REG_FILE._01026_ ),
    .A2(\u_cpu.REG_FILE._01811_ ),
    .B1(\u_cpu.REG_FILE._01835_ ),
    .C1(\u_cpu.REG_FILE._01737_ ),
    .X(\u_cpu.ALU.SrcA[12] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06515_  (.A(\u_cpu.REG_FILE.rf[15][13] ),
    .B_N(\u_cpu.REG_FILE._01034_ ),
    .X(\u_cpu.REG_FILE._01836_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06516_  (.A1(\u_cpu.REG_FILE._01351_ ),
    .A2(\u_cpu.REG_FILE.rf[14][13] ),
    .B1(\u_cpu.REG_FILE._01352_ ),
    .C1(\u_cpu.REG_FILE._01836_ ),
    .Y(\u_cpu.REG_FILE._01837_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06517_  (.A(\u_cpu.REG_FILE._01031_ ),
    .X(\u_cpu.REG_FILE._01838_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06518_  (.A1(\u_cpu.REG_FILE._01584_ ),
    .A2(\u_cpu.REG_FILE.rf[12][13] ),
    .B1_N(\u_cpu.REG_FILE._01838_ ),
    .X(\u_cpu.REG_FILE._01839_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06519_  (.A1(\u_cpu.REG_FILE._01787_ ),
    .A2(\u_cpu.REG_FILE.rf[13][13] ),
    .B1(\u_cpu.REG_FILE._01839_ ),
    .Y(\u_cpu.REG_FILE._01840_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06520_  (.A(\u_cpu.REG_FILE._01837_ ),
    .B(\u_cpu.REG_FILE._01840_ ),
    .C(\u_cpu.REG_FILE._01690_ ),
    .Y(\u_cpu.REG_FILE._01841_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06521_  (.A_N(\u_cpu.REG_FILE.rf[9][13] ),
    .B(\u_cpu.REG_FILE._01050_ ),
    .X(\u_cpu.REG_FILE._01842_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06522_  (.A(\u_cpu.REG_FILE._01054_ ),
    .X(\u_cpu.REG_FILE._01843_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06523_  (.A1(\u_cpu.REG_FILE._01475_ ),
    .A2(\u_cpu.REG_FILE.rf[8][13] ),
    .B1_N(\u_cpu.REG_FILE._01843_ ),
    .Y(\u_cpu.REG_FILE._01844_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06524_  (.A(\u_cpu.REG_FILE.rf[11][13] ),
    .B_N(\u_cpu.REG_FILE._01590_ ),
    .X(\u_cpu.REG_FILE._01845_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06525_  (.A1(\u_cpu.REG_FILE._01425_ ),
    .A2(\u_cpu.REG_FILE.rf[10][13] ),
    .B1(\u_cpu.REG_FILE._01360_ ),
    .C1(\u_cpu.REG_FILE._01845_ ),
    .Y(\u_cpu.REG_FILE._01846_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06526_  (.A1(\u_cpu.REG_FILE._01842_ ),
    .A2(\u_cpu.REG_FILE._01844_ ),
    .B1(\u_cpu.REG_FILE._01424_ ),
    .C1(\u_cpu.REG_FILE._01846_ ),
    .Y(\u_cpu.REG_FILE._01847_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06527_  (.A(\u_cpu.REG_FILE._01841_ ),
    .B(\u_cpu.REG_FILE._01847_ ),
    .C(\u_cpu.REG_FILE._01796_ ),
    .Y(\u_cpu.REG_FILE._01848_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06528_  (.A(\u_cpu.REG_FILE.rf[5][13] ),
    .Y(\u_cpu.REG_FILE._01849_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06529_  (.A(\u_cpu.REG_FILE._01074_ ),
    .X(\u_cpu.REG_FILE._01850_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06530_  (.A1(\u_cpu.REG_FILE._01431_ ),
    .A2(\u_cpu.REG_FILE.rf[4][13] ),
    .B1_N(\u_cpu.REG_FILE._01482_ ),
    .Y(\u_cpu.REG_FILE._01851_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._06531_  (.A1(\u_cpu.REG_FILE._01849_ ),
    .A2(\u_cpu.REG_FILE._01850_ ),
    .B1(\u_cpu.REG_FILE._01851_ ),
    .Y(\u_cpu.REG_FILE._01852_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06532_  (.A1(\u_cpu.REG_FILE._01434_ ),
    .A2(\u_cpu.REG_FILE.rf[6][13] ),
    .B1(\u_cpu.REG_FILE._01598_ ),
    .Y(\u_cpu.REG_FILE._01853_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06533_  (.A_N(\u_cpu.REG_FILE.rf[7][13] ),
    .B(\u_cpu.REG_FILE._01085_ ),
    .X(\u_cpu.REG_FILE._01854_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06534_  (.A1(\u_cpu.REG_FILE._01853_ ),
    .A2(\u_cpu.REG_FILE._01854_ ),
    .B1(\u_cpu.REG_FILE._01601_ ),
    .Y(\u_cpu.REG_FILE._01855_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06535_  (.A_N(\u_cpu.REG_FILE.rf[1][13] ),
    .B(\u_cpu.REG_FILE._01804_ ),
    .X(\u_cpu.REG_FILE._01856_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06536_  (.A1(\u_cpu.REG_FILE._01372_ ),
    .A2(\u_cpu.REG_FILE.rf[0][13] ),
    .B1_N(\u_cpu.REG_FILE._01705_ ),
    .Y(\u_cpu.REG_FILE._01857_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06537_  (.A(\u_cpu.REG_FILE._01057_ ),
    .X(\u_cpu.REG_FILE._01858_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06538_  (.A(\u_cpu.REG_FILE.rf[3][13] ),
    .B_N(\u_cpu.REG_FILE._01241_ ),
    .X(\u_cpu.REG_FILE._01859_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06539_  (.A1(\u_cpu.REG_FILE._01707_ ),
    .A2(\u_cpu.REG_FILE.rf[2][13] ),
    .B1(\u_cpu.REG_FILE._01240_ ),
    .C1(\u_cpu.REG_FILE._01859_ ),
    .Y(\u_cpu.REG_FILE._01860_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06540_  (.A1(\u_cpu.REG_FILE._01856_ ),
    .A2(\u_cpu.REG_FILE._01857_ ),
    .B1(\u_cpu.REG_FILE._01858_ ),
    .C1(\u_cpu.REG_FILE._01860_ ),
    .Y(\u_cpu.REG_FILE._01861_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06541_  (.A1(\u_cpu.REG_FILE._01852_ ),
    .A2(\u_cpu.REG_FILE._01855_ ),
    .B1(\u_cpu.REG_FILE._01603_ ),
    .C1(\u_cpu.REG_FILE._01861_ ),
    .Y(\u_cpu.REG_FILE._01862_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._06542_  (.A(\u_cpu.REG_FILE._01848_ ),
    .B(\u_cpu.REG_FILE._01862_ ),
    .Y(\u_cpu.REG_FILE._01863_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06543_  (.A(\u_cpu.REG_FILE.rf[27][13] ),
    .B_N(\u_cpu.REG_FILE._01108_ ),
    .X(\u_cpu.REG_FILE._01864_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06544_  (.A1(\u_cpu.REG_FILE._01105_ ),
    .A2(\u_cpu.REG_FILE.rf[26][13] ),
    .B1(\u_cpu.REG_FILE._01660_ ),
    .C1(\u_cpu.REG_FILE._01864_ ),
    .X(\u_cpu.REG_FILE._01865_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06545_  (.A1(\u_cpu.REG_FILE._01447_ ),
    .A2(\u_cpu.REG_FILE.rf[24][13] ),
    .B1_N(\u_cpu.REG_FILE._01062_ ),
    .X(\u_cpu.REG_FILE._01866_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06546_  (.A(\u_cpu.REG_FILE.rf[25][13] ),
    .B_N(\u_cpu.REG_FILE._01194_ ),
    .X(\u_cpu.REG_FILE._01867_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._06547_  (.A1(\u_cpu.REG_FILE._01866_ ),
    .A2(\u_cpu.REG_FILE._01867_ ),
    .B1(\u_cpu.REG_FILE._01196_ ),
    .X(\u_cpu.REG_FILE._01868_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06548_  (.A(\u_cpu.M_AXI_WDATA[18] ),
    .X(\u_cpu.REG_FILE._01869_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06549_  (.A(\u_cpu.REG_FILE._01390_ ),
    .B(\u_cpu.REG_FILE.rf[30][13] ),
    .Y(\u_cpu.REG_FILE._01870_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06550_  (.A1(\u_cpu.REG_FILE.rf[31][13] ),
    .A2(\u_cpu.REG_FILE._01200_ ),
    .B1(\u_cpu.REG_FILE._01501_ ),
    .Y(\u_cpu.REG_FILE._01871_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06551_  (.A1(\u_cpu.REG_FILE._01503_ ),
    .A2(\u_cpu.REG_FILE.rf[28][13] ),
    .B1_N(\u_cpu.REG_FILE._01126_ ),
    .X(\u_cpu.REG_FILE._01872_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06552_  (.A1(\u_cpu.REG_FILE._01668_ ),
    .A2(\u_cpu.REG_FILE.rf[29][13] ),
    .B1(\u_cpu.REG_FILE._01872_ ),
    .Y(\u_cpu.REG_FILE._01873_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06553_  (.A1(\u_cpu.REG_FILE._01870_ ),
    .A2(\u_cpu.REG_FILE._01871_ ),
    .B1(\u_cpu.REG_FILE._01873_ ),
    .C1(\u_cpu.REG_FILE._01395_ ),
    .Y(\u_cpu.REG_FILE._01874_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06554_  (.A1(\u_cpu.REG_FILE._01865_ ),
    .A2(\u_cpu.REG_FILE._01868_ ),
    .B1(\u_cpu.REG_FILE._01869_ ),
    .C1(\u_cpu.REG_FILE._01874_ ),
    .Y(\u_cpu.REG_FILE._01875_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06555_  (.A1(\u_cpu.REG_FILE._01206_ ),
    .A2(\u_cpu.REG_FILE.rf[18][13] ),
    .B1(\u_cpu.REG_FILE._01135_ ),
    .Y(\u_cpu.REG_FILE._01876_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06556_  (.A(\u_cpu.REG_FILE.rf[19][13] ),
    .B(\u_cpu.REG_FILE._01509_ ),
    .Y(\u_cpu.REG_FILE._01877_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06557_  (.A1(\u_cpu.REG_FILE._01141_ ),
    .A2(\u_cpu.REG_FILE.rf[16][13] ),
    .B1_N(\u_cpu.REG_FILE._01153_ ),
    .X(\u_cpu.REG_FILE._01878_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06558_  (.A1(\u_cpu.REG_FILE._01726_ ),
    .A2(\u_cpu.REG_FILE.rf[17][13] ),
    .B1(\u_cpu.REG_FILE._01878_ ),
    .Y(\u_cpu.REG_FILE._01879_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06559_  (.A1(\u_cpu.REG_FILE._01876_ ),
    .A2(\u_cpu.REG_FILE._01877_ ),
    .B1(\u_cpu.REG_FILE._01264_ ),
    .C1(\u_cpu.REG_FILE._01879_ ),
    .Y(\u_cpu.REG_FILE._01880_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06560_  (.A(\u_cpu.REG_FILE._01269_ ),
    .B(\u_cpu.REG_FILE.rf[22][13] ),
    .X(\u_cpu.REG_FILE._01881_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06561_  (.A1(\u_cpu.REG_FILE._01321_ ),
    .A2(\u_cpu.REG_FILE.rf[23][13] ),
    .B1(\u_cpu.REG_FILE._01063_ ),
    .C1(\u_cpu.REG_FILE._01881_ ),
    .Y(\u_cpu.REG_FILE._01882_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06562_  (.A1(\u_cpu.REG_FILE._01632_ ),
    .A2(\u_cpu.REG_FILE.rf[20][13] ),
    .B1_N(\u_cpu.REG_FILE._01214_ ),
    .X(\u_cpu.REG_FILE._01883_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06563_  (.A1(\u_cpu.REG_FILE._01120_ ),
    .A2(\u_cpu.REG_FILE.rf[21][13] ),
    .B1(\u_cpu.REG_FILE._01883_ ),
    .Y(\u_cpu.REG_FILE._01884_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06564_  (.A(\u_cpu.REG_FILE._01882_ ),
    .B(\u_cpu.REG_FILE._01884_ ),
    .C(\u_cpu.REG_FILE._01552_ ),
    .Y(\u_cpu.REG_FILE._01885_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06565_  (.A(\u_cpu.REG_FILE._01569_ ),
    .B(\u_cpu.REG_FILE._01880_ ),
    .C(\u_cpu.REG_FILE._01885_ ),
    .Y(\u_cpu.REG_FILE._01886_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06566_  (.A(\u_cpu.REG_FILE._01875_ ),
    .B(\u_cpu.REG_FILE._01886_ ),
    .C(\u_cpu.REG_FILE._01684_ ),
    .Y(\u_cpu.REG_FILE._01887_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06567_  (.A1(\u_cpu.REG_FILE._01026_ ),
    .A2(\u_cpu.REG_FILE._01863_ ),
    .B1(\u_cpu.REG_FILE._01887_ ),
    .C1(\u_cpu.REG_FILE._01737_ ),
    .X(\u_cpu.ALU.SrcA[13] ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06568_  (.A(\u_cpu.REG_FILE._01024_ ),
    .X(\u_cpu.REG_FILE._01888_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06569_  (.A(\u_cpu.REG_FILE._01028_ ),
    .X(\u_cpu.REG_FILE._01889_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06570_  (.A(\u_cpu.REG_FILE.rf[15][14] ),
    .B_N(\u_cpu.REG_FILE._01889_ ),
    .X(\u_cpu.REG_FILE._01890_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06571_  (.A1(\u_cpu.REG_FILE._01351_ ),
    .A2(\u_cpu.REG_FILE.rf[14][14] ),
    .B1(\u_cpu.REG_FILE._01352_ ),
    .C1(\u_cpu.REG_FILE._01890_ ),
    .Y(\u_cpu.REG_FILE._01891_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06572_  (.A1(\u_cpu.REG_FILE._01584_ ),
    .A2(\u_cpu.REG_FILE.rf[12][14] ),
    .B1_N(\u_cpu.REG_FILE._01838_ ),
    .X(\u_cpu.REG_FILE._01892_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06573_  (.A1(\u_cpu.REG_FILE._01787_ ),
    .A2(\u_cpu.REG_FILE.rf[13][14] ),
    .B1(\u_cpu.REG_FILE._01892_ ),
    .Y(\u_cpu.REG_FILE._01893_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06574_  (.A(\u_cpu.REG_FILE._01891_ ),
    .B(\u_cpu.REG_FILE._01893_ ),
    .C(\u_cpu.REG_FILE._01690_ ),
    .Y(\u_cpu.REG_FILE._01894_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06575_  (.A(\u_cpu.REG_FILE._01073_ ),
    .X(\u_cpu.REG_FILE._01895_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06576_  (.A_N(\u_cpu.REG_FILE.rf[9][14] ),
    .B(\u_cpu.REG_FILE._01895_ ),
    .X(\u_cpu.REG_FILE._01896_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06577_  (.A1(\u_cpu.REG_FILE._01475_ ),
    .A2(\u_cpu.REG_FILE.rf[8][14] ),
    .B1_N(\u_cpu.REG_FILE._01843_ ),
    .Y(\u_cpu.REG_FILE._01897_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06578_  (.A(\u_cpu.REG_FILE.rf[11][14] ),
    .B_N(\u_cpu.REG_FILE._01590_ ),
    .X(\u_cpu.REG_FILE._01898_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06579_  (.A1(\u_cpu.REG_FILE._01425_ ),
    .A2(\u_cpu.REG_FILE.rf[10][14] ),
    .B1(\u_cpu.REG_FILE._01360_ ),
    .C1(\u_cpu.REG_FILE._01898_ ),
    .Y(\u_cpu.REG_FILE._01899_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06580_  (.A1(\u_cpu.REG_FILE._01896_ ),
    .A2(\u_cpu.REG_FILE._01897_ ),
    .B1(\u_cpu.REG_FILE._01424_ ),
    .C1(\u_cpu.REG_FILE._01899_ ),
    .Y(\u_cpu.REG_FILE._01900_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06581_  (.A(\u_cpu.REG_FILE._01894_ ),
    .B(\u_cpu.REG_FILE._01900_ ),
    .C(\u_cpu.REG_FILE._01796_ ),
    .Y(\u_cpu.REG_FILE._01901_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06582_  (.A(\u_cpu.REG_FILE.rf[5][14] ),
    .Y(\u_cpu.REG_FILE._01902_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06583_  (.A1(\u_cpu.REG_FILE._01431_ ),
    .A2(\u_cpu.REG_FILE.rf[4][14] ),
    .B1_N(\u_cpu.REG_FILE._01482_ ),
    .Y(\u_cpu.REG_FILE._01903_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._06584_  (.A1(\u_cpu.REG_FILE._01902_ ),
    .A2(\u_cpu.REG_FILE._01850_ ),
    .B1(\u_cpu.REG_FILE._01903_ ),
    .Y(\u_cpu.REG_FILE._01904_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06585_  (.A1(\u_cpu.REG_FILE._01434_ ),
    .A2(\u_cpu.REG_FILE.rf[6][14] ),
    .B1(\u_cpu.REG_FILE._01598_ ),
    .Y(\u_cpu.REG_FILE._01905_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06586_  (.A(\u_cpu.REG_FILE._01073_ ),
    .X(\u_cpu.REG_FILE._01906_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06587_  (.A_N(\u_cpu.REG_FILE.rf[7][14] ),
    .B(\u_cpu.REG_FILE._01906_ ),
    .X(\u_cpu.REG_FILE._01907_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06588_  (.A1(\u_cpu.REG_FILE._01905_ ),
    .A2(\u_cpu.REG_FILE._01907_ ),
    .B1(\u_cpu.REG_FILE._01601_ ),
    .Y(\u_cpu.REG_FILE._01908_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06589_  (.A_N(\u_cpu.REG_FILE.rf[1][14] ),
    .B(\u_cpu.REG_FILE._01804_ ),
    .X(\u_cpu.REG_FILE._01909_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06590_  (.A1(\u_cpu.REG_FILE._01372_ ),
    .A2(\u_cpu.REG_FILE.rf[0][14] ),
    .B1_N(\u_cpu.REG_FILE._01705_ ),
    .Y(\u_cpu.REG_FILE._01910_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06591_  (.A(\u_cpu.REG_FILE.rf[3][14] ),
    .B_N(\u_cpu.REG_FILE._01241_ ),
    .X(\u_cpu.REG_FILE._01911_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06592_  (.A1(\u_cpu.REG_FILE._01707_ ),
    .A2(\u_cpu.REG_FILE.rf[2][14] ),
    .B1(\u_cpu.REG_FILE._01240_ ),
    .C1(\u_cpu.REG_FILE._01911_ ),
    .Y(\u_cpu.REG_FILE._01912_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06593_  (.A1(\u_cpu.REG_FILE._01909_ ),
    .A2(\u_cpu.REG_FILE._01910_ ),
    .B1(\u_cpu.REG_FILE._01858_ ),
    .C1(\u_cpu.REG_FILE._01912_ ),
    .Y(\u_cpu.REG_FILE._01913_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06594_  (.A1(\u_cpu.REG_FILE._01904_ ),
    .A2(\u_cpu.REG_FILE._01908_ ),
    .B1(\u_cpu.REG_FILE._01603_ ),
    .C1(\u_cpu.REG_FILE._01913_ ),
    .Y(\u_cpu.REG_FILE._01914_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._06595_  (.A(\u_cpu.REG_FILE._01901_ ),
    .B(\u_cpu.REG_FILE._01914_ ),
    .Y(\u_cpu.REG_FILE._01915_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06596_  (.A(\u_cpu.REG_FILE.rf[27][14] ),
    .B_N(\u_cpu.REG_FILE._01528_ ),
    .X(\u_cpu.REG_FILE._01916_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06597_  (.A1(\u_cpu.REG_FILE._01105_ ),
    .A2(\u_cpu.REG_FILE.rf[26][14] ),
    .B1(\u_cpu.REG_FILE._01660_ ),
    .C1(\u_cpu.REG_FILE._01916_ ),
    .X(\u_cpu.REG_FILE._01917_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06598_  (.A1(\u_cpu.REG_FILE._01447_ ),
    .A2(\u_cpu.REG_FILE.rf[24][14] ),
    .B1_N(\u_cpu.REG_FILE._01062_ ),
    .X(\u_cpu.REG_FILE._01918_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06599_  (.A(\u_cpu.REG_FILE.rf[25][14] ),
    .B_N(\u_cpu.REG_FILE._01194_ ),
    .X(\u_cpu.REG_FILE._01919_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._06600_  (.A1(\u_cpu.REG_FILE._01918_ ),
    .A2(\u_cpu.REG_FILE._01919_ ),
    .B1(\u_cpu.REG_FILE._01196_ ),
    .X(\u_cpu.REG_FILE._01920_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06601_  (.A(\u_cpu.REG_FILE._01390_ ),
    .B(\u_cpu.REG_FILE.rf[30][14] ),
    .Y(\u_cpu.REG_FILE._01921_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06602_  (.A1(\u_cpu.REG_FILE.rf[31][14] ),
    .A2(\u_cpu.REG_FILE._01200_ ),
    .B1(\u_cpu.REG_FILE._01501_ ),
    .Y(\u_cpu.REG_FILE._01922_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06603_  (.A1(\u_cpu.REG_FILE._01503_ ),
    .A2(\u_cpu.REG_FILE.rf[28][14] ),
    .B1_N(\u_cpu.REG_FILE._01098_ ),
    .X(\u_cpu.REG_FILE._01923_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06604_  (.A1(\u_cpu.REG_FILE._01668_ ),
    .A2(\u_cpu.REG_FILE.rf[29][14] ),
    .B1(\u_cpu.REG_FILE._01923_ ),
    .Y(\u_cpu.REG_FILE._01924_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06605_  (.A1(\u_cpu.REG_FILE._01921_ ),
    .A2(\u_cpu.REG_FILE._01922_ ),
    .B1(\u_cpu.REG_FILE._01924_ ),
    .C1(\u_cpu.REG_FILE._01395_ ),
    .Y(\u_cpu.REG_FILE._01925_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06606_  (.A1(\u_cpu.REG_FILE._01917_ ),
    .A2(\u_cpu.REG_FILE._01920_ ),
    .B1(\u_cpu.REG_FILE._01869_ ),
    .C1(\u_cpu.REG_FILE._01925_ ),
    .Y(\u_cpu.REG_FILE._01926_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06607_  (.A1(\u_cpu.REG_FILE._01206_ ),
    .A2(\u_cpu.REG_FILE.rf[18][14] ),
    .B1(\u_cpu.REG_FILE._01135_ ),
    .Y(\u_cpu.REG_FILE._01927_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06608_  (.A(\u_cpu.REG_FILE.rf[19][14] ),
    .B(\u_cpu.REG_FILE._01509_ ),
    .Y(\u_cpu.REG_FILE._01928_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06609_  (.A1(\u_cpu.REG_FILE._01141_ ),
    .A2(\u_cpu.REG_FILE.rf[16][14] ),
    .B1_N(\u_cpu.REG_FILE._01153_ ),
    .X(\u_cpu.REG_FILE._01929_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06610_  (.A1(\u_cpu.REG_FILE._01726_ ),
    .A2(\u_cpu.REG_FILE.rf[17][14] ),
    .B1(\u_cpu.REG_FILE._01929_ ),
    .Y(\u_cpu.REG_FILE._01930_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06611_  (.A1(\u_cpu.REG_FILE._01927_ ),
    .A2(\u_cpu.REG_FILE._01928_ ),
    .B1(\u_cpu.REG_FILE._01264_ ),
    .C1(\u_cpu.REG_FILE._01930_ ),
    .Y(\u_cpu.REG_FILE._01931_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06612_  (.A(\u_cpu.REG_FILE._01260_ ),
    .B(\u_cpu.REG_FILE.rf[20][14] ),
    .Y(\u_cpu.REG_FILE._01932_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06613_  (.A_N(\u_cpu.REG_FILE.rf[21][14] ),
    .B(\u_cpu.REG_FILE._01262_ ),
    .X(\u_cpu.REG_FILE._01933_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06614_  (.A(\u_cpu.REG_FILE.rf[23][14] ),
    .B_N(\u_cpu.REG_FILE._01408_ ),
    .X(\u_cpu.REG_FILE._01934_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06615_  (.A1(\u_cpu.REG_FILE._01260_ ),
    .A2(\u_cpu.REG_FILE.rf[22][14] ),
    .B1(\u_cpu.REG_FILE._01400_ ),
    .C1(\u_cpu.REG_FILE._01934_ ),
    .Y(\u_cpu.REG_FILE._01935_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._06616_  (.A1(\u_cpu.REG_FILE._01259_ ),
    .A2(\u_cpu.REG_FILE._01932_ ),
    .A3(\u_cpu.REG_FILE._01933_ ),
    .B1(\u_cpu.REG_FILE._01115_ ),
    .C1(\u_cpu.REG_FILE._01935_ ),
    .Y(\u_cpu.REG_FILE._01936_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06617_  (.A(\u_cpu.REG_FILE._01569_ ),
    .B(\u_cpu.REG_FILE._01931_ ),
    .C(\u_cpu.REG_FILE._01936_ ),
    .Y(\u_cpu.REG_FILE._01937_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06618_  (.A(\u_cpu.REG_FILE._01926_ ),
    .B(\u_cpu.REG_FILE._01937_ ),
    .C(\u_cpu.REG_FILE._01684_ ),
    .Y(\u_cpu.REG_FILE._01938_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06619_  (.A1(\u_cpu.REG_FILE._01888_ ),
    .A2(\u_cpu.REG_FILE._01915_ ),
    .B1(\u_cpu.REG_FILE._01938_ ),
    .C1(\u_cpu.REG_FILE._01737_ ),
    .X(\u_cpu.ALU.SrcA[14] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06620_  (.A(\u_cpu.REG_FILE.rf[15][15] ),
    .B_N(\u_cpu.REG_FILE._01889_ ),
    .X(\u_cpu.REG_FILE._01939_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06621_  (.A1(\u_cpu.REG_FILE._01351_ ),
    .A2(\u_cpu.REG_FILE.rf[14][15] ),
    .B1(\u_cpu.REG_FILE._01352_ ),
    .C1(\u_cpu.REG_FILE._01939_ ),
    .Y(\u_cpu.REG_FILE._01940_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06622_  (.A1(\u_cpu.REG_FILE._01584_ ),
    .A2(\u_cpu.REG_FILE.rf[12][15] ),
    .B1_N(\u_cpu.REG_FILE._01838_ ),
    .X(\u_cpu.REG_FILE._01941_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06623_  (.A1(\u_cpu.REG_FILE._01787_ ),
    .A2(\u_cpu.REG_FILE.rf[13][15] ),
    .B1(\u_cpu.REG_FILE._01941_ ),
    .Y(\u_cpu.REG_FILE._01942_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06624_  (.A(\u_cpu.REG_FILE._01940_ ),
    .B(\u_cpu.REG_FILE._01942_ ),
    .C(\u_cpu.REG_FILE._01690_ ),
    .Y(\u_cpu.REG_FILE._01943_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06625_  (.A_N(\u_cpu.REG_FILE.rf[9][15] ),
    .B(\u_cpu.REG_FILE._01895_ ),
    .X(\u_cpu.REG_FILE._01944_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06626_  (.A1(\u_cpu.REG_FILE._01475_ ),
    .A2(\u_cpu.REG_FILE.rf[8][15] ),
    .B1_N(\u_cpu.REG_FILE._01843_ ),
    .Y(\u_cpu.REG_FILE._01945_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06627_  (.A(\u_cpu.REG_FILE.rf[11][15] ),
    .B_N(\u_cpu.REG_FILE._01590_ ),
    .X(\u_cpu.REG_FILE._01946_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06628_  (.A1(\u_cpu.REG_FILE._01425_ ),
    .A2(\u_cpu.REG_FILE.rf[10][15] ),
    .B1(\u_cpu.REG_FILE._01360_ ),
    .C1(\u_cpu.REG_FILE._01946_ ),
    .Y(\u_cpu.REG_FILE._01947_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06629_  (.A1(\u_cpu.REG_FILE._01944_ ),
    .A2(\u_cpu.REG_FILE._01945_ ),
    .B1(\u_cpu.REG_FILE._01424_ ),
    .C1(\u_cpu.REG_FILE._01947_ ),
    .Y(\u_cpu.REG_FILE._01948_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06630_  (.A(\u_cpu.REG_FILE._01943_ ),
    .B(\u_cpu.REG_FILE._01948_ ),
    .C(\u_cpu.REG_FILE._01796_ ),
    .Y(\u_cpu.REG_FILE._01949_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06631_  (.A(\u_cpu.REG_FILE.rf[5][15] ),
    .Y(\u_cpu.REG_FILE._01950_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06632_  (.A1(\u_cpu.REG_FILE._01431_ ),
    .A2(\u_cpu.REG_FILE.rf[4][15] ),
    .B1_N(\u_cpu.REG_FILE._01482_ ),
    .Y(\u_cpu.REG_FILE._01951_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._06633_  (.A1(\u_cpu.REG_FILE._01950_ ),
    .A2(\u_cpu.REG_FILE._01850_ ),
    .B1(\u_cpu.REG_FILE._01951_ ),
    .Y(\u_cpu.REG_FILE._01952_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06634_  (.A1(\u_cpu.REG_FILE._01434_ ),
    .A2(\u_cpu.REG_FILE.rf[6][15] ),
    .B1(\u_cpu.REG_FILE._01598_ ),
    .Y(\u_cpu.REG_FILE._01953_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06635_  (.A_N(\u_cpu.REG_FILE.rf[7][15] ),
    .B(\u_cpu.REG_FILE._01906_ ),
    .X(\u_cpu.REG_FILE._01954_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06636_  (.A1(\u_cpu.REG_FILE._01953_ ),
    .A2(\u_cpu.REG_FILE._01954_ ),
    .B1(\u_cpu.REG_FILE._01601_ ),
    .Y(\u_cpu.REG_FILE._01955_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06637_  (.A_N(\u_cpu.REG_FILE.rf[1][15] ),
    .B(\u_cpu.REG_FILE._01804_ ),
    .X(\u_cpu.REG_FILE._01956_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06638_  (.A1(\u_cpu.REG_FILE._01372_ ),
    .A2(\u_cpu.REG_FILE.rf[0][15] ),
    .B1_N(\u_cpu.REG_FILE._01705_ ),
    .Y(\u_cpu.REG_FILE._01957_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06639_  (.A(\u_cpu.REG_FILE.rf[3][15] ),
    .B_N(\u_cpu.REG_FILE._01241_ ),
    .X(\u_cpu.REG_FILE._01958_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06640_  (.A1(\u_cpu.REG_FILE._01707_ ),
    .A2(\u_cpu.REG_FILE.rf[2][15] ),
    .B1(\u_cpu.REG_FILE._01240_ ),
    .C1(\u_cpu.REG_FILE._01958_ ),
    .Y(\u_cpu.REG_FILE._01959_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06641_  (.A1(\u_cpu.REG_FILE._01956_ ),
    .A2(\u_cpu.REG_FILE._01957_ ),
    .B1(\u_cpu.REG_FILE._01858_ ),
    .C1(\u_cpu.REG_FILE._01959_ ),
    .Y(\u_cpu.REG_FILE._01960_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06642_  (.A1(\u_cpu.REG_FILE._01952_ ),
    .A2(\u_cpu.REG_FILE._01955_ ),
    .B1(\u_cpu.REG_FILE._01603_ ),
    .C1(\u_cpu.REG_FILE._01960_ ),
    .Y(\u_cpu.REG_FILE._01961_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._06643_  (.A(\u_cpu.REG_FILE._01949_ ),
    .B(\u_cpu.REG_FILE._01961_ ),
    .Y(\u_cpu.REG_FILE._01962_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06644_  (.A1(\u_cpu.REG_FILE._01379_ ),
    .A2(\u_cpu.REG_FILE.rf[24][15] ),
    .B1_N(\u_cpu.REG_FILE._01611_ ),
    .Y(\u_cpu.REG_FILE._01963_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06645_  (.A_N(\u_cpu.REG_FILE.rf[25][15] ),
    .B(\u_cpu.REG_FILE._01382_ ),
    .X(\u_cpu.REG_FILE._01964_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06646_  (.A1(\u_cpu.REG_FILE._01963_ ),
    .A2(\u_cpu.REG_FILE._01964_ ),
    .B1(\u_cpu.REG_FILE._01814_ ),
    .Y(\u_cpu.REG_FILE._01965_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06647_  (.A(\u_cpu.REG_FILE._01340_ ),
    .B(\u_cpu.REG_FILE.rf[26][15] ),
    .X(\u_cpu.REG_FILE._01966_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06648_  (.A1(\u_cpu.REG_FILE._01386_ ),
    .A2(\u_cpu.REG_FILE.rf[27][15] ),
    .B1(\u_cpu.REG_FILE._01387_ ),
    .C1(\u_cpu.REG_FILE._01966_ ),
    .X(\u_cpu.REG_FILE._01967_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06649_  (.A(\u_cpu.REG_FILE._01390_ ),
    .B(\u_cpu.REG_FILE.rf[30][15] ),
    .Y(\u_cpu.REG_FILE._01968_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06650_  (.A(\u_cpu.REG_FILE._01123_ ),
    .X(\u_cpu.REG_FILE._01969_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06651_  (.A1(\u_cpu.REG_FILE.rf[31][15] ),
    .A2(\u_cpu.REG_FILE._01969_ ),
    .B1(\u_cpu.REG_FILE._01501_ ),
    .Y(\u_cpu.REG_FILE._01970_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06652_  (.A1(\u_cpu.REG_FILE._01503_ ),
    .A2(\u_cpu.REG_FILE.rf[28][15] ),
    .B1_N(\u_cpu.REG_FILE._01098_ ),
    .X(\u_cpu.REG_FILE._01971_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06653_  (.A1(\u_cpu.REG_FILE._01668_ ),
    .A2(\u_cpu.REG_FILE.rf[29][15] ),
    .B1(\u_cpu.REG_FILE._01971_ ),
    .Y(\u_cpu.REG_FILE._01972_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06654_  (.A1(\u_cpu.REG_FILE._01968_ ),
    .A2(\u_cpu.REG_FILE._01970_ ),
    .B1(\u_cpu.REG_FILE._01972_ ),
    .C1(\u_cpu.REG_FILE._01395_ ),
    .Y(\u_cpu.REG_FILE._01973_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06655_  (.A1(\u_cpu.REG_FILE._01965_ ),
    .A2(\u_cpu.REG_FILE._01967_ ),
    .B1(\u_cpu.REG_FILE._01869_ ),
    .C1(\u_cpu.REG_FILE._01973_ ),
    .Y(\u_cpu.REG_FILE._01974_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06656_  (.A(\u_cpu.REG_FILE.rf[19][15] ),
    .Y(\u_cpu.REG_FILE._01975_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06657_  (.A1(\u_cpu.REG_FILE._01317_ ),
    .A2(\u_cpu.REG_FILE.rf[18][15] ),
    .B1(\u_cpu.REG_FILE._01533_ ),
    .Y(\u_cpu.REG_FILE._01976_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._06658_  (.A1(\u_cpu.REG_FILE._01975_ ),
    .A2(\u_cpu.REG_FILE._01399_ ),
    .B1(\u_cpu.REG_FILE._01976_ ),
    .Y(\u_cpu.REG_FILE._01977_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06659_  (.A(\u_cpu.REG_FILE.rf[17][15] ),
    .Y(\u_cpu.REG_FILE._01978_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06660_  (.A1(\u_cpu.REG_FILE._01404_ ),
    .A2(\u_cpu.REG_FILE.rf[16][15] ),
    .B1_N(\u_cpu.REG_FILE._01258_ ),
    .Y(\u_cpu.REG_FILE._01979_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._06661_  (.A1(\u_cpu.REG_FILE._01978_ ),
    .A2(\u_cpu.REG_FILE._01284_ ),
    .B1(\u_cpu.REG_FILE._01979_ ),
    .Y(\u_cpu.REG_FILE._01980_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06662_  (.A(\u_cpu.REG_FILE.rf[23][15] ),
    .B_N(\u_cpu.REG_FILE._01408_ ),
    .X(\u_cpu.REG_FILE._01981_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06663_  (.A1(\u_cpu.REG_FILE._01077_ ),
    .A2(\u_cpu.REG_FILE.rf[22][15] ),
    .B1(\u_cpu.REG_FILE._01407_ ),
    .C1(\u_cpu.REG_FILE._01981_ ),
    .Y(\u_cpu.REG_FILE._01982_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06664_  (.A1(\u_cpu.REG_FILE._01324_ ),
    .A2(\u_cpu.REG_FILE.rf[20][15] ),
    .B1_N(\u_cpu.REG_FILE._01304_ ),
    .X(\u_cpu.REG_FILE._01983_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06665_  (.A1(\u_cpu.REG_FILE._01038_ ),
    .A2(\u_cpu.REG_FILE.rf[21][15] ),
    .B1(\u_cpu.REG_FILE._01983_ ),
    .Y(\u_cpu.REG_FILE._01984_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06666_  (.A(\u_cpu.REG_FILE._01982_ ),
    .B(\u_cpu.REG_FILE._01984_ ),
    .C(\u_cpu.REG_FILE._01115_ ),
    .Y(\u_cpu.REG_FILE._01985_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._06667_  (.A1(\u_cpu.REG_FILE._01277_ ),
    .A2(\u_cpu.REG_FILE._01977_ ),
    .A3(\u_cpu.REG_FILE._01980_ ),
    .B1(\u_cpu.REG_FILE._01985_ ),
    .C1(\u_cpu.REG_FILE._01414_ ),
    .Y(\u_cpu.REG_FILE._01986_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06668_  (.A(\u_cpu.REG_FILE._01974_ ),
    .B(\u_cpu.REG_FILE._01986_ ),
    .C(\u_cpu.REG_FILE._01684_ ),
    .Y(\u_cpu.REG_FILE._01987_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06669_  (.A1(\u_cpu.REG_FILE._01888_ ),
    .A2(\u_cpu.REG_FILE._01962_ ),
    .B1(\u_cpu.REG_FILE._01987_ ),
    .C1(\u_cpu.REG_FILE._01737_ ),
    .X(\u_cpu.ALU.SrcA[15] ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06670_  (.A1(\u_cpu.REG_FILE._01404_ ),
    .A2(\u_cpu.REG_FILE.rf[16][16] ),
    .B1_N(\u_cpu.REG_FILE._01553_ ),
    .Y(\u_cpu.REG_FILE._01988_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06671_  (.A_N(\u_cpu.REG_FILE.rf[17][16] ),
    .B(\u_cpu.REG_FILE._01750_ ),
    .X(\u_cpu.REG_FILE._01989_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06672_  (.A1(\u_cpu.REG_FILE._01279_ ),
    .A2(\u_cpu.REG_FILE.rf[18][16] ),
    .B1(\u_cpu.REG_FILE._01280_ ),
    .Y(\u_cpu.REG_FILE._01990_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06673_  (.A_N(\u_cpu.REG_FILE.rf[19][16] ),
    .B(\u_cpu.REG_FILE._01523_ ),
    .X(\u_cpu.REG_FILE._01991_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.REG_FILE._06674_  (.A1(\u_cpu.REG_FILE._01988_ ),
    .A2(\u_cpu.REG_FILE._01989_ ),
    .B1(\u_cpu.REG_FILE._01990_ ),
    .B2(\u_cpu.REG_FILE._01991_ ),
    .Y(\u_cpu.REG_FILE._01992_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06675_  (.A(\u_cpu.REG_FILE._01118_ ),
    .B(\u_cpu.REG_FILE.rf[20][16] ),
    .Y(\u_cpu.REG_FILE._01993_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06676_  (.A1(\u_cpu.REG_FILE.rf[21][16] ),
    .A2(\u_cpu.REG_FILE._01287_ ),
    .B1_N(\u_cpu.REG_FILE._01305_ ),
    .Y(\u_cpu.REG_FILE._01994_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06677_  (.A(\u_cpu.REG_FILE._01536_ ),
    .B(\u_cpu.REG_FILE.rf[22][16] ),
    .X(\u_cpu.REG_FILE._01995_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06678_  (.A1(\u_cpu.REG_FILE._01535_ ),
    .A2(\u_cpu.REG_FILE.rf[23][16] ),
    .B1(\u_cpu.REG_FILE._01527_ ),
    .C1(\u_cpu.REG_FILE._01995_ ),
    .Y(\u_cpu.REG_FILE._01996_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06679_  (.A1(\u_cpu.REG_FILE._01993_ ),
    .A2(\u_cpu.REG_FILE._01994_ ),
    .B1(\u_cpu.REG_FILE._01129_ ),
    .C1(\u_cpu.REG_FILE._01996_ ),
    .Y(\u_cpu.REG_FILE._01997_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06680_  (.A1(\u_cpu.REG_FILE._01992_ ),
    .A2(\u_cpu.REG_FILE._01277_ ),
    .B1(\u_cpu.REG_FILE._01541_ ),
    .C1(\u_cpu.REG_FILE._01997_ ),
    .X(\u_cpu.REG_FILE._01998_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06681_  (.A(\u_cpu.REG_FILE.rf[31][16] ),
    .B_N(\u_cpu.REG_FILE._01111_ ),
    .X(\u_cpu.REG_FILE._01999_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06682_  (.A1(\u_cpu.REG_FILE._01030_ ),
    .A2(\u_cpu.REG_FILE.rf[30][16] ),
    .B1(\u_cpu.REG_FILE._01033_ ),
    .C1(\u_cpu.REG_FILE._01999_ ),
    .Y(\u_cpu.REG_FILE._02000_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06683_  (.A1(\u_cpu.REG_FILE._01299_ ),
    .A2(\u_cpu.REG_FILE.rf[28][16] ),
    .B1_N(\u_cpu.REG_FILE._01106_ ),
    .X(\u_cpu.REG_FILE._02001_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06684_  (.A1(\u_cpu.REG_FILE._01298_ ),
    .A2(\u_cpu.REG_FILE.rf[29][16] ),
    .B1(\u_cpu.REG_FILE._02001_ ),
    .Y(\u_cpu.REG_FILE._02002_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06685_  (.A(\u_cpu.REG_FILE._02000_ ),
    .B(\u_cpu.REG_FILE._02002_ ),
    .C(\u_cpu.REG_FILE._01293_ ),
    .Y(\u_cpu.REG_FILE._02003_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06686_  (.A_N(\u_cpu.REG_FILE.rf[25][16] ),
    .B(\u_cpu.REG_FILE._01547_ ),
    .X(\u_cpu.REG_FILE._02004_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06687_  (.A1(\u_cpu.REG_FILE._01093_ ),
    .A2(\u_cpu.REG_FILE.rf[24][16] ),
    .B1_N(\u_cpu.REG_FILE._01550_ ),
    .Y(\u_cpu.REG_FILE._02005_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06688_  (.A(\u_cpu.REG_FILE.rf[27][16] ),
    .B_N(\u_cpu.REG_FILE._01310_ ),
    .X(\u_cpu.REG_FILE._02006_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06689_  (.A1(\u_cpu.REG_FILE._01308_ ),
    .A2(\u_cpu.REG_FILE.rf[26][16] ),
    .B1(\u_cpu.REG_FILE._01309_ ),
    .C1(\u_cpu.REG_FILE._02006_ ),
    .Y(\u_cpu.REG_FILE._02007_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06690_  (.A1(\u_cpu.REG_FILE._02004_ ),
    .A2(\u_cpu.REG_FILE._02005_ ),
    .B1(\u_cpu.REG_FILE._01059_ ),
    .C1(\u_cpu.REG_FILE._02007_ ),
    .Y(\u_cpu.REG_FILE._02008_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._06691_  (.A1(\u_cpu.REG_FILE._02003_ ),
    .A2(\u_cpu.REG_FILE._02008_ ),
    .A3(\u_cpu.REG_FILE._01314_ ),
    .B1(\u_cpu.REG_FILE._01315_ ),
    .X(\u_cpu.REG_FILE._02009_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06692_  (.A(\u_cpu.REG_FILE._01330_ ),
    .X(\u_cpu.REG_FILE._02010_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06693_  (.A(\u_cpu.REG_FILE._02010_ ),
    .B(\u_cpu.REG_FILE.rf[14][16] ),
    .Y(\u_cpu.REG_FILE._02011_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06694_  (.A1(\u_cpu.REG_FILE.rf[15][16] ),
    .A2(\u_cpu.REG_FILE._01969_ ),
    .B1(\u_cpu.REG_FILE._01660_ ),
    .Y(\u_cpu.REG_FILE._02012_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06695_  (.A(\u_cpu.REG_FILE._01028_ ),
    .X(\u_cpu.REG_FILE._02013_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06696_  (.A1(\u_cpu.REG_FILE._02013_ ),
    .A2(\u_cpu.REG_FILE.rf[12][16] ),
    .B1_N(\u_cpu.REG_FILE._01142_ ),
    .X(\u_cpu.REG_FILE._02014_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06697_  (.A1(\u_cpu.REG_FILE._01140_ ),
    .A2(\u_cpu.REG_FILE.rf[13][16] ),
    .B1(\u_cpu.REG_FILE._02014_ ),
    .Y(\u_cpu.REG_FILE._02015_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06698_  (.A(\u_cpu.REG_FILE._01046_ ),
    .X(\u_cpu.REG_FILE._02016_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06699_  (.A1(\u_cpu.REG_FILE._02011_ ),
    .A2(\u_cpu.REG_FILE._02012_ ),
    .B1(\u_cpu.REG_FILE._02015_ ),
    .C1(\u_cpu.REG_FILE._02016_ ),
    .Y(\u_cpu.REG_FILE._02017_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06700_  (.A(\u_cpu.REG_FILE._01052_ ),
    .X(\u_cpu.REG_FILE._02018_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06701_  (.A(\u_cpu.REG_FILE.rf[11][16] ),
    .B_N(\u_cpu.REG_FILE._01148_ ),
    .X(\u_cpu.REG_FILE._02019_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06702_  (.A1(\u_cpu.REG_FILE._02018_ ),
    .A2(\u_cpu.REG_FILE.rf[10][16] ),
    .B1(\u_cpu.REG_FILE._01618_ ),
    .C1(\u_cpu.REG_FILE._02019_ ),
    .Y(\u_cpu.REG_FILE._02020_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06703_  (.A1(\u_cpu.REG_FILE._01536_ ),
    .A2(\u_cpu.REG_FILE.rf[8][16] ),
    .B1_N(\u_cpu.REG_FILE._01134_ ),
    .X(\u_cpu.REG_FILE._02021_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06704_  (.A1(\u_cpu.REG_FILE._01120_ ),
    .A2(\u_cpu.REG_FILE.rf[9][16] ),
    .B1(\u_cpu.REG_FILE._02021_ ),
    .Y(\u_cpu.REG_FILE._02022_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06705_  (.A(\u_cpu.REG_FILE._01525_ ),
    .B(\u_cpu.REG_FILE._02020_ ),
    .C(\u_cpu.REG_FILE._02022_ ),
    .Y(\u_cpu.REG_FILE._02023_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06706_  (.A(\u_cpu.REG_FILE._02017_ ),
    .B(\u_cpu.REG_FILE._02023_ ),
    .C(\u_cpu.REG_FILE._01314_ ),
    .Y(\u_cpu.REG_FILE._02024_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06707_  (.A(\u_cpu.REG_FILE.rf[3][16] ),
    .B_N(\u_cpu.REG_FILE._01148_ ),
    .X(\u_cpu.REG_FILE._02025_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06708_  (.A1(\u_cpu.REG_FILE._02018_ ),
    .A2(\u_cpu.REG_FILE.rf[2][16] ),
    .B1(\u_cpu.REG_FILE._01618_ ),
    .C1(\u_cpu.REG_FILE._02025_ ),
    .Y(\u_cpu.REG_FILE._02026_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06709_  (.A1(\u_cpu.REG_FILE._01152_ ),
    .A2(\u_cpu.REG_FILE.rf[0][16] ),
    .B1_N(\u_cpu.REG_FILE._01153_ ),
    .X(\u_cpu.REG_FILE._02027_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06710_  (.A1(\u_cpu.REG_FILE._01726_ ),
    .A2(\u_cpu.REG_FILE.rf[1][16] ),
    .B1(\u_cpu.REG_FILE._02027_ ),
    .Y(\u_cpu.REG_FILE._02028_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06711_  (.A(\u_cpu.REG_FILE._01525_ ),
    .B(\u_cpu.REG_FILE._02026_ ),
    .C(\u_cpu.REG_FILE._02028_ ),
    .Y(\u_cpu.REG_FILE._02029_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06712_  (.A1(\u_cpu.REG_FILE._01029_ ),
    .A2(\u_cpu.REG_FILE.rf[4][16] ),
    .B1_N(\u_cpu.REG_FILE._01239_ ),
    .X(\u_cpu.REG_FILE._02030_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06713_  (.A1(\u_cpu.REG_FILE._01137_ ),
    .A2(\u_cpu.REG_FILE.rf[5][16] ),
    .B1(\u_cpu.REG_FILE._02030_ ),
    .Y(\u_cpu.REG_FILE._02031_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.REG_FILE._06714_  (.A1(\u_cpu.REG_FILE._02013_ ),
    .A2(\u_cpu.REG_FILE.rf[6][16] ),
    .B1(\u_cpu.REG_FILE._01032_ ),
    .X(\u_cpu.REG_FILE._02032_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06715_  (.A1(\u_cpu.REG_FILE.rf[7][16] ),
    .A2(\u_cpu.REG_FILE._01386_ ),
    .B1(\u_cpu.REG_FILE._02032_ ),
    .Y(\u_cpu.REG_FILE._02033_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06716_  (.A(\u_cpu.REG_FILE._02031_ ),
    .B(\u_cpu.REG_FILE._01156_ ),
    .C(\u_cpu.REG_FILE._02033_ ),
    .Y(\u_cpu.REG_FILE._02034_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06717_  (.A(\u_cpu.REG_FILE._01132_ ),
    .B(\u_cpu.REG_FILE._02029_ ),
    .C(\u_cpu.REG_FILE._02034_ ),
    .Y(\u_cpu.REG_FILE._02035_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06718_  (.A(\u_cpu.REG_FILE._01315_ ),
    .B(\u_cpu.REG_FILE._02024_ ),
    .C(\u_cpu.REG_FILE._02035_ ),
    .Y(\u_cpu.REG_FILE._02036_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06719_  (.A1(\u_cpu.REG_FILE._01998_ ),
    .A2(\u_cpu.REG_FILE._02009_ ),
    .B1(\u_cpu.REG_FILE._02036_ ),
    .C1(\u_cpu.REG_FILE._01737_ ),
    .X(\u_cpu.ALU.SrcA[16] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06720_  (.A(\u_cpu.REG_FILE.rf[15][17] ),
    .B_N(\u_cpu.REG_FILE._01889_ ),
    .X(\u_cpu.REG_FILE._02037_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06721_  (.A1(\u_cpu.REG_FILE._01351_ ),
    .A2(\u_cpu.REG_FILE.rf[14][17] ),
    .B1(\u_cpu.REG_FILE._01352_ ),
    .C1(\u_cpu.REG_FILE._02037_ ),
    .Y(\u_cpu.REG_FILE._02038_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06722_  (.A1(\u_cpu.REG_FILE._01584_ ),
    .A2(\u_cpu.REG_FILE.rf[12][17] ),
    .B1_N(\u_cpu.REG_FILE._01838_ ),
    .X(\u_cpu.REG_FILE._02039_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06723_  (.A1(\u_cpu.REG_FILE._01787_ ),
    .A2(\u_cpu.REG_FILE.rf[13][17] ),
    .B1(\u_cpu.REG_FILE._02039_ ),
    .Y(\u_cpu.REG_FILE._02040_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06724_  (.A(\u_cpu.REG_FILE._02038_ ),
    .B(\u_cpu.REG_FILE._02040_ ),
    .C(\u_cpu.REG_FILE._01690_ ),
    .Y(\u_cpu.REG_FILE._02041_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06725_  (.A_N(\u_cpu.REG_FILE.rf[9][17] ),
    .B(\u_cpu.REG_FILE._01895_ ),
    .X(\u_cpu.REG_FILE._02042_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06726_  (.A1(\u_cpu.REG_FILE._01475_ ),
    .A2(\u_cpu.REG_FILE.rf[8][17] ),
    .B1_N(\u_cpu.REG_FILE._01843_ ),
    .Y(\u_cpu.REG_FILE._02043_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06727_  (.A(\u_cpu.REG_FILE.rf[11][17] ),
    .B_N(\u_cpu.REG_FILE._01590_ ),
    .X(\u_cpu.REG_FILE._02044_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06728_  (.A1(\u_cpu.REG_FILE._01425_ ),
    .A2(\u_cpu.REG_FILE.rf[10][17] ),
    .B1(\u_cpu.REG_FILE._01360_ ),
    .C1(\u_cpu.REG_FILE._02044_ ),
    .Y(\u_cpu.REG_FILE._02045_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06729_  (.A1(\u_cpu.REG_FILE._02042_ ),
    .A2(\u_cpu.REG_FILE._02043_ ),
    .B1(\u_cpu.REG_FILE._01424_ ),
    .C1(\u_cpu.REG_FILE._02045_ ),
    .Y(\u_cpu.REG_FILE._02046_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06730_  (.A(\u_cpu.REG_FILE._02041_ ),
    .B(\u_cpu.REG_FILE._02046_ ),
    .C(\u_cpu.REG_FILE._01796_ ),
    .Y(\u_cpu.REG_FILE._02047_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06731_  (.A(\u_cpu.REG_FILE.rf[5][17] ),
    .Y(\u_cpu.REG_FILE._02048_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06732_  (.A1(\u_cpu.REG_FILE._01431_ ),
    .A2(\u_cpu.REG_FILE.rf[4][17] ),
    .B1_N(\u_cpu.REG_FILE._01482_ ),
    .Y(\u_cpu.REG_FILE._02049_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._06733_  (.A1(\u_cpu.REG_FILE._02048_ ),
    .A2(\u_cpu.REG_FILE._01850_ ),
    .B1(\u_cpu.REG_FILE._02049_ ),
    .Y(\u_cpu.REG_FILE._02050_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06734_  (.A1(\u_cpu.REG_FILE._01434_ ),
    .A2(\u_cpu.REG_FILE.rf[6][17] ),
    .B1(\u_cpu.REG_FILE._01598_ ),
    .Y(\u_cpu.REG_FILE._02051_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06735_  (.A_N(\u_cpu.REG_FILE.rf[7][17] ),
    .B(\u_cpu.REG_FILE._01906_ ),
    .X(\u_cpu.REG_FILE._02052_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06736_  (.A1(\u_cpu.REG_FILE._02051_ ),
    .A2(\u_cpu.REG_FILE._02052_ ),
    .B1(\u_cpu.REG_FILE._01601_ ),
    .Y(\u_cpu.REG_FILE._02053_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06737_  (.A_N(\u_cpu.REG_FILE.rf[1][17] ),
    .B(\u_cpu.REG_FILE._01804_ ),
    .X(\u_cpu.REG_FILE._02054_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06738_  (.A1(\u_cpu.REG_FILE._01372_ ),
    .A2(\u_cpu.REG_FILE.rf[0][17] ),
    .B1_N(\u_cpu.REG_FILE._01705_ ),
    .Y(\u_cpu.REG_FILE._02055_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06739_  (.A(\u_cpu.REG_FILE._01239_ ),
    .X(\u_cpu.REG_FILE._02056_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06740_  (.A(\u_cpu.REG_FILE._01040_ ),
    .X(\u_cpu.REG_FILE._02057_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06741_  (.A(\u_cpu.REG_FILE.rf[3][17] ),
    .B_N(\u_cpu.REG_FILE._02057_ ),
    .X(\u_cpu.REG_FILE._02058_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06742_  (.A1(\u_cpu.REG_FILE._01707_ ),
    .A2(\u_cpu.REG_FILE.rf[2][17] ),
    .B1(\u_cpu.REG_FILE._02056_ ),
    .C1(\u_cpu.REG_FILE._02058_ ),
    .Y(\u_cpu.REG_FILE._02059_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06743_  (.A1(\u_cpu.REG_FILE._02054_ ),
    .A2(\u_cpu.REG_FILE._02055_ ),
    .B1(\u_cpu.REG_FILE._01858_ ),
    .C1(\u_cpu.REG_FILE._02059_ ),
    .Y(\u_cpu.REG_FILE._02060_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06744_  (.A1(\u_cpu.REG_FILE._02050_ ),
    .A2(\u_cpu.REG_FILE._02053_ ),
    .B1(\u_cpu.REG_FILE._01603_ ),
    .C1(\u_cpu.REG_FILE._02060_ ),
    .Y(\u_cpu.REG_FILE._02061_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._06745_  (.A(\u_cpu.REG_FILE._02047_ ),
    .B(\u_cpu.REG_FILE._02061_ ),
    .Y(\u_cpu.REG_FILE._02062_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06746_  (.A1(\u_cpu.REG_FILE._01379_ ),
    .A2(\u_cpu.REG_FILE.rf[24][17] ),
    .B1_N(\u_cpu.REG_FILE._01611_ ),
    .Y(\u_cpu.REG_FILE._02063_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06747_  (.A_N(\u_cpu.REG_FILE.rf[25][17] ),
    .B(\u_cpu.REG_FILE._01382_ ),
    .X(\u_cpu.REG_FILE._02064_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06748_  (.A1(\u_cpu.REG_FILE._02063_ ),
    .A2(\u_cpu.REG_FILE._02064_ ),
    .B1(\u_cpu.REG_FILE._01814_ ),
    .Y(\u_cpu.REG_FILE._02065_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06749_  (.A(\u_cpu.REG_FILE._01340_ ),
    .B(\u_cpu.REG_FILE.rf[26][17] ),
    .X(\u_cpu.REG_FILE._02066_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06750_  (.A1(\u_cpu.REG_FILE._01386_ ),
    .A2(\u_cpu.REG_FILE.rf[27][17] ),
    .B1(\u_cpu.REG_FILE._01387_ ),
    .C1(\u_cpu.REG_FILE._02066_ ),
    .X(\u_cpu.REG_FILE._02067_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06751_  (.A(\u_cpu.REG_FILE._01390_ ),
    .B(\u_cpu.REG_FILE.rf[30][17] ),
    .Y(\u_cpu.REG_FILE._02068_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06752_  (.A1(\u_cpu.REG_FILE.rf[31][17] ),
    .A2(\u_cpu.REG_FILE._01969_ ),
    .B1(\u_cpu.REG_FILE._01501_ ),
    .Y(\u_cpu.REG_FILE._02069_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06753_  (.A1(\u_cpu.REG_FILE._01503_ ),
    .A2(\u_cpu.REG_FILE.rf[28][17] ),
    .B1_N(\u_cpu.REG_FILE._01098_ ),
    .X(\u_cpu.REG_FILE._02070_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06754_  (.A1(\u_cpu.REG_FILE._01668_ ),
    .A2(\u_cpu.REG_FILE.rf[29][17] ),
    .B1(\u_cpu.REG_FILE._02070_ ),
    .Y(\u_cpu.REG_FILE._02071_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06755_  (.A1(\u_cpu.REG_FILE._02068_ ),
    .A2(\u_cpu.REG_FILE._02069_ ),
    .B1(\u_cpu.REG_FILE._02071_ ),
    .C1(\u_cpu.REG_FILE._01395_ ),
    .Y(\u_cpu.REG_FILE._02072_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06756_  (.A1(\u_cpu.REG_FILE._02065_ ),
    .A2(\u_cpu.REG_FILE._02067_ ),
    .B1(\u_cpu.REG_FILE._01869_ ),
    .C1(\u_cpu.REG_FILE._02072_ ),
    .Y(\u_cpu.REG_FILE._02073_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06757_  (.A(\u_cpu.REG_FILE.rf[19][17] ),
    .Y(\u_cpu.REG_FILE._02074_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06758_  (.A1(\u_cpu.REG_FILE._01523_ ),
    .A2(\u_cpu.REG_FILE.rf[18][17] ),
    .B1(\u_cpu.REG_FILE._01533_ ),
    .Y(\u_cpu.REG_FILE._02075_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._06759_  (.A1(\u_cpu.REG_FILE._02074_ ),
    .A2(\u_cpu.REG_FILE._01399_ ),
    .B1(\u_cpu.REG_FILE._02075_ ),
    .Y(\u_cpu.REG_FILE._02076_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06760_  (.A(\u_cpu.REG_FILE.rf[17][17] ),
    .Y(\u_cpu.REG_FILE._02077_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06761_  (.A1(\u_cpu.REG_FILE._01404_ ),
    .A2(\u_cpu.REG_FILE.rf[16][17] ),
    .B1_N(\u_cpu.REG_FILE._01258_ ),
    .Y(\u_cpu.REG_FILE._02078_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._06762_  (.A1(\u_cpu.REG_FILE._02077_ ),
    .A2(\u_cpu.REG_FILE._01399_ ),
    .B1(\u_cpu.REG_FILE._02078_ ),
    .Y(\u_cpu.REG_FILE._02079_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06763_  (.A(\u_cpu.REG_FILE.rf[23][17] ),
    .B_N(\u_cpu.REG_FILE._01408_ ),
    .X(\u_cpu.REG_FILE._02080_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06764_  (.A1(\u_cpu.REG_FILE._01077_ ),
    .A2(\u_cpu.REG_FILE.rf[22][17] ),
    .B1(\u_cpu.REG_FILE._01407_ ),
    .C1(\u_cpu.REG_FILE._02080_ ),
    .Y(\u_cpu.REG_FILE._02081_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06765_  (.A1(\u_cpu.REG_FILE._01324_ ),
    .A2(\u_cpu.REG_FILE.rf[20][17] ),
    .B1_N(\u_cpu.REG_FILE._01304_ ),
    .X(\u_cpu.REG_FILE._02082_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06766_  (.A1(\u_cpu.REG_FILE._01038_ ),
    .A2(\u_cpu.REG_FILE.rf[21][17] ),
    .B1(\u_cpu.REG_FILE._02082_ ),
    .Y(\u_cpu.REG_FILE._02083_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06767_  (.A(\u_cpu.REG_FILE._02081_ ),
    .B(\u_cpu.REG_FILE._02083_ ),
    .C(\u_cpu.REG_FILE._01115_ ),
    .Y(\u_cpu.REG_FILE._02084_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._06768_  (.A1(\u_cpu.REG_FILE._01277_ ),
    .A2(\u_cpu.REG_FILE._02076_ ),
    .A3(\u_cpu.REG_FILE._02079_ ),
    .B1(\u_cpu.REG_FILE._02084_ ),
    .C1(\u_cpu.REG_FILE._01414_ ),
    .Y(\u_cpu.REG_FILE._02085_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06769_  (.A(\u_cpu.REG_FILE._02073_ ),
    .B(\u_cpu.REG_FILE._02085_ ),
    .C(\u_cpu.REG_FILE._01684_ ),
    .Y(\u_cpu.REG_FILE._02086_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06770_  (.A1(\u_cpu.REG_FILE._01888_ ),
    .A2(\u_cpu.REG_FILE._02062_ ),
    .B1(\u_cpu.REG_FILE._02086_ ),
    .C1(\u_cpu.REG_FILE._01737_ ),
    .X(\u_cpu.ALU.SrcA[17] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06771_  (.A(\u_cpu.REG_FILE.rf[15][18] ),
    .B_N(\u_cpu.REG_FILE._01889_ ),
    .X(\u_cpu.REG_FILE._02087_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06772_  (.A1(\u_cpu.REG_FILE._01531_ ),
    .A2(\u_cpu.REG_FILE.rf[14][18] ),
    .B1(\u_cpu.REG_FILE._01288_ ),
    .C1(\u_cpu.REG_FILE._02087_ ),
    .Y(\u_cpu.REG_FILE._02088_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06773_  (.A1(\u_cpu.REG_FILE._01584_ ),
    .A2(\u_cpu.REG_FILE.rf[12][18] ),
    .B1_N(\u_cpu.REG_FILE._01838_ ),
    .X(\u_cpu.REG_FILE._02089_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06774_  (.A1(\u_cpu.REG_FILE._01787_ ),
    .A2(\u_cpu.REG_FILE.rf[13][18] ),
    .B1(\u_cpu.REG_FILE._02089_ ),
    .Y(\u_cpu.REG_FILE._02090_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06775_  (.A(\u_cpu.REG_FILE._02088_ ),
    .B(\u_cpu.REG_FILE._02090_ ),
    .C(\u_cpu.REG_FILE._01690_ ),
    .Y(\u_cpu.REG_FILE._02091_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06776_  (.A_N(\u_cpu.REG_FILE.rf[9][18] ),
    .B(\u_cpu.REG_FILE._01895_ ),
    .X(\u_cpu.REG_FILE._02092_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06777_  (.A1(\u_cpu.REG_FILE._01475_ ),
    .A2(\u_cpu.REG_FILE.rf[8][18] ),
    .B1_N(\u_cpu.REG_FILE._01843_ ),
    .Y(\u_cpu.REG_FILE._02093_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06778_  (.A(\u_cpu.REG_FILE.rf[11][18] ),
    .B_N(\u_cpu.REG_FILE._01590_ ),
    .X(\u_cpu.REG_FILE._02094_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06779_  (.A1(\u_cpu.REG_FILE._01425_ ),
    .A2(\u_cpu.REG_FILE.rf[10][18] ),
    .B1(\u_cpu.REG_FILE._01339_ ),
    .C1(\u_cpu.REG_FILE._02094_ ),
    .Y(\u_cpu.REG_FILE._02095_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06780_  (.A1(\u_cpu.REG_FILE._02092_ ),
    .A2(\u_cpu.REG_FILE._02093_ ),
    .B1(\u_cpu.REG_FILE._01424_ ),
    .C1(\u_cpu.REG_FILE._02095_ ),
    .Y(\u_cpu.REG_FILE._02096_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06781_  (.A(\u_cpu.REG_FILE._02091_ ),
    .B(\u_cpu.REG_FILE._02096_ ),
    .C(\u_cpu.REG_FILE._01796_ ),
    .Y(\u_cpu.REG_FILE._02097_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06782_  (.A(\u_cpu.REG_FILE.rf[5][18] ),
    .Y(\u_cpu.REG_FILE._02098_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06783_  (.A1(\u_cpu.REG_FILE._01431_ ),
    .A2(\u_cpu.REG_FILE.rf[4][18] ),
    .B1_N(\u_cpu.REG_FILE._01482_ ),
    .Y(\u_cpu.REG_FILE._02099_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._06784_  (.A1(\u_cpu.REG_FILE._02098_ ),
    .A2(\u_cpu.REG_FILE._01850_ ),
    .B1(\u_cpu.REG_FILE._02099_ ),
    .Y(\u_cpu.REG_FILE._02100_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06785_  (.A1(\u_cpu.REG_FILE._01434_ ),
    .A2(\u_cpu.REG_FILE.rf[6][18] ),
    .B1(\u_cpu.REG_FILE._01598_ ),
    .Y(\u_cpu.REG_FILE._02101_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06786_  (.A_N(\u_cpu.REG_FILE.rf[7][18] ),
    .B(\u_cpu.REG_FILE._01906_ ),
    .X(\u_cpu.REG_FILE._02102_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06787_  (.A1(\u_cpu.REG_FILE._02101_ ),
    .A2(\u_cpu.REG_FILE._02102_ ),
    .B1(\u_cpu.REG_FILE._01601_ ),
    .Y(\u_cpu.REG_FILE._02103_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06788_  (.A_N(\u_cpu.REG_FILE.rf[1][18] ),
    .B(\u_cpu.REG_FILE._01804_ ),
    .X(\u_cpu.REG_FILE._02104_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06789_  (.A(\u_cpu.REG_FILE._01076_ ),
    .X(\u_cpu.REG_FILE._02105_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06790_  (.A1(\u_cpu.REG_FILE._02105_ ),
    .A2(\u_cpu.REG_FILE.rf[0][18] ),
    .B1_N(\u_cpu.REG_FILE._01705_ ),
    .Y(\u_cpu.REG_FILE._02106_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06791_  (.A(\u_cpu.REG_FILE.rf[3][18] ),
    .B_N(\u_cpu.REG_FILE._02057_ ),
    .X(\u_cpu.REG_FILE._02107_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06792_  (.A1(\u_cpu.REG_FILE._01707_ ),
    .A2(\u_cpu.REG_FILE.rf[2][18] ),
    .B1(\u_cpu.REG_FILE._02056_ ),
    .C1(\u_cpu.REG_FILE._02107_ ),
    .Y(\u_cpu.REG_FILE._02108_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06793_  (.A1(\u_cpu.REG_FILE._02104_ ),
    .A2(\u_cpu.REG_FILE._02106_ ),
    .B1(\u_cpu.REG_FILE._01858_ ),
    .C1(\u_cpu.REG_FILE._02108_ ),
    .Y(\u_cpu.REG_FILE._02109_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06794_  (.A1(\u_cpu.REG_FILE._02100_ ),
    .A2(\u_cpu.REG_FILE._02103_ ),
    .B1(\u_cpu.REG_FILE._01603_ ),
    .C1(\u_cpu.REG_FILE._02109_ ),
    .Y(\u_cpu.REG_FILE._02110_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._06795_  (.A(\u_cpu.REG_FILE._02097_ ),
    .B(\u_cpu.REG_FILE._02110_ ),
    .Y(\u_cpu.REG_FILE._02111_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06796_  (.A(\u_cpu.REG_FILE.rf[19][18] ),
    .Y(\u_cpu.REG_FILE._02112_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06797_  (.A1(\u_cpu.REG_FILE._01081_ ),
    .A2(\u_cpu.REG_FILE.rf[18][18] ),
    .B1(\u_cpu.REG_FILE._01083_ ),
    .Y(\u_cpu.REG_FILE._02113_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._06798_  (.A1(\u_cpu.REG_FILE._02112_ ),
    .A2(\u_cpu.REG_FILE._01284_ ),
    .B1(\u_cpu.REG_FILE._02113_ ),
    .Y(\u_cpu.REG_FILE._02114_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06799_  (.A(\u_cpu.REG_FILE.rf[17][18] ),
    .Y(\u_cpu.REG_FILE._02115_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06800_  (.A(\u_cpu.REG_FILE._01184_ ),
    .B(\u_cpu.REG_FILE.rf[16][18] ),
    .Y(\u_cpu.REG_FILE._02116_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._06801_  (.A1(\u_cpu.REG_FILE._02115_ ),
    .A2(\u_cpu.REG_FILE._01030_ ),
    .B1(\u_cpu.REG_FILE._01259_ ),
    .C1(\u_cpu.REG_FILE._02116_ ),
    .Y(\u_cpu.REG_FILE._02117_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06802_  (.A(\u_cpu.REG_FILE._01408_ ),
    .B(\u_cpu.REG_FILE.rf[22][18] ),
    .X(\u_cpu.REG_FILE._02118_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06803_  (.A1(\u_cpu.REG_FILE._01327_ ),
    .A2(\u_cpu.REG_FILE.rf[23][18] ),
    .B1(\u_cpu.REG_FILE._01618_ ),
    .C1(\u_cpu.REG_FILE._02118_ ),
    .Y(\u_cpu.REG_FILE._02119_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06804_  (.A1(\u_cpu.REG_FILE._01330_ ),
    .A2(\u_cpu.REG_FILE.rf[20][18] ),
    .B1_N(\u_cpu.REG_FILE._01082_ ),
    .X(\u_cpu.REG_FILE._02120_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06805_  (.A1(\u_cpu.REG_FILE._01329_ ),
    .A2(\u_cpu.REG_FILE.rf[21][18] ),
    .B1(\u_cpu.REG_FILE._02120_ ),
    .Y(\u_cpu.REG_FILE._02121_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06806_  (.A(\u_cpu.REG_FILE._01045_ ),
    .X(\u_cpu.REG_FILE._02122_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06807_  (.A(\u_cpu.REG_FILE._02119_ ),
    .B(\u_cpu.REG_FILE._02121_ ),
    .C(\u_cpu.REG_FILE._02122_ ),
    .Y(\u_cpu.REG_FILE._02123_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._06808_  (.A1(\u_cpu.REG_FILE._01277_ ),
    .A2(\u_cpu.REG_FILE._02114_ ),
    .A3(\u_cpu.REG_FILE._02117_ ),
    .B1(\u_cpu.REG_FILE._02123_ ),
    .C1(\u_cpu.REG_FILE._01090_ ),
    .Y(\u_cpu.REG_FILE._02124_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06809_  (.A(\u_cpu.REG_FILE.rf[27][18] ),
    .B_N(\u_cpu.REG_FILE._01330_ ),
    .X(\u_cpu.REG_FILE._02125_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06810_  (.A1(\u_cpu.REG_FILE._01093_ ),
    .A2(\u_cpu.REG_FILE.rf[26][18] ),
    .B1(\u_cpu.REG_FILE._01099_ ),
    .C1(\u_cpu.REG_FILE._02125_ ),
    .X(\u_cpu.REG_FILE._02126_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06811_  (.A1(\u_cpu.REG_FILE._01774_ ),
    .A2(\u_cpu.REG_FILE.rf[24][18] ),
    .B1_N(\u_cpu.REG_FILE._01553_ ),
    .Y(\u_cpu.REG_FILE._02127_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06812_  (.A_N(\u_cpu.REG_FILE.rf[25][18] ),
    .B(\u_cpu.REG_FILE._01750_ ),
    .X(\u_cpu.REG_FILE._02128_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06813_  (.A1(\u_cpu.REG_FILE._02127_ ),
    .A2(\u_cpu.REG_FILE._02128_ ),
    .B1(\u_cpu.REG_FILE._01814_ ),
    .Y(\u_cpu.REG_FILE._02129_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06814_  (.A(\u_cpu.REG_FILE._01325_ ),
    .B(\u_cpu.REG_FILE.rf[30][18] ),
    .Y(\u_cpu.REG_FILE._02130_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06815_  (.A1(\u_cpu.REG_FILE.rf[31][18] ),
    .A2(\u_cpu.REG_FILE._01329_ ),
    .B1(\u_cpu.REG_FILE._01099_ ),
    .Y(\u_cpu.REG_FILE._02131_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06816_  (.A1(\u_cpu.REG_FILE._01345_ ),
    .A2(\u_cpu.REG_FILE.rf[28][18] ),
    .B1_N(\u_cpu.REG_FILE._01082_ ),
    .X(\u_cpu.REG_FILE._02132_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06817_  (.A1(\u_cpu.REG_FILE._01265_ ),
    .A2(\u_cpu.REG_FILE.rf[29][18] ),
    .B1(\u_cpu.REG_FILE._02132_ ),
    .Y(\u_cpu.REG_FILE._02133_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06818_  (.A1(\u_cpu.REG_FILE._02130_ ),
    .A2(\u_cpu.REG_FILE._02131_ ),
    .B1(\u_cpu.REG_FILE._02133_ ),
    .C1(\u_cpu.REG_FILE._01333_ ),
    .Y(\u_cpu.REG_FILE._02134_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06819_  (.A1(\u_cpu.REG_FILE._02126_ ),
    .A2(\u_cpu.REG_FILE._02129_ ),
    .B1(\u_cpu.REG_FILE._01069_ ),
    .C1(\u_cpu.REG_FILE._02134_ ),
    .Y(\u_cpu.REG_FILE._02135_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06820_  (.A(\u_cpu.REG_FILE._02124_ ),
    .B(\u_cpu.REG_FILE._01025_ ),
    .C(\u_cpu.REG_FILE._02135_ ),
    .Y(\u_cpu.REG_FILE._02136_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06821_  (.A1(\u_cpu.REG_FILE._01888_ ),
    .A2(\u_cpu.REG_FILE._02111_ ),
    .B1(\u_cpu.REG_FILE._02136_ ),
    .C1(\u_cpu.REG_FILE._01737_ ),
    .X(\u_cpu.ALU.SrcA[18] ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06822_  (.A1(\u_cpu.REG_FILE._01184_ ),
    .A2(\u_cpu.REG_FILE.rf[8][19] ),
    .B1_N(\u_cpu.REG_FILE._01521_ ),
    .Y(\u_cpu.REG_FILE._02137_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06823_  (.A_N(\u_cpu.REG_FILE.rf[9][19] ),
    .B(\u_cpu.REG_FILE._01074_ ),
    .X(\u_cpu.REG_FILE._02138_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06824_  (.A1(\u_cpu.REG_FILE._02137_ ),
    .A2(\u_cpu.REG_FILE._02138_ ),
    .B1(\u_cpu.REG_FILE._01525_ ),
    .Y(\u_cpu.REG_FILE._02139_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06825_  (.A(\u_cpu.REG_FILE._01528_ ),
    .B(\u_cpu.REG_FILE.rf[10][19] ),
    .X(\u_cpu.REG_FILE._02140_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06826_  (.A1(\u_cpu.REG_FILE._01137_ ),
    .A2(\u_cpu.REG_FILE.rf[11][19] ),
    .B1(\u_cpu.REG_FILE._01387_ ),
    .C1(\u_cpu.REG_FILE._02140_ ),
    .X(\u_cpu.REG_FILE._02141_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06827_  (.A(\u_cpu.REG_FILE._01118_ ),
    .B(\u_cpu.REG_FILE.rf[12][19] ),
    .Y(\u_cpu.REG_FILE._02142_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06828_  (.A1(\u_cpu.REG_FILE.rf[13][19] ),
    .A2(\u_cpu.REG_FILE._01287_ ),
    .B1_N(\u_cpu.REG_FILE._01305_ ),
    .Y(\u_cpu.REG_FILE._02143_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06829_  (.A(\u_cpu.REG_FILE._01536_ ),
    .B(\u_cpu.REG_FILE.rf[14][19] ),
    .X(\u_cpu.REG_FILE._02144_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06830_  (.A1(\u_cpu.REG_FILE._01535_ ),
    .A2(\u_cpu.REG_FILE.rf[15][19] ),
    .B1(\u_cpu.REG_FILE._01527_ ),
    .C1(\u_cpu.REG_FILE._02144_ ),
    .Y(\u_cpu.REG_FILE._02145_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06831_  (.A1(\u_cpu.REG_FILE._02142_ ),
    .A2(\u_cpu.REG_FILE._02143_ ),
    .B1(\u_cpu.REG_FILE._01129_ ),
    .C1(\u_cpu.REG_FILE._02145_ ),
    .Y(\u_cpu.REG_FILE._02146_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06832_  (.A1(\u_cpu.REG_FILE._02139_ ),
    .A2(\u_cpu.REG_FILE._02141_ ),
    .B1(\u_cpu.REG_FILE._01117_ ),
    .C1(\u_cpu.REG_FILE._02146_ ),
    .X(\u_cpu.REG_FILE._02147_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06833_  (.A_N(\u_cpu.REG_FILE.rf[1][19] ),
    .B(\u_cpu.REG_FILE._01547_ ),
    .X(\u_cpu.REG_FILE._02148_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06834_  (.A1(\u_cpu.REG_FILE._01093_ ),
    .A2(\u_cpu.REG_FILE.rf[0][19] ),
    .B1_N(\u_cpu.REG_FILE._01550_ ),
    .Y(\u_cpu.REG_FILE._02149_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06835_  (.A(\u_cpu.REG_FILE.rf[3][19] ),
    .B_N(\u_cpu.REG_FILE._01310_ ),
    .X(\u_cpu.REG_FILE._02150_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06836_  (.A1(\u_cpu.REG_FILE._01308_ ),
    .A2(\u_cpu.REG_FILE.rf[2][19] ),
    .B1(\u_cpu.REG_FILE._01309_ ),
    .C1(\u_cpu.REG_FILE._02150_ ),
    .Y(\u_cpu.REG_FILE._02151_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06837_  (.A1(\u_cpu.REG_FILE._02148_ ),
    .A2(\u_cpu.REG_FILE._02149_ ),
    .B1(\u_cpu.REG_FILE._01059_ ),
    .C1(\u_cpu.REG_FILE._02151_ ),
    .Y(\u_cpu.REG_FILE._02152_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06838_  (.A_N(\u_cpu.REG_FILE.rf[5][19] ),
    .B(\u_cpu.REG_FILE._01547_ ),
    .X(\u_cpu.REG_FILE._02153_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06839_  (.A1(\u_cpu.REG_FILE._01549_ ),
    .A2(\u_cpu.REG_FILE.rf[4][19] ),
    .B1_N(\u_cpu.REG_FILE._01550_ ),
    .Y(\u_cpu.REG_FILE._02154_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.REG_FILE._06840_  (.A1(\u_cpu.REG_FILE._01262_ ),
    .A2(\u_cpu.REG_FILE.rf[6][19] ),
    .B1(\u_cpu.REG_FILE._01553_ ),
    .X(\u_cpu.REG_FILE._02155_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06841_  (.A1(\u_cpu.REG_FILE.rf[7][19] ),
    .A2(\u_cpu.REG_FILE._01287_ ),
    .B1(\u_cpu.REG_FILE._02155_ ),
    .Y(\u_cpu.REG_FILE._02156_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06842_  (.A1(\u_cpu.REG_FILE._02153_ ),
    .A2(\u_cpu.REG_FILE._02154_ ),
    .B1(\u_cpu.REG_FILE._01087_ ),
    .C1(\u_cpu.REG_FILE._02156_ ),
    .Y(\u_cpu.REG_FILE._02157_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._06843_  (.A1(\u_cpu.REG_FILE._01541_ ),
    .A2(\u_cpu.REG_FILE._02152_ ),
    .A3(\u_cpu.REG_FILE._02157_ ),
    .B1(\u_cpu.REG_FILE._01024_ ),
    .X(\u_cpu.REG_FILE._02158_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06844_  (.A1(\u_cpu.REG_FILE._01279_ ),
    .A2(\u_cpu.REG_FILE.rf[18][19] ),
    .B1(\u_cpu.REG_FILE._01280_ ),
    .Y(\u_cpu.REG_FILE._02159_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06845_  (.A(\u_cpu.REG_FILE.rf[19][19] ),
    .B(\u_cpu.REG_FILE._01298_ ),
    .Y(\u_cpu.REG_FILE._02160_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06846_  (.A1(\u_cpu.REG_FILE._01029_ ),
    .A2(\u_cpu.REG_FILE.rf[16][19] ),
    .B1_N(\u_cpu.REG_FILE._01239_ ),
    .X(\u_cpu.REG_FILE._02161_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06847_  (.A1(\u_cpu.REG_FILE._01137_ ),
    .A2(\u_cpu.REG_FILE.rf[17][19] ),
    .B1(\u_cpu.REG_FILE._02161_ ),
    .Y(\u_cpu.REG_FILE._02162_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06848_  (.A1(\u_cpu.REG_FILE._02159_ ),
    .A2(\u_cpu.REG_FILE._02160_ ),
    .B1(\u_cpu.REG_FILE._01307_ ),
    .C1(\u_cpu.REG_FILE._02162_ ),
    .Y(\u_cpu.REG_FILE._02163_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06849_  (.A(\u_cpu.REG_FILE._02010_ ),
    .B(\u_cpu.REG_FILE.rf[22][19] ),
    .Y(\u_cpu.REG_FILE._02164_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06850_  (.A1(\u_cpu.REG_FILE.rf[23][19] ),
    .A2(\u_cpu.REG_FILE._01146_ ),
    .B1(\u_cpu.REG_FILE._01660_ ),
    .Y(\u_cpu.REG_FILE._02165_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06851_  (.A1(\u_cpu.REG_FILE._02013_ ),
    .A2(\u_cpu.REG_FILE.rf[20][19] ),
    .B1_N(\u_cpu.REG_FILE._01142_ ),
    .X(\u_cpu.REG_FILE._02166_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06852_  (.A1(\u_cpu.REG_FILE._01140_ ),
    .A2(\u_cpu.REG_FILE.rf[21][19] ),
    .B1(\u_cpu.REG_FILE._02166_ ),
    .Y(\u_cpu.REG_FILE._02167_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06853_  (.A1(\u_cpu.REG_FILE._02164_ ),
    .A2(\u_cpu.REG_FILE._02165_ ),
    .B1(\u_cpu.REG_FILE._02167_ ),
    .C1(\u_cpu.REG_FILE._02016_ ),
    .Y(\u_cpu.REG_FILE._02168_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06854_  (.A(\u_cpu.REG_FILE._01132_ ),
    .B(\u_cpu.REG_FILE._02163_ ),
    .C(\u_cpu.REG_FILE._02168_ ),
    .Y(\u_cpu.REG_FILE._02169_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06855_  (.A(\u_cpu.REG_FILE.rf[27][19] ),
    .B_N(\u_cpu.REG_FILE._01330_ ),
    .X(\u_cpu.REG_FILE._02170_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06856_  (.A1(\u_cpu.REG_FILE._01093_ ),
    .A2(\u_cpu.REG_FILE.rf[26][19] ),
    .B1(\u_cpu.REG_FILE._01099_ ),
    .C1(\u_cpu.REG_FILE._02170_ ),
    .X(\u_cpu.REG_FILE._02171_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06857_  (.A1(\u_cpu.REG_FILE._01404_ ),
    .A2(\u_cpu.REG_FILE.rf[24][19] ),
    .B1_N(\u_cpu.REG_FILE._01553_ ),
    .Y(\u_cpu.REG_FILE._02172_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06858_  (.A_N(\u_cpu.REG_FILE.rf[25][19] ),
    .B(\u_cpu.REG_FILE._01750_ ),
    .X(\u_cpu.REG_FILE._02173_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06859_  (.A1(\u_cpu.REG_FILE._02172_ ),
    .A2(\u_cpu.REG_FILE._02173_ ),
    .B1(\u_cpu.REG_FILE._01814_ ),
    .Y(\u_cpu.REG_FILE._02174_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06860_  (.A(\u_cpu.REG_FILE._01325_ ),
    .B(\u_cpu.REG_FILE.rf[30][19] ),
    .Y(\u_cpu.REG_FILE._02175_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06861_  (.A1(\u_cpu.REG_FILE.rf[31][19] ),
    .A2(\u_cpu.REG_FILE._01327_ ),
    .B1(\u_cpu.REG_FILE._01099_ ),
    .Y(\u_cpu.REG_FILE._02176_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06862_  (.A1(\u_cpu.REG_FILE._01330_ ),
    .A2(\u_cpu.REG_FILE.rf[28][19] ),
    .B1_N(\u_cpu.REG_FILE._01082_ ),
    .X(\u_cpu.REG_FILE._02177_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06863_  (.A1(\u_cpu.REG_FILE._01265_ ),
    .A2(\u_cpu.REG_FILE.rf[29][19] ),
    .B1(\u_cpu.REG_FILE._02177_ ),
    .Y(\u_cpu.REG_FILE._02178_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06864_  (.A1(\u_cpu.REG_FILE._02175_ ),
    .A2(\u_cpu.REG_FILE._02176_ ),
    .B1(\u_cpu.REG_FILE._02178_ ),
    .C1(\u_cpu.REG_FILE._01333_ ),
    .Y(\u_cpu.REG_FILE._02179_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06865_  (.A1(\u_cpu.REG_FILE._02171_ ),
    .A2(\u_cpu.REG_FILE._02174_ ),
    .B1(\u_cpu.REG_FILE._01069_ ),
    .C1(\u_cpu.REG_FILE._02179_ ),
    .Y(\u_cpu.REG_FILE._02180_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06866_  (.A(\u_cpu.REG_FILE._02169_ ),
    .B(\u_cpu.REG_FILE._01025_ ),
    .C(\u_cpu.REG_FILE._02180_ ),
    .Y(\u_cpu.REG_FILE._02181_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06867_  (.A1(\u_cpu.REG_FILE._02147_ ),
    .A2(\u_cpu.REG_FILE._02158_ ),
    .B1(\u_cpu.REG_FILE._02181_ ),
    .C1(\u_cpu.REG_FILE._01737_ ),
    .X(\u_cpu.ALU.SrcA[19] ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06868_  (.A(\u_cpu.REG_FILE._01279_ ),
    .B(\u_cpu.REG_FILE.rf[22][20] ),
    .X(\u_cpu.REG_FILE._02182_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06869_  (.A1(\u_cpu.REG_FILE._01039_ ),
    .A2(\u_cpu.REG_FILE.rf[23][20] ),
    .B1(\u_cpu.REG_FILE._01259_ ),
    .C1(\u_cpu.REG_FILE._02182_ ),
    .Y(\u_cpu.REG_FILE._02183_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06870_  (.A1(\u_cpu.REG_FILE._01279_ ),
    .A2(\u_cpu.REG_FILE.rf[20][20] ),
    .B1_N(\u_cpu.REG_FILE._01533_ ),
    .X(\u_cpu.REG_FILE._02184_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06871_  (.A(\u_cpu.REG_FILE.rf[21][20] ),
    .B_N(\u_cpu.REG_FILE._01260_ ),
    .X(\u_cpu.REG_FILE._02185_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._06872_  (.A1(\u_cpu.REG_FILE._02184_ ),
    .A2(\u_cpu.REG_FILE._02185_ ),
    .B1(\u_cpu.REG_FILE._01525_ ),
    .Y(\u_cpu.REG_FILE._02186_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06873_  (.A1(\u_cpu.REG_FILE._01133_ ),
    .A2(\u_cpu.REG_FILE.rf[16][20] ),
    .B1_N(\u_cpu.REG_FILE._01380_ ),
    .Y(\u_cpu.REG_FILE._02187_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06874_  (.A_N(\u_cpu.REG_FILE.rf[17][20] ),
    .B(\u_cpu.REG_FILE._01161_ ),
    .X(\u_cpu.REG_FILE._02188_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06875_  (.A1(\u_cpu.REG_FILE._01279_ ),
    .A2(\u_cpu.REG_FILE.rf[18][20] ),
    .B1(\u_cpu.REG_FILE._01280_ ),
    .Y(\u_cpu.REG_FILE._02189_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06876_  (.A_N(\u_cpu.REG_FILE.rf[19][20] ),
    .B(\u_cpu.REG_FILE._01382_ ),
    .X(\u_cpu.REG_FILE._02190_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.REG_FILE._06877_  (.A1(\u_cpu.REG_FILE._02187_ ),
    .A2(\u_cpu.REG_FILE._02188_ ),
    .B1(\u_cpu.REG_FILE._02189_ ),
    .B2(\u_cpu.REG_FILE._02190_ ),
    .C1(\u_cpu.REG_FILE._01307_ ),
    .X(\u_cpu.REG_FILE._02191_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._06878_  (.A1(\u_cpu.REG_FILE._02183_ ),
    .A2(\u_cpu.REG_FILE._02186_ ),
    .B1(\u_cpu.REG_FILE._01070_ ),
    .C1(\u_cpu.REG_FILE._02191_ ),
    .Y(\u_cpu.REG_FILE._02192_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06879_  (.A(\u_cpu.REG_FILE.rf[31][20] ),
    .B_N(\u_cpu.REG_FILE._01111_ ),
    .X(\u_cpu.REG_FILE._02193_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06880_  (.A1(\u_cpu.REG_FILE._01030_ ),
    .A2(\u_cpu.REG_FILE.rf[30][20] ),
    .B1(\u_cpu.REG_FILE._01033_ ),
    .C1(\u_cpu.REG_FILE._02193_ ),
    .Y(\u_cpu.REG_FILE._02194_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06881_  (.A1(\u_cpu.REG_FILE._01299_ ),
    .A2(\u_cpu.REG_FILE.rf[28][20] ),
    .B1_N(\u_cpu.REG_FILE._01106_ ),
    .X(\u_cpu.REG_FILE._02195_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06882_  (.A1(\u_cpu.REG_FILE._01298_ ),
    .A2(\u_cpu.REG_FILE.rf[29][20] ),
    .B1(\u_cpu.REG_FILE._02195_ ),
    .Y(\u_cpu.REG_FILE._02196_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06883_  (.A(\u_cpu.REG_FILE._02194_ ),
    .B(\u_cpu.REG_FILE._02196_ ),
    .C(\u_cpu.REG_FILE._01293_ ),
    .Y(\u_cpu.REG_FILE._02197_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06884_  (.A_N(\u_cpu.REG_FILE.rf[25][20] ),
    .B(\u_cpu.REG_FILE._01547_ ),
    .X(\u_cpu.REG_FILE._02198_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06885_  (.A1(\u_cpu.REG_FILE._01549_ ),
    .A2(\u_cpu.REG_FILE.rf[24][20] ),
    .B1_N(\u_cpu.REG_FILE._01550_ ),
    .Y(\u_cpu.REG_FILE._02199_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06886_  (.A(\u_cpu.REG_FILE.rf[27][20] ),
    .B_N(\u_cpu.REG_FILE._01310_ ),
    .X(\u_cpu.REG_FILE._02200_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06887_  (.A1(\u_cpu.REG_FILE._01308_ ),
    .A2(\u_cpu.REG_FILE.rf[26][20] ),
    .B1(\u_cpu.REG_FILE._01309_ ),
    .C1(\u_cpu.REG_FILE._02200_ ),
    .Y(\u_cpu.REG_FILE._02201_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06888_  (.A1(\u_cpu.REG_FILE._02198_ ),
    .A2(\u_cpu.REG_FILE._02199_ ),
    .B1(\u_cpu.REG_FILE._01059_ ),
    .C1(\u_cpu.REG_FILE._02201_ ),
    .Y(\u_cpu.REG_FILE._02202_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._06889_  (.A1(\u_cpu.REG_FILE._02197_ ),
    .A2(\u_cpu.REG_FILE._02202_ ),
    .A3(\u_cpu.REG_FILE._01314_ ),
    .B1(\u_cpu.REG_FILE._01315_ ),
    .X(\u_cpu.REG_FILE._02203_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06890_  (.A(\u_cpu.REG_FILE._02010_ ),
    .B(\u_cpu.REG_FILE.rf[14][20] ),
    .Y(\u_cpu.REG_FILE._02204_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06891_  (.A1(\u_cpu.REG_FILE.rf[15][20] ),
    .A2(\u_cpu.REG_FILE._01146_ ),
    .B1(\u_cpu.REG_FILE._01660_ ),
    .Y(\u_cpu.REG_FILE._02205_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06892_  (.A1(\u_cpu.REG_FILE._02013_ ),
    .A2(\u_cpu.REG_FILE.rf[12][20] ),
    .B1_N(\u_cpu.REG_FILE._01142_ ),
    .X(\u_cpu.REG_FILE._02206_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06893_  (.A1(\u_cpu.REG_FILE._01140_ ),
    .A2(\u_cpu.REG_FILE.rf[13][20] ),
    .B1(\u_cpu.REG_FILE._02206_ ),
    .Y(\u_cpu.REG_FILE._02207_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06894_  (.A1(\u_cpu.REG_FILE._02204_ ),
    .A2(\u_cpu.REG_FILE._02205_ ),
    .B1(\u_cpu.REG_FILE._02207_ ),
    .C1(\u_cpu.REG_FILE._02016_ ),
    .Y(\u_cpu.REG_FILE._02208_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06895_  (.A(\u_cpu.REG_FILE.rf[11][20] ),
    .B_N(\u_cpu.REG_FILE._01148_ ),
    .X(\u_cpu.REG_FILE._02209_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06896_  (.A1(\u_cpu.REG_FILE._01279_ ),
    .A2(\u_cpu.REG_FILE.rf[10][20] ),
    .B1(\u_cpu.REG_FILE._01618_ ),
    .C1(\u_cpu.REG_FILE._02209_ ),
    .Y(\u_cpu.REG_FILE._02210_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06897_  (.A1(\u_cpu.REG_FILE._01536_ ),
    .A2(\u_cpu.REG_FILE.rf[8][20] ),
    .B1_N(\u_cpu.REG_FILE._01134_ ),
    .X(\u_cpu.REG_FILE._02211_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06898_  (.A1(\u_cpu.REG_FILE._01120_ ),
    .A2(\u_cpu.REG_FILE.rf[9][20] ),
    .B1(\u_cpu.REG_FILE._02211_ ),
    .Y(\u_cpu.REG_FILE._02212_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06899_  (.A(\u_cpu.REG_FILE._01307_ ),
    .B(\u_cpu.REG_FILE._02210_ ),
    .C(\u_cpu.REG_FILE._02212_ ),
    .Y(\u_cpu.REG_FILE._02213_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06900_  (.A(\u_cpu.REG_FILE._02208_ ),
    .B(\u_cpu.REG_FILE._02213_ ),
    .C(\u_cpu.REG_FILE._01314_ ),
    .Y(\u_cpu.REG_FILE._02214_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06901_  (.A(\u_cpu.REG_FILE.rf[3][20] ),
    .B_N(\u_cpu.REG_FILE._01148_ ),
    .X(\u_cpu.REG_FILE._02215_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06902_  (.A1(\u_cpu.REG_FILE._02018_ ),
    .A2(\u_cpu.REG_FILE.rf[2][20] ),
    .B1(\u_cpu.REG_FILE._01618_ ),
    .C1(\u_cpu.REG_FILE._02215_ ),
    .Y(\u_cpu.REG_FILE._02216_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06903_  (.A1(\u_cpu.REG_FILE._01152_ ),
    .A2(\u_cpu.REG_FILE.rf[0][20] ),
    .B1_N(\u_cpu.REG_FILE._01153_ ),
    .X(\u_cpu.REG_FILE._02217_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06904_  (.A1(\u_cpu.REG_FILE._01726_ ),
    .A2(\u_cpu.REG_FILE.rf[1][20] ),
    .B1(\u_cpu.REG_FILE._02217_ ),
    .Y(\u_cpu.REG_FILE._02218_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06905_  (.A(\u_cpu.REG_FILE._01525_ ),
    .B(\u_cpu.REG_FILE._02216_ ),
    .C(\u_cpu.REG_FILE._02218_ ),
    .Y(\u_cpu.REG_FILE._02219_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06906_  (.A1(\u_cpu.REG_FILE._01029_ ),
    .A2(\u_cpu.REG_FILE.rf[4][20] ),
    .B1_N(\u_cpu.REG_FILE._01239_ ),
    .X(\u_cpu.REG_FILE._02220_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06907_  (.A1(\u_cpu.REG_FILE._01137_ ),
    .A2(\u_cpu.REG_FILE.rf[5][20] ),
    .B1(\u_cpu.REG_FILE._02220_ ),
    .Y(\u_cpu.REG_FILE._02221_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.REG_FILE._06908_  (.A1(\u_cpu.REG_FILE._02013_ ),
    .A2(\u_cpu.REG_FILE.rf[6][20] ),
    .B1(\u_cpu.REG_FILE._01032_ ),
    .X(\u_cpu.REG_FILE._02222_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06909_  (.A1(\u_cpu.REG_FILE.rf[7][20] ),
    .A2(\u_cpu.REG_FILE._01386_ ),
    .B1(\u_cpu.REG_FILE._02222_ ),
    .Y(\u_cpu.REG_FILE._02223_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06910_  (.A(\u_cpu.REG_FILE._02221_ ),
    .B(\u_cpu.REG_FILE._01156_ ),
    .C(\u_cpu.REG_FILE._02223_ ),
    .Y(\u_cpu.REG_FILE._02224_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06911_  (.A(\u_cpu.REG_FILE._01132_ ),
    .B(\u_cpu.REG_FILE._02219_ ),
    .C(\u_cpu.REG_FILE._02224_ ),
    .Y(\u_cpu.REG_FILE._02225_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06912_  (.A(\u_cpu.REG_FILE._01315_ ),
    .B(\u_cpu.REG_FILE._02214_ ),
    .C(\u_cpu.REG_FILE._02225_ ),
    .Y(\u_cpu.REG_FILE._02226_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._06913_  (.A(\u_cpu.REG_FILE._01164_ ),
    .X(\u_cpu.REG_FILE._02227_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06914_  (.A1(\u_cpu.REG_FILE._02192_ ),
    .A2(\u_cpu.REG_FILE._02203_ ),
    .B1(\u_cpu.REG_FILE._02226_ ),
    .C1(\u_cpu.REG_FILE._02227_ ),
    .X(\u_cpu.ALU.SrcA[20] ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06915_  (.A1(\u_cpu.REG_FILE._01184_ ),
    .A2(\u_cpu.REG_FILE.rf[8][21] ),
    .B1_N(\u_cpu.REG_FILE._01094_ ),
    .Y(\u_cpu.REG_FILE._02228_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06916_  (.A_N(\u_cpu.REG_FILE.rf[9][21] ),
    .B(\u_cpu.REG_FILE._01074_ ),
    .X(\u_cpu.REG_FILE._02229_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06917_  (.A1(\u_cpu.REG_FILE._02228_ ),
    .A2(\u_cpu.REG_FILE._02229_ ),
    .B1(\u_cpu.REG_FILE._01525_ ),
    .Y(\u_cpu.REG_FILE._02230_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06918_  (.A(\u_cpu.REG_FILE._01528_ ),
    .B(\u_cpu.REG_FILE.rf[10][21] ),
    .X(\u_cpu.REG_FILE._02231_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06919_  (.A1(\u_cpu.REG_FILE._01137_ ),
    .A2(\u_cpu.REG_FILE.rf[11][21] ),
    .B1(\u_cpu.REG_FILE._01387_ ),
    .C1(\u_cpu.REG_FILE._02231_ ),
    .X(\u_cpu.REG_FILE._02232_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06920_  (.A(\u_cpu.REG_FILE._01118_ ),
    .B(\u_cpu.REG_FILE.rf[12][21] ),
    .Y(\u_cpu.REG_FILE._02233_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06921_  (.A1(\u_cpu.REG_FILE.rf[13][21] ),
    .A2(\u_cpu.REG_FILE._01535_ ),
    .B1_N(\u_cpu.REG_FILE._01305_ ),
    .Y(\u_cpu.REG_FILE._02234_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06922_  (.A(\u_cpu.REG_FILE._01536_ ),
    .B(\u_cpu.REG_FILE.rf[14][21] ),
    .X(\u_cpu.REG_FILE._02235_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06923_  (.A1(\u_cpu.REG_FILE._01535_ ),
    .A2(\u_cpu.REG_FILE.rf[15][21] ),
    .B1(\u_cpu.REG_FILE._01527_ ),
    .C1(\u_cpu.REG_FILE._02235_ ),
    .Y(\u_cpu.REG_FILE._02236_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06924_  (.A1(\u_cpu.REG_FILE._02233_ ),
    .A2(\u_cpu.REG_FILE._02234_ ),
    .B1(\u_cpu.REG_FILE._01129_ ),
    .C1(\u_cpu.REG_FILE._02236_ ),
    .Y(\u_cpu.REG_FILE._02237_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06925_  (.A1(\u_cpu.REG_FILE._02230_ ),
    .A2(\u_cpu.REG_FILE._02232_ ),
    .B1(\u_cpu.REG_FILE._01117_ ),
    .C1(\u_cpu.REG_FILE._02237_ ),
    .X(\u_cpu.REG_FILE._02238_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06926_  (.A_N(\u_cpu.REG_FILE.rf[1][21] ),
    .B(\u_cpu.REG_FILE._01547_ ),
    .X(\u_cpu.REG_FILE._02239_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06927_  (.A1(\u_cpu.REG_FILE._01549_ ),
    .A2(\u_cpu.REG_FILE.rf[0][21] ),
    .B1_N(\u_cpu.REG_FILE._01550_ ),
    .Y(\u_cpu.REG_FILE._02240_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06928_  (.A(\u_cpu.REG_FILE.rf[3][21] ),
    .B_N(\u_cpu.REG_FILE._01310_ ),
    .X(\u_cpu.REG_FILE._02241_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06929_  (.A1(\u_cpu.REG_FILE._01061_ ),
    .A2(\u_cpu.REG_FILE.rf[2][21] ),
    .B1(\u_cpu.REG_FILE._01309_ ),
    .C1(\u_cpu.REG_FILE._02241_ ),
    .Y(\u_cpu.REG_FILE._02242_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06930_  (.A1(\u_cpu.REG_FILE._02239_ ),
    .A2(\u_cpu.REG_FILE._02240_ ),
    .B1(\u_cpu.REG_FILE._01059_ ),
    .C1(\u_cpu.REG_FILE._02242_ ),
    .Y(\u_cpu.REG_FILE._02243_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06931_  (.A1(\u_cpu.REG_FILE._01161_ ),
    .A2(\u_cpu.REG_FILE.rf[4][21] ),
    .B1_N(\u_cpu.REG_FILE._01042_ ),
    .X(\u_cpu.REG_FILE._02244_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06932_  (.A1(\u_cpu.REG_FILE._01039_ ),
    .A2(\u_cpu.REG_FILE.rf[5][21] ),
    .B1(\u_cpu.REG_FILE._02244_ ),
    .Y(\u_cpu.REG_FILE._02245_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.REG_FILE._06933_  (.A1(\u_cpu.REG_FILE._01029_ ),
    .A2(\u_cpu.REG_FILE.rf[6][21] ),
    .B1(\u_cpu.REG_FILE._01258_ ),
    .X(\u_cpu.REG_FILE._02246_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06934_  (.A1(\u_cpu.REG_FILE.rf[7][21] ),
    .A2(\u_cpu.REG_FILE._01287_ ),
    .B1(\u_cpu.REG_FILE._02246_ ),
    .Y(\u_cpu.REG_FILE._02247_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06935_  (.A(\u_cpu.REG_FILE._02245_ ),
    .B(\u_cpu.REG_FILE._02247_ ),
    .C(\u_cpu.REG_FILE._02016_ ),
    .Y(\u_cpu.REG_FILE._02248_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._06936_  (.A1(\u_cpu.REG_FILE._01541_ ),
    .A2(\u_cpu.REG_FILE._02243_ ),
    .A3(\u_cpu.REG_FILE._02248_ ),
    .B1(\u_cpu.REG_FILE._01024_ ),
    .X(\u_cpu.REG_FILE._02249_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06937_  (.A(\u_cpu.REG_FILE.rf[19][21] ),
    .Y(\u_cpu.REG_FILE._02250_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06938_  (.A1(\u_cpu.REG_FILE._01081_ ),
    .A2(\u_cpu.REG_FILE.rf[18][21] ),
    .B1(\u_cpu.REG_FILE._01083_ ),
    .Y(\u_cpu.REG_FILE._02251_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._06939_  (.A1(\u_cpu.REG_FILE._02250_ ),
    .A2(\u_cpu.REG_FILE._01284_ ),
    .B1(\u_cpu.REG_FILE._02251_ ),
    .Y(\u_cpu.REG_FILE._02252_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06940_  (.A(\u_cpu.REG_FILE.rf[17][21] ),
    .Y(\u_cpu.REG_FILE._02253_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06941_  (.A(\u_cpu.REG_FILE._01184_ ),
    .B(\u_cpu.REG_FILE.rf[16][21] ),
    .Y(\u_cpu.REG_FILE._02254_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._06942_  (.A1(\u_cpu.REG_FILE._02253_ ),
    .A2(\u_cpu.REG_FILE._01030_ ),
    .B1(\u_cpu.REG_FILE._01259_ ),
    .C1(\u_cpu.REG_FILE._02254_ ),
    .Y(\u_cpu.REG_FILE._02255_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06943_  (.A(\u_cpu.REG_FILE._01317_ ),
    .B(\u_cpu.REG_FILE.rf[20][21] ),
    .Y(\u_cpu.REG_FILE._02256_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06944_  (.A_N(\u_cpu.REG_FILE.rf[21][21] ),
    .B(\u_cpu.REG_FILE._02013_ ),
    .X(\u_cpu.REG_FILE._02257_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06945_  (.A(\u_cpu.REG_FILE.rf[23][21] ),
    .B_N(\u_cpu.REG_FILE._01049_ ),
    .X(\u_cpu.REG_FILE._02258_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06946_  (.A1(\u_cpu.REG_FILE._01317_ ),
    .A2(\u_cpu.REG_FILE.rf[22][21] ),
    .B1(\u_cpu.REG_FILE._01533_ ),
    .C1(\u_cpu.REG_FILE._02258_ ),
    .Y(\u_cpu.REG_FILE._02259_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._06947_  (.A1(\u_cpu.REG_FILE._01387_ ),
    .A2(\u_cpu.REG_FILE._02256_ ),
    .A3(\u_cpu.REG_FILE._02257_ ),
    .B1(\u_cpu.REG_FILE._01115_ ),
    .C1(\u_cpu.REG_FILE._02259_ ),
    .Y(\u_cpu.REG_FILE._02260_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._06948_  (.A1(\u_cpu.REG_FILE._01277_ ),
    .A2(\u_cpu.REG_FILE._02252_ ),
    .A3(\u_cpu.REG_FILE._02255_ ),
    .B1(\u_cpu.REG_FILE._02260_ ),
    .C1(\u_cpu.REG_FILE._01090_ ),
    .Y(\u_cpu.REG_FILE._02261_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06949_  (.A(\u_cpu.REG_FILE._02010_ ),
    .B(\u_cpu.REG_FILE.rf[24][21] ),
    .Y(\u_cpu.REG_FILE._02262_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06950_  (.A1(\u_cpu.REG_FILE.rf[25][21] ),
    .A2(\u_cpu.REG_FILE._01151_ ),
    .B1_N(\u_cpu.REG_FILE._01305_ ),
    .Y(\u_cpu.REG_FILE._02263_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06951_  (.A(\u_cpu.REG_FILE._01148_ ),
    .B(\u_cpu.REG_FILE.rf[26][21] ),
    .X(\u_cpu.REG_FILE._02264_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06952_  (.A1(\u_cpu.REG_FILE._01969_ ),
    .A2(\u_cpu.REG_FILE.rf[27][21] ),
    .B1(\u_cpu.REG_FILE._01309_ ),
    .C1(\u_cpu.REG_FILE._02264_ ),
    .Y(\u_cpu.REG_FILE._02265_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06953_  (.A1(\u_cpu.REG_FILE._02262_ ),
    .A2(\u_cpu.REG_FILE._02263_ ),
    .B1(\u_cpu.REG_FILE._01307_ ),
    .C1(\u_cpu.REG_FILE._02265_ ),
    .Y(\u_cpu.REG_FILE._02266_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06954_  (.A(\u_cpu.REG_FILE.rf[31][21] ),
    .B_N(\u_cpu.REG_FILE._01065_ ),
    .X(\u_cpu.REG_FILE._02267_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06955_  (.A1(\u_cpu.REG_FILE._01061_ ),
    .A2(\u_cpu.REG_FILE.rf[30][21] ),
    .B1(\u_cpu.REG_FILE._01147_ ),
    .C1(\u_cpu.REG_FILE._02267_ ),
    .Y(\u_cpu.REG_FILE._02268_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06956_  (.A1(\u_cpu.REG_FILE._01152_ ),
    .A2(\u_cpu.REG_FILE.rf[28][21] ),
    .B1_N(\u_cpu.REG_FILE._01153_ ),
    .X(\u_cpu.REG_FILE._02269_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06957_  (.A1(\u_cpu.REG_FILE._01726_ ),
    .A2(\u_cpu.REG_FILE.rf[29][21] ),
    .B1(\u_cpu.REG_FILE._02269_ ),
    .Y(\u_cpu.REG_FILE._02270_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06958_  (.A(\u_cpu.REG_FILE._02268_ ),
    .B(\u_cpu.REG_FILE._02270_ ),
    .C(\u_cpu.REG_FILE._01156_ ),
    .Y(\u_cpu.REG_FILE._02271_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06959_  (.A(\u_cpu.REG_FILE._02266_ ),
    .B(\u_cpu.REG_FILE._01314_ ),
    .C(\u_cpu.REG_FILE._02271_ ),
    .Y(\u_cpu.REG_FILE._02272_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06960_  (.A(\u_cpu.REG_FILE._02261_ ),
    .B(\u_cpu.REG_FILE._01025_ ),
    .C(\u_cpu.REG_FILE._02272_ ),
    .Y(\u_cpu.REG_FILE._02273_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06961_  (.A1(\u_cpu.REG_FILE._02238_ ),
    .A2(\u_cpu.REG_FILE._02249_ ),
    .B1(\u_cpu.REG_FILE._02273_ ),
    .C1(\u_cpu.REG_FILE._02227_ ),
    .X(\u_cpu.ALU.SrcA[21] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06962_  (.A(\u_cpu.REG_FILE.rf[15][22] ),
    .B_N(\u_cpu.REG_FILE._01889_ ),
    .X(\u_cpu.REG_FILE._02274_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06963_  (.A1(\u_cpu.REG_FILE._01531_ ),
    .A2(\u_cpu.REG_FILE.rf[14][22] ),
    .B1(\u_cpu.REG_FILE._01288_ ),
    .C1(\u_cpu.REG_FILE._02274_ ),
    .Y(\u_cpu.REG_FILE._02275_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06964_  (.A1(\u_cpu.REG_FILE._01584_ ),
    .A2(\u_cpu.REG_FILE.rf[12][22] ),
    .B1_N(\u_cpu.REG_FILE._01838_ ),
    .X(\u_cpu.REG_FILE._02276_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06965_  (.A1(\u_cpu.REG_FILE._01787_ ),
    .A2(\u_cpu.REG_FILE.rf[13][22] ),
    .B1(\u_cpu.REG_FILE._02276_ ),
    .Y(\u_cpu.REG_FILE._02277_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06966_  (.A(\u_cpu.REG_FILE._02275_ ),
    .B(\u_cpu.REG_FILE._02277_ ),
    .C(\u_cpu.REG_FILE._01690_ ),
    .Y(\u_cpu.REG_FILE._02278_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06967_  (.A_N(\u_cpu.REG_FILE.rf[9][22] ),
    .B(\u_cpu.REG_FILE._01895_ ),
    .X(\u_cpu.REG_FILE._02279_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06968_  (.A1(\u_cpu.REG_FILE._01475_ ),
    .A2(\u_cpu.REG_FILE.rf[8][22] ),
    .B1_N(\u_cpu.REG_FILE._01843_ ),
    .Y(\u_cpu.REG_FILE._02280_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06969_  (.A(\u_cpu.REG_FILE.rf[11][22] ),
    .B_N(\u_cpu.REG_FILE._01590_ ),
    .X(\u_cpu.REG_FILE._02281_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06970_  (.A1(\u_cpu.REG_FILE._01620_ ),
    .A2(\u_cpu.REG_FILE.rf[10][22] ),
    .B1(\u_cpu.REG_FILE._01339_ ),
    .C1(\u_cpu.REG_FILE._02281_ ),
    .Y(\u_cpu.REG_FILE._02282_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06971_  (.A1(\u_cpu.REG_FILE._02279_ ),
    .A2(\u_cpu.REG_FILE._02280_ ),
    .B1(\u_cpu.REG_FILE._01384_ ),
    .C1(\u_cpu.REG_FILE._02282_ ),
    .Y(\u_cpu.REG_FILE._02283_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._06972_  (.A(\u_cpu.REG_FILE._02278_ ),
    .B(\u_cpu.REG_FILE._02283_ ),
    .C(\u_cpu.REG_FILE._01796_ ),
    .Y(\u_cpu.REG_FILE._02284_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._06973_  (.A(\u_cpu.REG_FILE.rf[5][22] ),
    .Y(\u_cpu.REG_FILE._02285_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06974_  (.A1(\u_cpu.REG_FILE._01133_ ),
    .A2(\u_cpu.REG_FILE.rf[4][22] ),
    .B1_N(\u_cpu.REG_FILE._01482_ ),
    .Y(\u_cpu.REG_FILE._02286_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._06975_  (.A1(\u_cpu.REG_FILE._02285_ ),
    .A2(\u_cpu.REG_FILE._01850_ ),
    .B1(\u_cpu.REG_FILE._02286_ ),
    .Y(\u_cpu.REG_FILE._02287_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06976_  (.A1(\u_cpu.REG_FILE._01774_ ),
    .A2(\u_cpu.REG_FILE.rf[6][22] ),
    .B1(\u_cpu.REG_FILE._01598_ ),
    .Y(\u_cpu.REG_FILE._02288_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06977_  (.A_N(\u_cpu.REG_FILE.rf[7][22] ),
    .B(\u_cpu.REG_FILE._01906_ ),
    .X(\u_cpu.REG_FILE._02289_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06978_  (.A1(\u_cpu.REG_FILE._02288_ ),
    .A2(\u_cpu.REG_FILE._02289_ ),
    .B1(\u_cpu.REG_FILE._01601_ ),
    .Y(\u_cpu.REG_FILE._02290_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06979_  (.A_N(\u_cpu.REG_FILE.rf[1][22] ),
    .B(\u_cpu.REG_FILE._01804_ ),
    .X(\u_cpu.REG_FILE._02291_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06980_  (.A1(\u_cpu.REG_FILE._02105_ ),
    .A2(\u_cpu.REG_FILE.rf[0][22] ),
    .B1_N(\u_cpu.REG_FILE._01705_ ),
    .Y(\u_cpu.REG_FILE._02292_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._06981_  (.A(\u_cpu.REG_FILE.rf[3][22] ),
    .B_N(\u_cpu.REG_FILE._02057_ ),
    .X(\u_cpu.REG_FILE._02293_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06982_  (.A1(\u_cpu.REG_FILE._01707_ ),
    .A2(\u_cpu.REG_FILE.rf[2][22] ),
    .B1(\u_cpu.REG_FILE._02056_ ),
    .C1(\u_cpu.REG_FILE._02293_ ),
    .Y(\u_cpu.REG_FILE._02294_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06983_  (.A1(\u_cpu.REG_FILE._02291_ ),
    .A2(\u_cpu.REG_FILE._02292_ ),
    .B1(\u_cpu.REG_FILE._01858_ ),
    .C1(\u_cpu.REG_FILE._02294_ ),
    .Y(\u_cpu.REG_FILE._02295_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06984_  (.A1(\u_cpu.REG_FILE._02287_ ),
    .A2(\u_cpu.REG_FILE._02290_ ),
    .B1(\u_cpu.REG_FILE._01603_ ),
    .C1(\u_cpu.REG_FILE._02295_ ),
    .Y(\u_cpu.REG_FILE._02296_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._06985_  (.A(\u_cpu.REG_FILE._02284_ ),
    .B(\u_cpu.REG_FILE._02296_ ),
    .Y(\u_cpu.REG_FILE._02297_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06986_  (.A1(\u_cpu.REG_FILE._01379_ ),
    .A2(\u_cpu.REG_FILE.rf[24][22] ),
    .B1_N(\u_cpu.REG_FILE._01611_ ),
    .Y(\u_cpu.REG_FILE._02298_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._06987_  (.A_N(\u_cpu.REG_FILE.rf[25][22] ),
    .B(\u_cpu.REG_FILE._01382_ ),
    .X(\u_cpu.REG_FILE._02299_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06988_  (.A1(\u_cpu.REG_FILE._02298_ ),
    .A2(\u_cpu.REG_FILE._02299_ ),
    .B1(\u_cpu.REG_FILE._01814_ ),
    .Y(\u_cpu.REG_FILE._02300_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._06989_  (.A(\u_cpu.REG_FILE._01340_ ),
    .B(\u_cpu.REG_FILE.rf[26][22] ),
    .X(\u_cpu.REG_FILE._02301_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._06990_  (.A1(\u_cpu.REG_FILE._01386_ ),
    .A2(\u_cpu.REG_FILE.rf[27][22] ),
    .B1(\u_cpu.REG_FILE._01387_ ),
    .C1(\u_cpu.REG_FILE._02301_ ),
    .X(\u_cpu.REG_FILE._02302_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06991_  (.A(\u_cpu.REG_FILE._01097_ ),
    .B(\u_cpu.REG_FILE.rf[30][22] ),
    .Y(\u_cpu.REG_FILE._02303_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06992_  (.A1(\u_cpu.REG_FILE.rf[31][22] ),
    .A2(\u_cpu.REG_FILE._01327_ ),
    .B1(\u_cpu.REG_FILE._01618_ ),
    .Y(\u_cpu.REG_FILE._02304_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._06993_  (.A(\u_cpu.REG_FILE._01325_ ),
    .B(\u_cpu.REG_FILE.rf[28][22] ),
    .Y(\u_cpu.REG_FILE._02305_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._06994_  (.A1(\u_cpu.REG_FILE.rf[29][22] ),
    .A2(\u_cpu.REG_FILE._01265_ ),
    .B1_N(\u_cpu.REG_FILE._01521_ ),
    .Y(\u_cpu.REG_FILE._02306_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._06995_  (.A1(\u_cpu.REG_FILE._02303_ ),
    .A2(\u_cpu.REG_FILE._02304_ ),
    .B1(\u_cpu.REG_FILE._02305_ ),
    .B2(\u_cpu.REG_FILE._02306_ ),
    .C1(\u_cpu.REG_FILE._01333_ ),
    .Y(\u_cpu.REG_FILE._02307_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._06996_  (.A1(\u_cpu.REG_FILE._02300_ ),
    .A2(\u_cpu.REG_FILE._02302_ ),
    .B1(\u_cpu.REG_FILE._01869_ ),
    .C1(\u_cpu.REG_FILE._02307_ ),
    .Y(\u_cpu.REG_FILE._02308_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.REG_FILE._06997_  (.A1(\u_cpu.REG_FILE._01528_ ),
    .A2(\u_cpu.REG_FILE.rf[18][22] ),
    .B1(\u_cpu.REG_FILE._01032_ ),
    .X(\u_cpu.REG_FILE._02309_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._06998_  (.A1(\u_cpu.REG_FILE.rf[19][22] ),
    .A2(\u_cpu.REG_FILE._01124_ ),
    .B1(\u_cpu.REG_FILE._02309_ ),
    .Y(\u_cpu.REG_FILE._02310_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._06999_  (.A1(\u_cpu.REG_FILE._01536_ ),
    .A2(\u_cpu.REG_FILE.rf[16][22] ),
    .B1_N(\u_cpu.REG_FILE._01134_ ),
    .X(\u_cpu.REG_FILE._02311_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07000_  (.A1(\u_cpu.REG_FILE._01120_ ),
    .A2(\u_cpu.REG_FILE.rf[17][22] ),
    .B1(\u_cpu.REG_FILE._02311_ ),
    .Y(\u_cpu.REG_FILE._02312_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07001_  (.A(\u_cpu.REG_FILE._01307_ ),
    .B(\u_cpu.REG_FILE._02310_ ),
    .C(\u_cpu.REG_FILE._02312_ ),
    .Y(\u_cpu.REG_FILE._02313_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._07002_  (.A(\u_cpu.REG_FILE._01269_ ),
    .B(\u_cpu.REG_FILE.rf[22][22] ),
    .X(\u_cpu.REG_FILE._02314_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07003_  (.A1(\u_cpu.REG_FILE._01321_ ),
    .A2(\u_cpu.REG_FILE.rf[23][22] ),
    .B1(\u_cpu.REG_FILE._01063_ ),
    .C1(\u_cpu.REG_FILE._02314_ ),
    .Y(\u_cpu.REG_FILE._02315_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07004_  (.A1(\u_cpu.REG_FILE._01632_ ),
    .A2(\u_cpu.REG_FILE.rf[20][22] ),
    .B1_N(\u_cpu.REG_FILE._01214_ ),
    .X(\u_cpu.REG_FILE._02316_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07005_  (.A1(\u_cpu.REG_FILE._01120_ ),
    .A2(\u_cpu.REG_FILE.rf[21][22] ),
    .B1(\u_cpu.REG_FILE._02316_ ),
    .Y(\u_cpu.REG_FILE._02317_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07006_  (.A(\u_cpu.REG_FILE._02315_ ),
    .B(\u_cpu.REG_FILE._02317_ ),
    .C(\u_cpu.REG_FILE._01552_ ),
    .Y(\u_cpu.REG_FILE._02318_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07007_  (.A(\u_cpu.REG_FILE._01569_ ),
    .B(\u_cpu.REG_FILE._02313_ ),
    .C(\u_cpu.REG_FILE._02318_ ),
    .Y(\u_cpu.REG_FILE._02319_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07008_  (.A(\u_cpu.REG_FILE._02308_ ),
    .B(\u_cpu.REG_FILE._02319_ ),
    .C(\u_cpu.REG_FILE._01684_ ),
    .Y(\u_cpu.REG_FILE._02320_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07009_  (.A1(\u_cpu.REG_FILE._01888_ ),
    .A2(\u_cpu.REG_FILE._02297_ ),
    .B1(\u_cpu.REG_FILE._02320_ ),
    .C1(\u_cpu.REG_FILE._02227_ ),
    .X(\u_cpu.ALU.SrcA[22] ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07010_  (.A1(\u_cpu.REG_FILE._01404_ ),
    .A2(\u_cpu.REG_FILE.rf[16][23] ),
    .B1_N(\u_cpu.REG_FILE._01553_ ),
    .Y(\u_cpu.REG_FILE._02321_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07011_  (.A_N(\u_cpu.REG_FILE.rf[17][23] ),
    .B(\u_cpu.REG_FILE._01750_ ),
    .X(\u_cpu.REG_FILE._02322_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07012_  (.A1(\u_cpu.REG_FILE._01279_ ),
    .A2(\u_cpu.REG_FILE.rf[18][23] ),
    .B1(\u_cpu.REG_FILE._01280_ ),
    .Y(\u_cpu.REG_FILE._02323_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07013_  (.A_N(\u_cpu.REG_FILE.rf[19][23] ),
    .B(\u_cpu.REG_FILE._01523_ ),
    .X(\u_cpu.REG_FILE._02324_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.REG_FILE._07014_  (.A1(\u_cpu.REG_FILE._02321_ ),
    .A2(\u_cpu.REG_FILE._02322_ ),
    .B1(\u_cpu.REG_FILE._02323_ ),
    .B2(\u_cpu.REG_FILE._02324_ ),
    .Y(\u_cpu.REG_FILE._02325_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07015_  (.A(\u_cpu.REG_FILE._01118_ ),
    .B(\u_cpu.REG_FILE.rf[20][23] ),
    .Y(\u_cpu.REG_FILE._02326_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07016_  (.A1(\u_cpu.REG_FILE.rf[21][23] ),
    .A2(\u_cpu.REG_FILE._01535_ ),
    .B1_N(\u_cpu.REG_FILE._01305_ ),
    .Y(\u_cpu.REG_FILE._02327_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._07017_  (.A(\u_cpu.REG_FILE._01536_ ),
    .B(\u_cpu.REG_FILE.rf[22][23] ),
    .X(\u_cpu.REG_FILE._02328_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07018_  (.A1(\u_cpu.REG_FILE._01535_ ),
    .A2(\u_cpu.REG_FILE.rf[23][23] ),
    .B1(\u_cpu.REG_FILE._01527_ ),
    .C1(\u_cpu.REG_FILE._02328_ ),
    .Y(\u_cpu.REG_FILE._02329_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07019_  (.A1(\u_cpu.REG_FILE._02326_ ),
    .A2(\u_cpu.REG_FILE._02327_ ),
    .B1(\u_cpu.REG_FILE._01129_ ),
    .C1(\u_cpu.REG_FILE._02329_ ),
    .Y(\u_cpu.REG_FILE._02330_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07020_  (.A1(\u_cpu.REG_FILE._02325_ ),
    .A2(\u_cpu.REG_FILE._01277_ ),
    .B1(\u_cpu.REG_FILE._01541_ ),
    .C1(\u_cpu.REG_FILE._02330_ ),
    .X(\u_cpu.REG_FILE._02331_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07021_  (.A(\u_cpu.REG_FILE.rf[31][23] ),
    .B_N(\u_cpu.REG_FILE._01111_ ),
    .X(\u_cpu.REG_FILE._02332_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07022_  (.A1(\u_cpu.REG_FILE._01030_ ),
    .A2(\u_cpu.REG_FILE.rf[30][23] ),
    .B1(\u_cpu.REG_FILE._01033_ ),
    .C1(\u_cpu.REG_FILE._02332_ ),
    .Y(\u_cpu.REG_FILE._02333_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07023_  (.A1(\u_cpu.REG_FILE._01299_ ),
    .A2(\u_cpu.REG_FILE.rf[28][23] ),
    .B1_N(\u_cpu.REG_FILE._01106_ ),
    .X(\u_cpu.REG_FILE._02334_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07024_  (.A1(\u_cpu.REG_FILE._01298_ ),
    .A2(\u_cpu.REG_FILE.rf[29][23] ),
    .B1(\u_cpu.REG_FILE._02334_ ),
    .Y(\u_cpu.REG_FILE._02335_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07025_  (.A(\u_cpu.REG_FILE._02333_ ),
    .B(\u_cpu.REG_FILE._02335_ ),
    .C(\u_cpu.REG_FILE._01293_ ),
    .Y(\u_cpu.REG_FILE._02336_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07026_  (.A_N(\u_cpu.REG_FILE.rf[25][23] ),
    .B(\u_cpu.REG_FILE._01547_ ),
    .X(\u_cpu.REG_FILE._02337_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07027_  (.A1(\u_cpu.REG_FILE._01549_ ),
    .A2(\u_cpu.REG_FILE.rf[24][23] ),
    .B1_N(\u_cpu.REG_FILE._01550_ ),
    .Y(\u_cpu.REG_FILE._02338_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07028_  (.A(\u_cpu.REG_FILE.rf[27][23] ),
    .B_N(\u_cpu.REG_FILE._01310_ ),
    .X(\u_cpu.REG_FILE._02339_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07029_  (.A1(\u_cpu.REG_FILE._01061_ ),
    .A2(\u_cpu.REG_FILE.rf[26][23] ),
    .B1(\u_cpu.REG_FILE._01309_ ),
    .C1(\u_cpu.REG_FILE._02339_ ),
    .Y(\u_cpu.REG_FILE._02340_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07030_  (.A1(\u_cpu.REG_FILE._02337_ ),
    .A2(\u_cpu.REG_FILE._02338_ ),
    .B1(\u_cpu.REG_FILE._01059_ ),
    .C1(\u_cpu.REG_FILE._02340_ ),
    .Y(\u_cpu.REG_FILE._02341_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._07031_  (.A1(\u_cpu.REG_FILE._02336_ ),
    .A2(\u_cpu.REG_FILE._02341_ ),
    .A3(\u_cpu.REG_FILE._01314_ ),
    .B1(\u_cpu.REG_FILE._01315_ ),
    .X(\u_cpu.REG_FILE._02342_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07032_  (.A(\u_cpu.REG_FILE.rf[5][23] ),
    .Y(\u_cpu.REG_FILE._02343_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07033_  (.A1(\u_cpu.REG_FILE._01260_ ),
    .A2(\u_cpu.REG_FILE.rf[4][23] ),
    .B1_N(\u_cpu.REG_FILE._01611_ ),
    .Y(\u_cpu.REG_FILE._02344_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07034_  (.A1(\u_cpu.REG_FILE._02343_ ),
    .A2(\u_cpu.REG_FILE._01284_ ),
    .B1(\u_cpu.REG_FILE._02344_ ),
    .Y(\u_cpu.REG_FILE._02345_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07035_  (.A1(\u_cpu.REG_FILE._01317_ ),
    .A2(\u_cpu.REG_FILE.rf[6][23] ),
    .B1(\u_cpu.REG_FILE._01400_ ),
    .Y(\u_cpu.REG_FILE._02346_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07036_  (.A_N(\u_cpu.REG_FILE.rf[7][23] ),
    .B(\u_cpu.REG_FILE._01161_ ),
    .X(\u_cpu.REG_FILE._02347_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07037_  (.A1(\u_cpu.REG_FILE._02346_ ),
    .A2(\u_cpu.REG_FILE._02347_ ),
    .B1(\u_cpu.REG_FILE._02122_ ),
    .Y(\u_cpu.REG_FILE._02348_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07038_  (.A_N(\u_cpu.REG_FILE.rf[1][23] ),
    .B(\u_cpu.REG_FILE._01041_ ),
    .X(\u_cpu.REG_FILE._02349_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07039_  (.A1(\u_cpu.REG_FILE._01260_ ),
    .A2(\u_cpu.REG_FILE.rf[0][23] ),
    .B1_N(\u_cpu.REG_FILE._01380_ ),
    .Y(\u_cpu.REG_FILE._02350_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07040_  (.A(\u_cpu.REG_FILE.rf[3][23] ),
    .B_N(\u_cpu.REG_FILE._01052_ ),
    .X(\u_cpu.REG_FILE._02351_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07041_  (.A1(\u_cpu.REG_FILE._01184_ ),
    .A2(\u_cpu.REG_FILE.rf[2][23] ),
    .B1(\u_cpu.REG_FILE._01407_ ),
    .C1(\u_cpu.REG_FILE._02351_ ),
    .Y(\u_cpu.REG_FILE._02352_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07042_  (.A1(\u_cpu.REG_FILE._02349_ ),
    .A2(\u_cpu.REG_FILE._02350_ ),
    .B1(\u_cpu.REG_FILE._01264_ ),
    .C1(\u_cpu.REG_FILE._02352_ ),
    .Y(\u_cpu.REG_FILE._02353_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07043_  (.A1(\u_cpu.REG_FILE._02345_ ),
    .A2(\u_cpu.REG_FILE._02348_ ),
    .B1(\u_cpu.REG_FILE._02353_ ),
    .Y(\u_cpu.REG_FILE._02354_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07044_  (.A(\u_cpu.REG_FILE._01620_ ),
    .B(\u_cpu.REG_FILE.rf[14][23] ),
    .Y(\u_cpu.REG_FILE._02355_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07045_  (.A1(\u_cpu.REG_FILE.rf[15][23] ),
    .A2(\u_cpu.REG_FILE._01329_ ),
    .B1(\u_cpu.REG_FILE._01280_ ),
    .Y(\u_cpu.REG_FILE._02356_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07046_  (.A1(\u_cpu.REG_FILE._01345_ ),
    .A2(\u_cpu.REG_FILE.rf[12][23] ),
    .B1_N(\u_cpu.REG_FILE._01134_ ),
    .X(\u_cpu.REG_FILE._02357_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07047_  (.A1(\u_cpu.REG_FILE._01265_ ),
    .A2(\u_cpu.REG_FILE.rf[13][23] ),
    .B1(\u_cpu.REG_FILE._02357_ ),
    .Y(\u_cpu.REG_FILE._02358_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07048_  (.A1(\u_cpu.REG_FILE._02355_ ),
    .A2(\u_cpu.REG_FILE._02356_ ),
    .B1(\u_cpu.REG_FILE._02358_ ),
    .C1(\u_cpu.REG_FILE._01333_ ),
    .Y(\u_cpu.REG_FILE._02359_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07049_  (.A(\u_cpu.REG_FILE.rf[11][23] ),
    .B_N(\u_cpu.REG_FILE._01052_ ),
    .X(\u_cpu.REG_FILE._02360_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07050_  (.A1(\u_cpu.REG_FILE._02105_ ),
    .A2(\u_cpu.REG_FILE.rf[10][23] ),
    .B1(\u_cpu.REG_FILE._01407_ ),
    .C1(\u_cpu.REG_FILE._02360_ ),
    .Y(\u_cpu.REG_FILE._02361_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07051_  (.A1(\u_cpu.REG_FILE._01330_ ),
    .A2(\u_cpu.REG_FILE.rf[8][23] ),
    .B1_N(\u_cpu.REG_FILE._01082_ ),
    .X(\u_cpu.REG_FILE._02362_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07052_  (.A1(\u_cpu.REG_FILE._01329_ ),
    .A2(\u_cpu.REG_FILE.rf[9][23] ),
    .B1(\u_cpu.REG_FILE._02362_ ),
    .Y(\u_cpu.REG_FILE._02363_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07053_  (.A(\u_cpu.REG_FILE._01307_ ),
    .B(\u_cpu.REG_FILE._02361_ ),
    .C(\u_cpu.REG_FILE._02363_ ),
    .Y(\u_cpu.REG_FILE._02364_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07054_  (.A(\u_cpu.REG_FILE._02359_ ),
    .B(\u_cpu.REG_FILE._02364_ ),
    .C(\u_cpu.REG_FILE._01069_ ),
    .Y(\u_cpu.REG_FILE._02365_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07055_  (.A1(\u_cpu.REG_FILE._01070_ ),
    .A2(\u_cpu.REG_FILE._02354_ ),
    .B1(\u_cpu.REG_FILE._02365_ ),
    .C1(\u_cpu.REG_FILE._01315_ ),
    .Y(\u_cpu.REG_FILE._02366_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07056_  (.A1(\u_cpu.REG_FILE._02331_ ),
    .A2(\u_cpu.REG_FILE._02342_ ),
    .B1(\u_cpu.REG_FILE._02366_ ),
    .C1(\u_cpu.REG_FILE._02227_ ),
    .X(\u_cpu.ALU.SrcA[23] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07057_  (.A(\u_cpu.REG_FILE.rf[15][24] ),
    .B_N(\u_cpu.REG_FILE._01889_ ),
    .X(\u_cpu.REG_FILE._02367_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07058_  (.A1(\u_cpu.REG_FILE._01531_ ),
    .A2(\u_cpu.REG_FILE.rf[14][24] ),
    .B1(\u_cpu.REG_FILE._01288_ ),
    .C1(\u_cpu.REG_FILE._02367_ ),
    .Y(\u_cpu.REG_FILE._02368_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07059_  (.A1(\u_cpu.REG_FILE._01584_ ),
    .A2(\u_cpu.REG_FILE.rf[12][24] ),
    .B1_N(\u_cpu.REG_FILE._01838_ ),
    .X(\u_cpu.REG_FILE._02369_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07060_  (.A1(\u_cpu.REG_FILE._01787_ ),
    .A2(\u_cpu.REG_FILE.rf[13][24] ),
    .B1(\u_cpu.REG_FILE._02369_ ),
    .Y(\u_cpu.REG_FILE._02370_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07061_  (.A(\u_cpu.REG_FILE._02368_ ),
    .B(\u_cpu.REG_FILE._02370_ ),
    .C(\u_cpu.REG_FILE._01690_ ),
    .Y(\u_cpu.REG_FILE._02371_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07062_  (.A_N(\u_cpu.REG_FILE.rf[9][24] ),
    .B(\u_cpu.REG_FILE._01895_ ),
    .X(\u_cpu.REG_FILE._02372_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07063_  (.A1(\u_cpu.REG_FILE._02018_ ),
    .A2(\u_cpu.REG_FILE.rf[8][24] ),
    .B1_N(\u_cpu.REG_FILE._01843_ ),
    .Y(\u_cpu.REG_FILE._02373_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07064_  (.A(\u_cpu.REG_FILE.rf[11][24] ),
    .B_N(\u_cpu.REG_FILE._01590_ ),
    .X(\u_cpu.REG_FILE._02374_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07065_  (.A1(\u_cpu.REG_FILE._01620_ ),
    .A2(\u_cpu.REG_FILE.rf[10][24] ),
    .B1(\u_cpu.REG_FILE._01339_ ),
    .C1(\u_cpu.REG_FILE._02374_ ),
    .Y(\u_cpu.REG_FILE._02375_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07066_  (.A1(\u_cpu.REG_FILE._02372_ ),
    .A2(\u_cpu.REG_FILE._02373_ ),
    .B1(\u_cpu.REG_FILE._01384_ ),
    .C1(\u_cpu.REG_FILE._02375_ ),
    .Y(\u_cpu.REG_FILE._02376_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07067_  (.A(\u_cpu.REG_FILE._02371_ ),
    .B(\u_cpu.REG_FILE._02376_ ),
    .C(\u_cpu.REG_FILE._01796_ ),
    .Y(\u_cpu.REG_FILE._02377_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07068_  (.A(\u_cpu.REG_FILE.rf[5][24] ),
    .Y(\u_cpu.REG_FILE._02378_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07069_  (.A1(\u_cpu.REG_FILE._01133_ ),
    .A2(\u_cpu.REG_FILE.rf[4][24] ),
    .B1_N(\u_cpu.REG_FILE._01380_ ),
    .Y(\u_cpu.REG_FILE._02379_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07070_  (.A1(\u_cpu.REG_FILE._02378_ ),
    .A2(\u_cpu.REG_FILE._01850_ ),
    .B1(\u_cpu.REG_FILE._02379_ ),
    .Y(\u_cpu.REG_FILE._02380_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07071_  (.A1(\u_cpu.REG_FILE._01774_ ),
    .A2(\u_cpu.REG_FILE.rf[6][24] ),
    .B1(\u_cpu.REG_FILE._01598_ ),
    .Y(\u_cpu.REG_FILE._02381_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07072_  (.A_N(\u_cpu.REG_FILE.rf[7][24] ),
    .B(\u_cpu.REG_FILE._01906_ ),
    .X(\u_cpu.REG_FILE._02382_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07073_  (.A1(\u_cpu.REG_FILE._02381_ ),
    .A2(\u_cpu.REG_FILE._02382_ ),
    .B1(\u_cpu.REG_FILE._01601_ ),
    .Y(\u_cpu.REG_FILE._02383_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07074_  (.A_N(\u_cpu.REG_FILE.rf[1][24] ),
    .B(\u_cpu.REG_FILE._01804_ ),
    .X(\u_cpu.REG_FILE._02384_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07075_  (.A1(\u_cpu.REG_FILE._02105_ ),
    .A2(\u_cpu.REG_FILE.rf[0][24] ),
    .B1_N(\u_cpu.REG_FILE._01705_ ),
    .Y(\u_cpu.REG_FILE._02385_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07076_  (.A(\u_cpu.REG_FILE.rf[3][24] ),
    .B_N(\u_cpu.REG_FILE._02057_ ),
    .X(\u_cpu.REG_FILE._02386_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07077_  (.A1(\u_cpu.REG_FILE._01707_ ),
    .A2(\u_cpu.REG_FILE.rf[2][24] ),
    .B1(\u_cpu.REG_FILE._02056_ ),
    .C1(\u_cpu.REG_FILE._02386_ ),
    .Y(\u_cpu.REG_FILE._02387_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07078_  (.A1(\u_cpu.REG_FILE._02384_ ),
    .A2(\u_cpu.REG_FILE._02385_ ),
    .B1(\u_cpu.REG_FILE._01858_ ),
    .C1(\u_cpu.REG_FILE._02387_ ),
    .Y(\u_cpu.REG_FILE._02388_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07079_  (.A1(\u_cpu.REG_FILE._02380_ ),
    .A2(\u_cpu.REG_FILE._02383_ ),
    .B1(\u_cpu.REG_FILE._01603_ ),
    .C1(\u_cpu.REG_FILE._02388_ ),
    .Y(\u_cpu.REG_FILE._02389_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._07080_  (.A(\u_cpu.REG_FILE._02377_ ),
    .B(\u_cpu.REG_FILE._02389_ ),
    .Y(\u_cpu.REG_FILE._02390_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07081_  (.A1(\u_cpu.REG_FILE._01379_ ),
    .A2(\u_cpu.REG_FILE.rf[24][24] ),
    .B1_N(\u_cpu.REG_FILE._01611_ ),
    .Y(\u_cpu.REG_FILE._02391_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07082_  (.A_N(\u_cpu.REG_FILE.rf[25][24] ),
    .B(\u_cpu.REG_FILE._01750_ ),
    .X(\u_cpu.REG_FILE._02392_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07083_  (.A1(\u_cpu.REG_FILE._02391_ ),
    .A2(\u_cpu.REG_FILE._02392_ ),
    .B1(\u_cpu.REG_FILE._01814_ ),
    .Y(\u_cpu.REG_FILE._02393_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._07084_  (.A(\u_cpu.REG_FILE._01340_ ),
    .B(\u_cpu.REG_FILE.rf[26][24] ),
    .X(\u_cpu.REG_FILE._02394_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07085_  (.A1(\u_cpu.REG_FILE._01386_ ),
    .A2(\u_cpu.REG_FILE.rf[27][24] ),
    .B1(\u_cpu.REG_FILE._01121_ ),
    .C1(\u_cpu.REG_FILE._02394_ ),
    .X(\u_cpu.REG_FILE._02395_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07086_  (.A(\u_cpu.REG_FILE._02010_ ),
    .B(\u_cpu.REG_FILE.rf[30][24] ),
    .Y(\u_cpu.REG_FILE._02396_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07087_  (.A1(\u_cpu.REG_FILE.rf[31][24] ),
    .A2(\u_cpu.REG_FILE._01969_ ),
    .B1(\u_cpu.REG_FILE._01501_ ),
    .Y(\u_cpu.REG_FILE._02397_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07088_  (.A1(\u_cpu.REG_FILE._01503_ ),
    .A2(\u_cpu.REG_FILE.rf[28][24] ),
    .B1_N(\u_cpu.REG_FILE._01098_ ),
    .X(\u_cpu.REG_FILE._02398_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07089_  (.A1(\u_cpu.REG_FILE._01668_ ),
    .A2(\u_cpu.REG_FILE.rf[29][24] ),
    .B1(\u_cpu.REG_FILE._02398_ ),
    .Y(\u_cpu.REG_FILE._02399_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07090_  (.A1(\u_cpu.REG_FILE._02396_ ),
    .A2(\u_cpu.REG_FILE._02397_ ),
    .B1(\u_cpu.REG_FILE._02399_ ),
    .C1(\u_cpu.REG_FILE._02016_ ),
    .Y(\u_cpu.REG_FILE._02400_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07091_  (.A1(\u_cpu.REG_FILE._02393_ ),
    .A2(\u_cpu.REG_FILE._02395_ ),
    .B1(\u_cpu.REG_FILE._01869_ ),
    .C1(\u_cpu.REG_FILE._02400_ ),
    .Y(\u_cpu.REG_FILE._02401_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07092_  (.A(\u_cpu.REG_FILE.rf[19][24] ),
    .Y(\u_cpu.REG_FILE._02402_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07093_  (.A1(\u_cpu.REG_FILE._01523_ ),
    .A2(\u_cpu.REG_FILE.rf[18][24] ),
    .B1(\u_cpu.REG_FILE._01533_ ),
    .Y(\u_cpu.REG_FILE._02403_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07094_  (.A1(\u_cpu.REG_FILE._02402_ ),
    .A2(\u_cpu.REG_FILE._01399_ ),
    .B1(\u_cpu.REG_FILE._02403_ ),
    .Y(\u_cpu.REG_FILE._02404_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07095_  (.A(\u_cpu.REG_FILE.rf[17][24] ),
    .Y(\u_cpu.REG_FILE._02405_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07096_  (.A1(\u_cpu.REG_FILE._01404_ ),
    .A2(\u_cpu.REG_FILE.rf[16][24] ),
    .B1_N(\u_cpu.REG_FILE._01258_ ),
    .Y(\u_cpu.REG_FILE._02406_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07097_  (.A1(\u_cpu.REG_FILE._02405_ ),
    .A2(\u_cpu.REG_FILE._01399_ ),
    .B1(\u_cpu.REG_FILE._02406_ ),
    .Y(\u_cpu.REG_FILE._02407_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07098_  (.A(\u_cpu.REG_FILE.rf[23][24] ),
    .B_N(\u_cpu.REG_FILE._01408_ ),
    .X(\u_cpu.REG_FILE._02408_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07099_  (.A1(\u_cpu.REG_FILE._01077_ ),
    .A2(\u_cpu.REG_FILE.rf[22][24] ),
    .B1(\u_cpu.REG_FILE._01407_ ),
    .C1(\u_cpu.REG_FILE._02408_ ),
    .Y(\u_cpu.REG_FILE._02409_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07100_  (.A1(\u_cpu.REG_FILE._01324_ ),
    .A2(\u_cpu.REG_FILE.rf[20][24] ),
    .B1_N(\u_cpu.REG_FILE._01304_ ),
    .X(\u_cpu.REG_FILE._02410_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07101_  (.A1(\u_cpu.REG_FILE._01038_ ),
    .A2(\u_cpu.REG_FILE.rf[21][24] ),
    .B1(\u_cpu.REG_FILE._02410_ ),
    .Y(\u_cpu.REG_FILE._02411_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07102_  (.A(\u_cpu.REG_FILE._02409_ ),
    .B(\u_cpu.REG_FILE._02411_ ),
    .C(\u_cpu.REG_FILE._01115_ ),
    .Y(\u_cpu.REG_FILE._02412_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._07103_  (.A1(\u_cpu.REG_FILE._01047_ ),
    .A2(\u_cpu.REG_FILE._02404_ ),
    .A3(\u_cpu.REG_FILE._02407_ ),
    .B1(\u_cpu.REG_FILE._02412_ ),
    .C1(\u_cpu.REG_FILE._01414_ ),
    .Y(\u_cpu.REG_FILE._02413_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07104_  (.A(\u_cpu.REG_FILE._02401_ ),
    .B(\u_cpu.REG_FILE._02413_ ),
    .C(\u_cpu.REG_FILE._01684_ ),
    .Y(\u_cpu.REG_FILE._02414_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07105_  (.A1(\u_cpu.REG_FILE._01888_ ),
    .A2(\u_cpu.REG_FILE._02390_ ),
    .B1(\u_cpu.REG_FILE._02414_ ),
    .C1(\u_cpu.REG_FILE._02227_ ),
    .X(\u_cpu.ALU.SrcA[24] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07106_  (.A(\u_cpu.REG_FILE.rf[15][25] ),
    .B_N(\u_cpu.REG_FILE._01889_ ),
    .X(\u_cpu.REG_FILE._02415_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07107_  (.A1(\u_cpu.REG_FILE._01531_ ),
    .A2(\u_cpu.REG_FILE.rf[14][25] ),
    .B1(\u_cpu.REG_FILE._01288_ ),
    .C1(\u_cpu.REG_FILE._02415_ ),
    .Y(\u_cpu.REG_FILE._02416_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07108_  (.A1(\u_cpu.REG_FILE._01299_ ),
    .A2(\u_cpu.REG_FILE.rf[12][25] ),
    .B1_N(\u_cpu.REG_FILE._01838_ ),
    .X(\u_cpu.REG_FILE._02417_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07109_  (.A1(\u_cpu.REG_FILE._01787_ ),
    .A2(\u_cpu.REG_FILE.rf[13][25] ),
    .B1(\u_cpu.REG_FILE._02417_ ),
    .Y(\u_cpu.REG_FILE._02418_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07110_  (.A(\u_cpu.REG_FILE._02416_ ),
    .B(\u_cpu.REG_FILE._02418_ ),
    .C(\u_cpu.REG_FILE._01690_ ),
    .Y(\u_cpu.REG_FILE._02419_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07111_  (.A_N(\u_cpu.REG_FILE.rf[9][25] ),
    .B(\u_cpu.REG_FILE._01895_ ),
    .X(\u_cpu.REG_FILE._02420_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07112_  (.A1(\u_cpu.REG_FILE._02018_ ),
    .A2(\u_cpu.REG_FILE.rf[8][25] ),
    .B1_N(\u_cpu.REG_FILE._01843_ ),
    .Y(\u_cpu.REG_FILE._02421_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07113_  (.A(\u_cpu.REG_FILE.rf[11][25] ),
    .B_N(\u_cpu.REG_FILE._01345_ ),
    .X(\u_cpu.REG_FILE._02422_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07114_  (.A1(\u_cpu.REG_FILE._01620_ ),
    .A2(\u_cpu.REG_FILE.rf[10][25] ),
    .B1(\u_cpu.REG_FILE._01339_ ),
    .C1(\u_cpu.REG_FILE._02422_ ),
    .Y(\u_cpu.REG_FILE._02423_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07115_  (.A1(\u_cpu.REG_FILE._02420_ ),
    .A2(\u_cpu.REG_FILE._02421_ ),
    .B1(\u_cpu.REG_FILE._01384_ ),
    .C1(\u_cpu.REG_FILE._02423_ ),
    .Y(\u_cpu.REG_FILE._02424_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07116_  (.A(\u_cpu.REG_FILE._02419_ ),
    .B(\u_cpu.REG_FILE._02424_ ),
    .C(\u_cpu.REG_FILE._01796_ ),
    .Y(\u_cpu.REG_FILE._02425_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07117_  (.A(\u_cpu.REG_FILE.rf[5][25] ),
    .Y(\u_cpu.REG_FILE._02426_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07118_  (.A1(\u_cpu.REG_FILE._01133_ ),
    .A2(\u_cpu.REG_FILE.rf[4][25] ),
    .B1_N(\u_cpu.REG_FILE._01380_ ),
    .Y(\u_cpu.REG_FILE._02427_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07119_  (.A1(\u_cpu.REG_FILE._02426_ ),
    .A2(\u_cpu.REG_FILE._01850_ ),
    .B1(\u_cpu.REG_FILE._02427_ ),
    .Y(\u_cpu.REG_FILE._02428_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07120_  (.A1(\u_cpu.REG_FILE._01774_ ),
    .A2(\u_cpu.REG_FILE.rf[6][25] ),
    .B1(\u_cpu.REG_FILE._01400_ ),
    .Y(\u_cpu.REG_FILE._02429_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07121_  (.A_N(\u_cpu.REG_FILE.rf[7][25] ),
    .B(\u_cpu.REG_FILE._01906_ ),
    .X(\u_cpu.REG_FILE._02430_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07122_  (.A1(\u_cpu.REG_FILE._02429_ ),
    .A2(\u_cpu.REG_FILE._02430_ ),
    .B1(\u_cpu.REG_FILE._02122_ ),
    .Y(\u_cpu.REG_FILE._02431_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07123_  (.A_N(\u_cpu.REG_FILE.rf[1][25] ),
    .B(\u_cpu.REG_FILE._01804_ ),
    .X(\u_cpu.REG_FILE._02432_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07124_  (.A1(\u_cpu.REG_FILE._02105_ ),
    .A2(\u_cpu.REG_FILE.rf[0][25] ),
    .B1_N(\u_cpu.REG_FILE._01705_ ),
    .Y(\u_cpu.REG_FILE._02433_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07125_  (.A(\u_cpu.REG_FILE.rf[3][25] ),
    .B_N(\u_cpu.REG_FILE._02057_ ),
    .X(\u_cpu.REG_FILE._02434_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07126_  (.A1(\u_cpu.REG_FILE._01707_ ),
    .A2(\u_cpu.REG_FILE.rf[2][25] ),
    .B1(\u_cpu.REG_FILE._02056_ ),
    .C1(\u_cpu.REG_FILE._02434_ ),
    .Y(\u_cpu.REG_FILE._02435_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07127_  (.A1(\u_cpu.REG_FILE._02432_ ),
    .A2(\u_cpu.REG_FILE._02433_ ),
    .B1(\u_cpu.REG_FILE._01858_ ),
    .C1(\u_cpu.REG_FILE._02435_ ),
    .Y(\u_cpu.REG_FILE._02436_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07128_  (.A1(\u_cpu.REG_FILE._02428_ ),
    .A2(\u_cpu.REG_FILE._02431_ ),
    .B1(\u_cpu.REG_FILE._01414_ ),
    .C1(\u_cpu.REG_FILE._02436_ ),
    .Y(\u_cpu.REG_FILE._02437_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._07129_  (.A(\u_cpu.REG_FILE._02425_ ),
    .B(\u_cpu.REG_FILE._02437_ ),
    .Y(\u_cpu.REG_FILE._02438_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07130_  (.A1(\u_cpu.REG_FILE._01081_ ),
    .A2(\u_cpu.REG_FILE.rf[24][25] ),
    .B1_N(\u_cpu.REG_FILE._01611_ ),
    .Y(\u_cpu.REG_FILE._02439_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07131_  (.A_N(\u_cpu.REG_FILE.rf[25][25] ),
    .B(\u_cpu.REG_FILE._01750_ ),
    .X(\u_cpu.REG_FILE._02440_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07132_  (.A1(\u_cpu.REG_FILE._02439_ ),
    .A2(\u_cpu.REG_FILE._02440_ ),
    .B1(\u_cpu.REG_FILE._01814_ ),
    .Y(\u_cpu.REG_FILE._02441_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._07133_  (.A(\u_cpu.REG_FILE._01340_ ),
    .B(\u_cpu.REG_FILE.rf[26][25] ),
    .X(\u_cpu.REG_FILE._02442_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07134_  (.A1(\u_cpu.REG_FILE._01386_ ),
    .A2(\u_cpu.REG_FILE.rf[27][25] ),
    .B1(\u_cpu.REG_FILE._01121_ ),
    .C1(\u_cpu.REG_FILE._02442_ ),
    .X(\u_cpu.REG_FILE._02443_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07135_  (.A(\u_cpu.REG_FILE._01097_ ),
    .B(\u_cpu.REG_FILE.rf[30][25] ),
    .Y(\u_cpu.REG_FILE._02444_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07136_  (.A1(\u_cpu.REG_FILE.rf[31][25] ),
    .A2(\u_cpu.REG_FILE._01327_ ),
    .B1(\u_cpu.REG_FILE._01618_ ),
    .Y(\u_cpu.REG_FILE._02445_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07137_  (.A(\u_cpu.REG_FILE._01325_ ),
    .B(\u_cpu.REG_FILE.rf[28][25] ),
    .Y(\u_cpu.REG_FILE._02446_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07138_  (.A1(\u_cpu.REG_FILE.rf[29][25] ),
    .A2(\u_cpu.REG_FILE._01265_ ),
    .B1_N(\u_cpu.REG_FILE._01521_ ),
    .Y(\u_cpu.REG_FILE._02447_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._07139_  (.A1(\u_cpu.REG_FILE._02444_ ),
    .A2(\u_cpu.REG_FILE._02445_ ),
    .B1(\u_cpu.REG_FILE._02446_ ),
    .B2(\u_cpu.REG_FILE._02447_ ),
    .C1(\u_cpu.REG_FILE._01333_ ),
    .Y(\u_cpu.REG_FILE._02448_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07140_  (.A1(\u_cpu.REG_FILE._02441_ ),
    .A2(\u_cpu.REG_FILE._02443_ ),
    .B1(\u_cpu.REG_FILE._01869_ ),
    .C1(\u_cpu.REG_FILE._02448_ ),
    .Y(\u_cpu.REG_FILE._02449_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07141_  (.A1(\u_cpu.REG_FILE._01206_ ),
    .A2(\u_cpu.REG_FILE.rf[18][25] ),
    .B1(\u_cpu.REG_FILE._01135_ ),
    .Y(\u_cpu.REG_FILE._02450_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07142_  (.A(\u_cpu.REG_FILE.rf[19][25] ),
    .B(\u_cpu.REG_FILE._01509_ ),
    .Y(\u_cpu.REG_FILE._02451_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07143_  (.A1(\u_cpu.REG_FILE._01141_ ),
    .A2(\u_cpu.REG_FILE.rf[16][25] ),
    .B1_N(\u_cpu.REG_FILE._01153_ ),
    .X(\u_cpu.REG_FILE._02452_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07144_  (.A1(\u_cpu.REG_FILE._01726_ ),
    .A2(\u_cpu.REG_FILE.rf[17][25] ),
    .B1(\u_cpu.REG_FILE._02452_ ),
    .Y(\u_cpu.REG_FILE._02453_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07145_  (.A1(\u_cpu.REG_FILE._02450_ ),
    .A2(\u_cpu.REG_FILE._02451_ ),
    .B1(\u_cpu.REG_FILE._01264_ ),
    .C1(\u_cpu.REG_FILE._02453_ ),
    .Y(\u_cpu.REG_FILE._02454_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._07146_  (.A(\u_cpu.REG_FILE._01269_ ),
    .B(\u_cpu.REG_FILE.rf[22][25] ),
    .X(\u_cpu.REG_FILE._02455_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07147_  (.A1(\u_cpu.REG_FILE._01321_ ),
    .A2(\u_cpu.REG_FILE.rf[23][25] ),
    .B1(\u_cpu.REG_FILE._01063_ ),
    .C1(\u_cpu.REG_FILE._02455_ ),
    .Y(\u_cpu.REG_FILE._02456_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07148_  (.A1(\u_cpu.REG_FILE._01632_ ),
    .A2(\u_cpu.REG_FILE.rf[20][25] ),
    .B1_N(\u_cpu.REG_FILE._01134_ ),
    .X(\u_cpu.REG_FILE._02457_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07149_  (.A1(\u_cpu.REG_FILE._01120_ ),
    .A2(\u_cpu.REG_FILE.rf[21][25] ),
    .B1(\u_cpu.REG_FILE._02457_ ),
    .Y(\u_cpu.REG_FILE._02458_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07150_  (.A(\u_cpu.REG_FILE._02456_ ),
    .B(\u_cpu.REG_FILE._02458_ ),
    .C(\u_cpu.REG_FILE._01552_ ),
    .Y(\u_cpu.REG_FILE._02459_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07151_  (.A(\u_cpu.REG_FILE._01569_ ),
    .B(\u_cpu.REG_FILE._02454_ ),
    .C(\u_cpu.REG_FILE._02459_ ),
    .Y(\u_cpu.REG_FILE._02460_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07152_  (.A(\u_cpu.REG_FILE._02449_ ),
    .B(\u_cpu.REG_FILE._02460_ ),
    .C(\u_cpu.REG_FILE._01684_ ),
    .Y(\u_cpu.REG_FILE._02461_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07153_  (.A1(\u_cpu.REG_FILE._01888_ ),
    .A2(\u_cpu.REG_FILE._02438_ ),
    .B1(\u_cpu.REG_FILE._02461_ ),
    .C1(\u_cpu.REG_FILE._02227_ ),
    .X(\u_cpu.ALU.SrcA[25] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07154_  (.A(\u_cpu.REG_FILE.rf[15][26] ),
    .B_N(\u_cpu.REG_FILE._01889_ ),
    .X(\u_cpu.REG_FILE._02462_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07155_  (.A1(\u_cpu.REG_FILE._01531_ ),
    .A2(\u_cpu.REG_FILE.rf[14][26] ),
    .B1(\u_cpu.REG_FILE._01288_ ),
    .C1(\u_cpu.REG_FILE._02462_ ),
    .Y(\u_cpu.REG_FILE._02463_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07156_  (.A1(\u_cpu.REG_FILE._01299_ ),
    .A2(\u_cpu.REG_FILE.rf[12][26] ),
    .B1_N(\u_cpu.REG_FILE._01838_ ),
    .X(\u_cpu.REG_FILE._02464_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07157_  (.A1(\u_cpu.REG_FILE._01787_ ),
    .A2(\u_cpu.REG_FILE.rf[13][26] ),
    .B1(\u_cpu.REG_FILE._02464_ ),
    .Y(\u_cpu.REG_FILE._02465_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07158_  (.A(\u_cpu.REG_FILE._02463_ ),
    .B(\u_cpu.REG_FILE._02465_ ),
    .C(\u_cpu.REG_FILE._01293_ ),
    .Y(\u_cpu.REG_FILE._02466_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07159_  (.A_N(\u_cpu.REG_FILE.rf[9][26] ),
    .B(\u_cpu.REG_FILE._01895_ ),
    .X(\u_cpu.REG_FILE._02467_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07160_  (.A1(\u_cpu.REG_FILE._02018_ ),
    .A2(\u_cpu.REG_FILE.rf[8][26] ),
    .B1_N(\u_cpu.REG_FILE._01843_ ),
    .Y(\u_cpu.REG_FILE._02468_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07161_  (.A(\u_cpu.REG_FILE.rf[11][26] ),
    .B_N(\u_cpu.REG_FILE._01345_ ),
    .X(\u_cpu.REG_FILE._02469_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07162_  (.A1(\u_cpu.REG_FILE._01620_ ),
    .A2(\u_cpu.REG_FILE.rf[10][26] ),
    .B1(\u_cpu.REG_FILE._01339_ ),
    .C1(\u_cpu.REG_FILE._02469_ ),
    .Y(\u_cpu.REG_FILE._02470_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07163_  (.A1(\u_cpu.REG_FILE._02467_ ),
    .A2(\u_cpu.REG_FILE._02468_ ),
    .B1(\u_cpu.REG_FILE._01384_ ),
    .C1(\u_cpu.REG_FILE._02470_ ),
    .Y(\u_cpu.REG_FILE._02471_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07164_  (.A(\u_cpu.REG_FILE._02466_ ),
    .B(\u_cpu.REG_FILE._02471_ ),
    .C(\u_cpu.REG_FILE._01796_ ),
    .Y(\u_cpu.REG_FILE._02472_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07165_  (.A(\u_cpu.REG_FILE.rf[5][26] ),
    .Y(\u_cpu.REG_FILE._02473_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07166_  (.A1(\u_cpu.REG_FILE._01133_ ),
    .A2(\u_cpu.REG_FILE.rf[4][26] ),
    .B1_N(\u_cpu.REG_FILE._01380_ ),
    .Y(\u_cpu.REG_FILE._02474_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07167_  (.A1(\u_cpu.REG_FILE._02473_ ),
    .A2(\u_cpu.REG_FILE._01850_ ),
    .B1(\u_cpu.REG_FILE._02474_ ),
    .Y(\u_cpu.REG_FILE._02475_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07168_  (.A1(\u_cpu.REG_FILE._01774_ ),
    .A2(\u_cpu.REG_FILE.rf[6][26] ),
    .B1(\u_cpu.REG_FILE._01400_ ),
    .Y(\u_cpu.REG_FILE._02476_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07169_  (.A_N(\u_cpu.REG_FILE.rf[7][26] ),
    .B(\u_cpu.REG_FILE._01906_ ),
    .X(\u_cpu.REG_FILE._02477_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07170_  (.A1(\u_cpu.REG_FILE._02476_ ),
    .A2(\u_cpu.REG_FILE._02477_ ),
    .B1(\u_cpu.REG_FILE._02122_ ),
    .Y(\u_cpu.REG_FILE._02478_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07171_  (.A_N(\u_cpu.REG_FILE.rf[1][26] ),
    .B(\u_cpu.REG_FILE._01804_ ),
    .X(\u_cpu.REG_FILE._02479_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07172_  (.A1(\u_cpu.REG_FILE._02105_ ),
    .A2(\u_cpu.REG_FILE.rf[0][26] ),
    .B1_N(\u_cpu.REG_FILE._01078_ ),
    .Y(\u_cpu.REG_FILE._02480_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07173_  (.A(\u_cpu.REG_FILE.rf[3][26] ),
    .B_N(\u_cpu.REG_FILE._02057_ ),
    .X(\u_cpu.REG_FILE._02481_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07174_  (.A1(\u_cpu.REG_FILE._01053_ ),
    .A2(\u_cpu.REG_FILE.rf[2][26] ),
    .B1(\u_cpu.REG_FILE._02056_ ),
    .C1(\u_cpu.REG_FILE._02481_ ),
    .Y(\u_cpu.REG_FILE._02482_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07175_  (.A1(\u_cpu.REG_FILE._02479_ ),
    .A2(\u_cpu.REG_FILE._02480_ ),
    .B1(\u_cpu.REG_FILE._01858_ ),
    .C1(\u_cpu.REG_FILE._02482_ ),
    .Y(\u_cpu.REG_FILE._02483_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07176_  (.A1(\u_cpu.REG_FILE._02475_ ),
    .A2(\u_cpu.REG_FILE._02478_ ),
    .B1(\u_cpu.REG_FILE._01414_ ),
    .C1(\u_cpu.REG_FILE._02483_ ),
    .Y(\u_cpu.REG_FILE._02484_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._07177_  (.A(\u_cpu.REG_FILE._02472_ ),
    .B(\u_cpu.REG_FILE._02484_ ),
    .Y(\u_cpu.REG_FILE._02485_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07178_  (.A(\u_cpu.REG_FILE.rf[19][26] ),
    .Y(\u_cpu.REG_FILE._02486_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07179_  (.A1(\u_cpu.REG_FILE._01081_ ),
    .A2(\u_cpu.REG_FILE.rf[18][26] ),
    .B1(\u_cpu.REG_FILE._01083_ ),
    .Y(\u_cpu.REG_FILE._02487_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07180_  (.A1(\u_cpu.REG_FILE._02486_ ),
    .A2(\u_cpu.REG_FILE._01284_ ),
    .B1(\u_cpu.REG_FILE._02487_ ),
    .Y(\u_cpu.REG_FILE._02488_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07181_  (.A(\u_cpu.REG_FILE.rf[17][26] ),
    .Y(\u_cpu.REG_FILE._02489_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07182_  (.A(\u_cpu.REG_FILE._01184_ ),
    .B(\u_cpu.REG_FILE.rf[16][26] ),
    .Y(\u_cpu.REG_FILE._02490_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._07183_  (.A1(\u_cpu.REG_FILE._02489_ ),
    .A2(\u_cpu.REG_FILE._01030_ ),
    .B1(\u_cpu.REG_FILE._01259_ ),
    .C1(\u_cpu.REG_FILE._02490_ ),
    .Y(\u_cpu.REG_FILE._02491_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._07184_  (.A(\u_cpu.REG_FILE._01408_ ),
    .B(\u_cpu.REG_FILE.rf[22][26] ),
    .X(\u_cpu.REG_FILE._02492_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07185_  (.A1(\u_cpu.REG_FILE._01327_ ),
    .A2(\u_cpu.REG_FILE.rf[23][26] ),
    .B1(\u_cpu.REG_FILE._01618_ ),
    .C1(\u_cpu.REG_FILE._02492_ ),
    .Y(\u_cpu.REG_FILE._02493_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07186_  (.A1(\u_cpu.REG_FILE._01330_ ),
    .A2(\u_cpu.REG_FILE.rf[20][26] ),
    .B1_N(\u_cpu.REG_FILE._01082_ ),
    .X(\u_cpu.REG_FILE._02494_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07187_  (.A1(\u_cpu.REG_FILE._01329_ ),
    .A2(\u_cpu.REG_FILE.rf[21][26] ),
    .B1(\u_cpu.REG_FILE._02494_ ),
    .Y(\u_cpu.REG_FILE._02495_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07188_  (.A(\u_cpu.REG_FILE._02493_ ),
    .B(\u_cpu.REG_FILE._02495_ ),
    .C(\u_cpu.REG_FILE._02122_ ),
    .Y(\u_cpu.REG_FILE._02496_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._07189_  (.A1(\u_cpu.REG_FILE._01277_ ),
    .A2(\u_cpu.REG_FILE._02488_ ),
    .A3(\u_cpu.REG_FILE._02491_ ),
    .B1(\u_cpu.REG_FILE._02496_ ),
    .C1(\u_cpu.REG_FILE._01090_ ),
    .Y(\u_cpu.REG_FILE._02497_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07190_  (.A(\u_cpu.REG_FILE.rf[27][26] ),
    .B_N(\u_cpu.REG_FILE._01330_ ),
    .X(\u_cpu.REG_FILE._02498_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07191_  (.A1(\u_cpu.REG_FILE._01093_ ),
    .A2(\u_cpu.REG_FILE.rf[26][26] ),
    .B1(\u_cpu.REG_FILE._01099_ ),
    .C1(\u_cpu.REG_FILE._02498_ ),
    .X(\u_cpu.REG_FILE._02499_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07192_  (.A1(\u_cpu.REG_FILE._01404_ ),
    .A2(\u_cpu.REG_FILE.rf[24][26] ),
    .B1_N(\u_cpu.REG_FILE._01553_ ),
    .Y(\u_cpu.REG_FILE._02500_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07193_  (.A_N(\u_cpu.REG_FILE.rf[25][26] ),
    .B(\u_cpu.REG_FILE._01750_ ),
    .X(\u_cpu.REG_FILE._02501_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07194_  (.A1(\u_cpu.REG_FILE._02500_ ),
    .A2(\u_cpu.REG_FILE._02501_ ),
    .B1(\u_cpu.REG_FILE._01096_ ),
    .Y(\u_cpu.REG_FILE._02502_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07195_  (.A(\u_cpu.REG_FILE._01325_ ),
    .B(\u_cpu.REG_FILE.rf[28][26] ),
    .Y(\u_cpu.REG_FILE._02503_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07196_  (.A1(\u_cpu.REG_FILE.rf[29][26] ),
    .A2(\u_cpu.REG_FILE._01329_ ),
    .B1_N(\u_cpu.REG_FILE._01094_ ),
    .Y(\u_cpu.REG_FILE._02504_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._07197_  (.A(\u_cpu.REG_FILE._01052_ ),
    .B(\u_cpu.REG_FILE.rf[30][26] ),
    .X(\u_cpu.REG_FILE._02505_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07198_  (.A1(\u_cpu.REG_FILE._01327_ ),
    .A2(\u_cpu.REG_FILE.rf[31][26] ),
    .B1(\u_cpu.REG_FILE._01099_ ),
    .C1(\u_cpu.REG_FILE._02505_ ),
    .Y(\u_cpu.REG_FILE._02506_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07199_  (.A1(\u_cpu.REG_FILE._02503_ ),
    .A2(\u_cpu.REG_FILE._02504_ ),
    .B1(\u_cpu.REG_FILE._02122_ ),
    .C1(\u_cpu.REG_FILE._02506_ ),
    .Y(\u_cpu.REG_FILE._02507_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07200_  (.A1(\u_cpu.REG_FILE._02499_ ),
    .A2(\u_cpu.REG_FILE._02502_ ),
    .B1(\u_cpu.REG_FILE._01069_ ),
    .C1(\u_cpu.REG_FILE._02507_ ),
    .Y(\u_cpu.REG_FILE._02508_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07201_  (.A(\u_cpu.REG_FILE._02497_ ),
    .B(\u_cpu.REG_FILE._01025_ ),
    .C(\u_cpu.REG_FILE._02508_ ),
    .Y(\u_cpu.REG_FILE._02509_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07202_  (.A1(\u_cpu.REG_FILE._01888_ ),
    .A2(\u_cpu.REG_FILE._02485_ ),
    .B1(\u_cpu.REG_FILE._02509_ ),
    .C1(\u_cpu.REG_FILE._02227_ ),
    .X(\u_cpu.ALU.SrcA[26] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07203_  (.A(\u_cpu.REG_FILE.rf[15][27] ),
    .B_N(\u_cpu.REG_FILE._01889_ ),
    .X(\u_cpu.REG_FILE._02510_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07204_  (.A1(\u_cpu.REG_FILE._01531_ ),
    .A2(\u_cpu.REG_FILE.rf[14][27] ),
    .B1(\u_cpu.REG_FILE._01288_ ),
    .C1(\u_cpu.REG_FILE._02510_ ),
    .Y(\u_cpu.REG_FILE._02511_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07205_  (.A1(\u_cpu.REG_FILE._01299_ ),
    .A2(\u_cpu.REG_FILE.rf[12][27] ),
    .B1_N(\u_cpu.REG_FILE._01838_ ),
    .X(\u_cpu.REG_FILE._02512_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07206_  (.A1(\u_cpu.REG_FILE._01298_ ),
    .A2(\u_cpu.REG_FILE.rf[13][27] ),
    .B1(\u_cpu.REG_FILE._02512_ ),
    .Y(\u_cpu.REG_FILE._02513_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07207_  (.A(\u_cpu.REG_FILE._02511_ ),
    .B(\u_cpu.REG_FILE._02513_ ),
    .C(\u_cpu.REG_FILE._01293_ ),
    .Y(\u_cpu.REG_FILE._02514_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07208_  (.A_N(\u_cpu.REG_FILE.rf[9][27] ),
    .B(\u_cpu.REG_FILE._01895_ ),
    .X(\u_cpu.REG_FILE._02515_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07209_  (.A1(\u_cpu.REG_FILE._02018_ ),
    .A2(\u_cpu.REG_FILE.rf[8][27] ),
    .B1_N(\u_cpu.REG_FILE._01843_ ),
    .Y(\u_cpu.REG_FILE._02516_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07210_  (.A(\u_cpu.REG_FILE.rf[11][27] ),
    .B_N(\u_cpu.REG_FILE._01345_ ),
    .X(\u_cpu.REG_FILE._02517_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07211_  (.A1(\u_cpu.REG_FILE._01620_ ),
    .A2(\u_cpu.REG_FILE.rf[10][27] ),
    .B1(\u_cpu.REG_FILE._01339_ ),
    .C1(\u_cpu.REG_FILE._02517_ ),
    .Y(\u_cpu.REG_FILE._02518_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07212_  (.A1(\u_cpu.REG_FILE._02515_ ),
    .A2(\u_cpu.REG_FILE._02516_ ),
    .B1(\u_cpu.REG_FILE._01384_ ),
    .C1(\u_cpu.REG_FILE._02518_ ),
    .Y(\u_cpu.REG_FILE._02519_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07213_  (.A(\u_cpu.REG_FILE._02514_ ),
    .B(\u_cpu.REG_FILE._02519_ ),
    .C(\u_cpu.REG_FILE._01117_ ),
    .Y(\u_cpu.REG_FILE._02520_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07214_  (.A(\u_cpu.REG_FILE.rf[5][27] ),
    .Y(\u_cpu.REG_FILE._02521_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07215_  (.A1(\u_cpu.REG_FILE._01133_ ),
    .A2(\u_cpu.REG_FILE.rf[4][27] ),
    .B1_N(\u_cpu.REG_FILE._01380_ ),
    .Y(\u_cpu.REG_FILE._02522_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07216_  (.A1(\u_cpu.REG_FILE._02521_ ),
    .A2(\u_cpu.REG_FILE._01850_ ),
    .B1(\u_cpu.REG_FILE._02522_ ),
    .Y(\u_cpu.REG_FILE._02523_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07217_  (.A1(\u_cpu.REG_FILE._01774_ ),
    .A2(\u_cpu.REG_FILE.rf[6][27] ),
    .B1(\u_cpu.REG_FILE._01400_ ),
    .Y(\u_cpu.REG_FILE._02524_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07218_  (.A_N(\u_cpu.REG_FILE.rf[7][27] ),
    .B(\u_cpu.REG_FILE._01906_ ),
    .X(\u_cpu.REG_FILE._02525_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07219_  (.A1(\u_cpu.REG_FILE._02524_ ),
    .A2(\u_cpu.REG_FILE._02525_ ),
    .B1(\u_cpu.REG_FILE._02122_ ),
    .Y(\u_cpu.REG_FILE._02526_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07220_  (.A_N(\u_cpu.REG_FILE.rf[1][27] ),
    .B(\u_cpu.REG_FILE._01161_ ),
    .X(\u_cpu.REG_FILE._02527_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07221_  (.A1(\u_cpu.REG_FILE._02105_ ),
    .A2(\u_cpu.REG_FILE.rf[0][27] ),
    .B1_N(\u_cpu.REG_FILE._01078_ ),
    .Y(\u_cpu.REG_FILE._02528_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07222_  (.A(\u_cpu.REG_FILE.rf[3][27] ),
    .B_N(\u_cpu.REG_FILE._02057_ ),
    .X(\u_cpu.REG_FILE._02529_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07223_  (.A1(\u_cpu.REG_FILE._01053_ ),
    .A2(\u_cpu.REG_FILE.rf[2][27] ),
    .B1(\u_cpu.REG_FILE._02056_ ),
    .C1(\u_cpu.REG_FILE._02529_ ),
    .Y(\u_cpu.REG_FILE._02530_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07224_  (.A1(\u_cpu.REG_FILE._02527_ ),
    .A2(\u_cpu.REG_FILE._02528_ ),
    .B1(\u_cpu.REG_FILE._01858_ ),
    .C1(\u_cpu.REG_FILE._02530_ ),
    .Y(\u_cpu.REG_FILE._02531_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07225_  (.A1(\u_cpu.REG_FILE._02523_ ),
    .A2(\u_cpu.REG_FILE._02526_ ),
    .B1(\u_cpu.REG_FILE._01414_ ),
    .C1(\u_cpu.REG_FILE._02531_ ),
    .Y(\u_cpu.REG_FILE._02532_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._07226_  (.A(\u_cpu.REG_FILE._02520_ ),
    .B(\u_cpu.REG_FILE._02532_ ),
    .Y(\u_cpu.REG_FILE._02533_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07227_  (.A(\u_cpu.REG_FILE.rf[27][27] ),
    .B_N(\u_cpu.REG_FILE._01528_ ),
    .X(\u_cpu.REG_FILE._02534_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07228_  (.A1(\u_cpu.REG_FILE._01308_ ),
    .A2(\u_cpu.REG_FILE.rf[26][27] ),
    .B1(\u_cpu.REG_FILE._01660_ ),
    .C1(\u_cpu.REG_FILE._02534_ ),
    .X(\u_cpu.REG_FILE._02535_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07229_  (.A1(\u_cpu.REG_FILE._01447_ ),
    .A2(\u_cpu.REG_FILE.rf[24][27] ),
    .B1_N(\u_cpu.REG_FILE._01062_ ),
    .X(\u_cpu.REG_FILE._02536_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07230_  (.A(\u_cpu.REG_FILE.rf[25][27] ),
    .B_N(\u_cpu.REG_FILE._01194_ ),
    .X(\u_cpu.REG_FILE._02537_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._07231_  (.A1(\u_cpu.REG_FILE._02536_ ),
    .A2(\u_cpu.REG_FILE._02537_ ),
    .B1(\u_cpu.REG_FILE._01196_ ),
    .X(\u_cpu.REG_FILE._02538_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07232_  (.A(\u_cpu.REG_FILE._02010_ ),
    .B(\u_cpu.REG_FILE.rf[30][27] ),
    .Y(\u_cpu.REG_FILE._02539_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07233_  (.A1(\u_cpu.REG_FILE.rf[31][27] ),
    .A2(\u_cpu.REG_FILE._01969_ ),
    .B1(\u_cpu.REG_FILE._01501_ ),
    .Y(\u_cpu.REG_FILE._02540_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07234_  (.A1(\u_cpu.REG_FILE._01503_ ),
    .A2(\u_cpu.REG_FILE.rf[28][27] ),
    .B1_N(\u_cpu.REG_FILE._01098_ ),
    .X(\u_cpu.REG_FILE._02541_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07235_  (.A1(\u_cpu.REG_FILE._01668_ ),
    .A2(\u_cpu.REG_FILE.rf[29][27] ),
    .B1(\u_cpu.REG_FILE._02541_ ),
    .Y(\u_cpu.REG_FILE._02542_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07236_  (.A1(\u_cpu.REG_FILE._02539_ ),
    .A2(\u_cpu.REG_FILE._02540_ ),
    .B1(\u_cpu.REG_FILE._02542_ ),
    .C1(\u_cpu.REG_FILE._02016_ ),
    .Y(\u_cpu.REG_FILE._02543_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07237_  (.A1(\u_cpu.REG_FILE._02535_ ),
    .A2(\u_cpu.REG_FILE._02538_ ),
    .B1(\u_cpu.REG_FILE._01869_ ),
    .C1(\u_cpu.REG_FILE._02543_ ),
    .Y(\u_cpu.REG_FILE._02544_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07238_  (.A(\u_cpu.REG_FILE._01379_ ),
    .B(\u_cpu.REG_FILE.rf[16][27] ),
    .Y(\u_cpu.REG_FILE._02545_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07239_  (.A_N(\u_cpu.REG_FILE.rf[17][27] ),
    .B(\u_cpu.REG_FILE._01029_ ),
    .X(\u_cpu.REG_FILE._02546_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.REG_FILE._07240_  (.A1(\u_cpu.REG_FILE._01060_ ),
    .A2(\u_cpu.REG_FILE.rf[18][27] ),
    .B1(\u_cpu.REG_FILE._01239_ ),
    .X(\u_cpu.REG_FILE._02547_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07241_  (.A1(\u_cpu.REG_FILE.rf[19][27] ),
    .A2(\u_cpu.REG_FILE._01329_ ),
    .B1(\u_cpu.REG_FILE._02547_ ),
    .Y(\u_cpu.REG_FILE._02548_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._07242_  (.A1(\u_cpu.REG_FILE._01033_ ),
    .A2(\u_cpu.REG_FILE._02545_ ),
    .A3(\u_cpu.REG_FILE._02546_ ),
    .B1(\u_cpu.REG_FILE._01058_ ),
    .C1(\u_cpu.REG_FILE._02548_ ),
    .Y(\u_cpu.REG_FILE._02549_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._07243_  (.A(\u_cpu.REG_FILE._01324_ ),
    .B(\u_cpu.REG_FILE.rf[22][27] ),
    .X(\u_cpu.REG_FILE._02550_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07244_  (.A1(\u_cpu.REG_FILE._01321_ ),
    .A2(\u_cpu.REG_FILE.rf[23][27] ),
    .B1(\u_cpu.REG_FILE._01063_ ),
    .C1(\u_cpu.REG_FILE._02550_ ),
    .Y(\u_cpu.REG_FILE._02551_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07245_  (.A1(\u_cpu.REG_FILE._01632_ ),
    .A2(\u_cpu.REG_FILE.rf[20][27] ),
    .B1_N(\u_cpu.REG_FILE._01134_ ),
    .X(\u_cpu.REG_FILE._02552_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07246_  (.A1(\u_cpu.REG_FILE._01120_ ),
    .A2(\u_cpu.REG_FILE.rf[21][27] ),
    .B1(\u_cpu.REG_FILE._02552_ ),
    .Y(\u_cpu.REG_FILE._02553_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07247_  (.A(\u_cpu.REG_FILE._02551_ ),
    .B(\u_cpu.REG_FILE._02553_ ),
    .C(\u_cpu.REG_FILE._01552_ ),
    .Y(\u_cpu.REG_FILE._02554_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07248_  (.A(\u_cpu.REG_FILE._01569_ ),
    .B(\u_cpu.REG_FILE._02549_ ),
    .C(\u_cpu.REG_FILE._02554_ ),
    .Y(\u_cpu.REG_FILE._02555_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07249_  (.A(\u_cpu.REG_FILE._02544_ ),
    .B(\u_cpu.REG_FILE._02555_ ),
    .C(\u_cpu.REG_FILE._01025_ ),
    .Y(\u_cpu.REG_FILE._02556_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07250_  (.A1(\u_cpu.REG_FILE._01888_ ),
    .A2(\u_cpu.REG_FILE._02533_ ),
    .B1(\u_cpu.REG_FILE._02556_ ),
    .C1(\u_cpu.REG_FILE._02227_ ),
    .X(\u_cpu.ALU.SrcA[27] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07251_  (.A(\u_cpu.REG_FILE.rf[15][28] ),
    .B_N(\u_cpu.REG_FILE._01889_ ),
    .X(\u_cpu.REG_FILE._02557_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07252_  (.A1(\u_cpu.REG_FILE._01531_ ),
    .A2(\u_cpu.REG_FILE.rf[14][28] ),
    .B1(\u_cpu.REG_FILE._01288_ ),
    .C1(\u_cpu.REG_FILE._02557_ ),
    .Y(\u_cpu.REG_FILE._02558_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07253_  (.A1(\u_cpu.REG_FILE._01299_ ),
    .A2(\u_cpu.REG_FILE.rf[12][28] ),
    .B1_N(\u_cpu.REG_FILE._01106_ ),
    .X(\u_cpu.REG_FILE._02559_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07254_  (.A1(\u_cpu.REG_FILE._01298_ ),
    .A2(\u_cpu.REG_FILE.rf[13][28] ),
    .B1(\u_cpu.REG_FILE._02559_ ),
    .Y(\u_cpu.REG_FILE._02560_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07255_  (.A(\u_cpu.REG_FILE._02558_ ),
    .B(\u_cpu.REG_FILE._02560_ ),
    .C(\u_cpu.REG_FILE._01293_ ),
    .Y(\u_cpu.REG_FILE._02561_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07256_  (.A_N(\u_cpu.REG_FILE.rf[9][28] ),
    .B(\u_cpu.REG_FILE._01895_ ),
    .X(\u_cpu.REG_FILE._02562_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07257_  (.A1(\u_cpu.REG_FILE._02018_ ),
    .A2(\u_cpu.REG_FILE.rf[8][28] ),
    .B1_N(\u_cpu.REG_FILE._01521_ ),
    .Y(\u_cpu.REG_FILE._02563_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07258_  (.A(\u_cpu.REG_FILE.rf[11][28] ),
    .B_N(\u_cpu.REG_FILE._01345_ ),
    .X(\u_cpu.REG_FILE._02564_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07259_  (.A1(\u_cpu.REG_FILE._01620_ ),
    .A2(\u_cpu.REG_FILE.rf[10][28] ),
    .B1(\u_cpu.REG_FILE._01339_ ),
    .C1(\u_cpu.REG_FILE._02564_ ),
    .Y(\u_cpu.REG_FILE._02565_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07260_  (.A1(\u_cpu.REG_FILE._02562_ ),
    .A2(\u_cpu.REG_FILE._02563_ ),
    .B1(\u_cpu.REG_FILE._01384_ ),
    .C1(\u_cpu.REG_FILE._02565_ ),
    .Y(\u_cpu.REG_FILE._02566_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07261_  (.A(\u_cpu.REG_FILE._02561_ ),
    .B(\u_cpu.REG_FILE._02566_ ),
    .C(\u_cpu.REG_FILE._01117_ ),
    .Y(\u_cpu.REG_FILE._02567_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07262_  (.A(\u_cpu.REG_FILE.rf[5][28] ),
    .Y(\u_cpu.REG_FILE._02568_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07263_  (.A1(\u_cpu.REG_FILE._01133_ ),
    .A2(\u_cpu.REG_FILE.rf[4][28] ),
    .B1_N(\u_cpu.REG_FILE._01380_ ),
    .Y(\u_cpu.REG_FILE._02569_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07264_  (.A1(\u_cpu.REG_FILE._02568_ ),
    .A2(\u_cpu.REG_FILE._01284_ ),
    .B1(\u_cpu.REG_FILE._02569_ ),
    .Y(\u_cpu.REG_FILE._02570_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07265_  (.A1(\u_cpu.REG_FILE._01774_ ),
    .A2(\u_cpu.REG_FILE.rf[6][28] ),
    .B1(\u_cpu.REG_FILE._01400_ ),
    .Y(\u_cpu.REG_FILE._02571_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07266_  (.A_N(\u_cpu.REG_FILE.rf[7][28] ),
    .B(\u_cpu.REG_FILE._01906_ ),
    .X(\u_cpu.REG_FILE._02572_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07267_  (.A1(\u_cpu.REG_FILE._02571_ ),
    .A2(\u_cpu.REG_FILE._02572_ ),
    .B1(\u_cpu.REG_FILE._02122_ ),
    .Y(\u_cpu.REG_FILE._02573_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07268_  (.A_N(\u_cpu.REG_FILE.rf[1][28] ),
    .B(\u_cpu.REG_FILE._01161_ ),
    .X(\u_cpu.REG_FILE._02574_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07269_  (.A1(\u_cpu.REG_FILE._02105_ ),
    .A2(\u_cpu.REG_FILE.rf[0][28] ),
    .B1_N(\u_cpu.REG_FILE._01078_ ),
    .Y(\u_cpu.REG_FILE._02575_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07270_  (.A(\u_cpu.REG_FILE.rf[3][28] ),
    .B_N(\u_cpu.REG_FILE._02057_ ),
    .X(\u_cpu.REG_FILE._02576_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07271_  (.A1(\u_cpu.REG_FILE._01053_ ),
    .A2(\u_cpu.REG_FILE.rf[2][28] ),
    .B1(\u_cpu.REG_FILE._02056_ ),
    .C1(\u_cpu.REG_FILE._02576_ ),
    .Y(\u_cpu.REG_FILE._02577_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07272_  (.A1(\u_cpu.REG_FILE._02574_ ),
    .A2(\u_cpu.REG_FILE._02575_ ),
    .B1(\u_cpu.REG_FILE._01139_ ),
    .C1(\u_cpu.REG_FILE._02577_ ),
    .Y(\u_cpu.REG_FILE._02578_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07273_  (.A1(\u_cpu.REG_FILE._02570_ ),
    .A2(\u_cpu.REG_FILE._02573_ ),
    .B1(\u_cpu.REG_FILE._01414_ ),
    .C1(\u_cpu.REG_FILE._02578_ ),
    .Y(\u_cpu.REG_FILE._02579_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._07274_  (.A(\u_cpu.REG_FILE._02567_ ),
    .B(\u_cpu.REG_FILE._02579_ ),
    .Y(\u_cpu.REG_FILE._02580_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07275_  (.A1(\u_cpu.REG_FILE._01081_ ),
    .A2(\u_cpu.REG_FILE.rf[24][28] ),
    .B1_N(\u_cpu.REG_FILE._01611_ ),
    .Y(\u_cpu.REG_FILE._02581_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07276_  (.A_N(\u_cpu.REG_FILE.rf[25][28] ),
    .B(\u_cpu.REG_FILE._01750_ ),
    .X(\u_cpu.REG_FILE._02582_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07277_  (.A1(\u_cpu.REG_FILE._02581_ ),
    .A2(\u_cpu.REG_FILE._02582_ ),
    .B1(\u_cpu.REG_FILE._01814_ ),
    .Y(\u_cpu.REG_FILE._02583_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._07278_  (.A(\u_cpu.REG_FILE._01340_ ),
    .B(\u_cpu.REG_FILE.rf[26][28] ),
    .X(\u_cpu.REG_FILE._02584_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07279_  (.A1(\u_cpu.REG_FILE._01124_ ),
    .A2(\u_cpu.REG_FILE.rf[27][28] ),
    .B1(\u_cpu.REG_FILE._01121_ ),
    .C1(\u_cpu.REG_FILE._02584_ ),
    .X(\u_cpu.REG_FILE._02585_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07280_  (.A(\u_cpu.REG_FILE._02010_ ),
    .B(\u_cpu.REG_FILE.rf[30][28] ),
    .Y(\u_cpu.REG_FILE._02586_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07281_  (.A1(\u_cpu.REG_FILE.rf[31][28] ),
    .A2(\u_cpu.REG_FILE._01969_ ),
    .B1(\u_cpu.REG_FILE._01107_ ),
    .Y(\u_cpu.REG_FILE._02587_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07282_  (.A1(\u_cpu.REG_FILE._02013_ ),
    .A2(\u_cpu.REG_FILE.rf[28][28] ),
    .B1_N(\u_cpu.REG_FILE._01098_ ),
    .X(\u_cpu.REG_FILE._02588_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07283_  (.A1(\u_cpu.REG_FILE._01668_ ),
    .A2(\u_cpu.REG_FILE.rf[29][28] ),
    .B1(\u_cpu.REG_FILE._02588_ ),
    .Y(\u_cpu.REG_FILE._02589_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07284_  (.A1(\u_cpu.REG_FILE._02586_ ),
    .A2(\u_cpu.REG_FILE._02587_ ),
    .B1(\u_cpu.REG_FILE._02589_ ),
    .C1(\u_cpu.REG_FILE._02016_ ),
    .Y(\u_cpu.REG_FILE._02590_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07285_  (.A1(\u_cpu.REG_FILE._02583_ ),
    .A2(\u_cpu.REG_FILE._02585_ ),
    .B1(\u_cpu.REG_FILE._01869_ ),
    .C1(\u_cpu.REG_FILE._02590_ ),
    .Y(\u_cpu.REG_FILE._02591_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07286_  (.A(\u_cpu.REG_FILE.rf[19][28] ),
    .Y(\u_cpu.REG_FILE._02592_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07287_  (.A1(\u_cpu.REG_FILE._01523_ ),
    .A2(\u_cpu.REG_FILE.rf[18][28] ),
    .B1(\u_cpu.REG_FILE._01533_ ),
    .Y(\u_cpu.REG_FILE._02593_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07288_  (.A1(\u_cpu.REG_FILE._02592_ ),
    .A2(\u_cpu.REG_FILE._01399_ ),
    .B1(\u_cpu.REG_FILE._02593_ ),
    .Y(\u_cpu.REG_FILE._02594_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07289_  (.A(\u_cpu.REG_FILE.rf[17][28] ),
    .Y(\u_cpu.REG_FILE._02595_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07290_  (.A1(\u_cpu.REG_FILE._01404_ ),
    .A2(\u_cpu.REG_FILE.rf[16][28] ),
    .B1_N(\u_cpu.REG_FILE._01258_ ),
    .Y(\u_cpu.REG_FILE._02596_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07291_  (.A1(\u_cpu.REG_FILE._02595_ ),
    .A2(\u_cpu.REG_FILE._01399_ ),
    .B1(\u_cpu.REG_FILE._02596_ ),
    .Y(\u_cpu.REG_FILE._02597_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07292_  (.A(\u_cpu.REG_FILE.rf[23][28] ),
    .B_N(\u_cpu.REG_FILE._01408_ ),
    .X(\u_cpu.REG_FILE._02598_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07293_  (.A1(\u_cpu.REG_FILE._01077_ ),
    .A2(\u_cpu.REG_FILE.rf[22][28] ),
    .B1(\u_cpu.REG_FILE._01407_ ),
    .C1(\u_cpu.REG_FILE._02598_ ),
    .Y(\u_cpu.REG_FILE._02599_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07294_  (.A1(\u_cpu.REG_FILE._01324_ ),
    .A2(\u_cpu.REG_FILE.rf[20][28] ),
    .B1_N(\u_cpu.REG_FILE._01304_ ),
    .X(\u_cpu.REG_FILE._02600_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07295_  (.A1(\u_cpu.REG_FILE._01038_ ),
    .A2(\u_cpu.REG_FILE.rf[21][28] ),
    .B1(\u_cpu.REG_FILE._02600_ ),
    .Y(\u_cpu.REG_FILE._02601_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07296_  (.A(\u_cpu.REG_FILE._02599_ ),
    .B(\u_cpu.REG_FILE._02601_ ),
    .C(\u_cpu.REG_FILE._01115_ ),
    .Y(\u_cpu.REG_FILE._02602_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._07297_  (.A1(\u_cpu.REG_FILE._01047_ ),
    .A2(\u_cpu.REG_FILE._02594_ ),
    .A3(\u_cpu.REG_FILE._02597_ ),
    .B1(\u_cpu.REG_FILE._02602_ ),
    .C1(\u_cpu.REG_FILE._01089_ ),
    .Y(\u_cpu.REG_FILE._02603_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07298_  (.A(\u_cpu.REG_FILE._02591_ ),
    .B(\u_cpu.REG_FILE._02603_ ),
    .C(\u_cpu.REG_FILE._01025_ ),
    .Y(\u_cpu.REG_FILE._02604_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07299_  (.A1(\u_cpu.REG_FILE._01888_ ),
    .A2(\u_cpu.REG_FILE._02580_ ),
    .B1(\u_cpu.REG_FILE._02604_ ),
    .C1(\u_cpu.REG_FILE._02227_ ),
    .X(\u_cpu.ALU.SrcA[28] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07300_  (.A(\u_cpu.REG_FILE.rf[15][29] ),
    .B_N(\u_cpu.REG_FILE._01262_ ),
    .X(\u_cpu.REG_FILE._02605_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07301_  (.A1(\u_cpu.REG_FILE._01531_ ),
    .A2(\u_cpu.REG_FILE.rf[14][29] ),
    .B1(\u_cpu.REG_FILE._01288_ ),
    .C1(\u_cpu.REG_FILE._02605_ ),
    .Y(\u_cpu.REG_FILE._02606_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07302_  (.A1(\u_cpu.REG_FILE._01299_ ),
    .A2(\u_cpu.REG_FILE.rf[12][29] ),
    .B1_N(\u_cpu.REG_FILE._01106_ ),
    .X(\u_cpu.REG_FILE._02607_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07303_  (.A1(\u_cpu.REG_FILE._01298_ ),
    .A2(\u_cpu.REG_FILE.rf[13][29] ),
    .B1(\u_cpu.REG_FILE._02607_ ),
    .Y(\u_cpu.REG_FILE._02608_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07304_  (.A(\u_cpu.REG_FILE._02606_ ),
    .B(\u_cpu.REG_FILE._02608_ ),
    .C(\u_cpu.REG_FILE._01293_ ),
    .Y(\u_cpu.REG_FILE._02609_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07305_  (.A_N(\u_cpu.REG_FILE.rf[9][29] ),
    .B(\u_cpu.REG_FILE._01382_ ),
    .X(\u_cpu.REG_FILE._02610_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07306_  (.A1(\u_cpu.REG_FILE._02018_ ),
    .A2(\u_cpu.REG_FILE.rf[8][29] ),
    .B1_N(\u_cpu.REG_FILE._01521_ ),
    .Y(\u_cpu.REG_FILE._02611_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07307_  (.A(\u_cpu.REG_FILE.rf[11][29] ),
    .B_N(\u_cpu.REG_FILE._01345_ ),
    .X(\u_cpu.REG_FILE._02612_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07308_  (.A1(\u_cpu.REG_FILE._01620_ ),
    .A2(\u_cpu.REG_FILE.rf[10][29] ),
    .B1(\u_cpu.REG_FILE._01339_ ),
    .C1(\u_cpu.REG_FILE._02612_ ),
    .Y(\u_cpu.REG_FILE._02613_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07309_  (.A1(\u_cpu.REG_FILE._02610_ ),
    .A2(\u_cpu.REG_FILE._02611_ ),
    .B1(\u_cpu.REG_FILE._01384_ ),
    .C1(\u_cpu.REG_FILE._02613_ ),
    .Y(\u_cpu.REG_FILE._02614_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07310_  (.A(\u_cpu.REG_FILE._02609_ ),
    .B(\u_cpu.REG_FILE._02614_ ),
    .C(\u_cpu.REG_FILE._01117_ ),
    .Y(\u_cpu.REG_FILE._02615_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07311_  (.A(\u_cpu.REG_FILE.rf[5][29] ),
    .Y(\u_cpu.REG_FILE._02616_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07312_  (.A1(\u_cpu.REG_FILE._01133_ ),
    .A2(\u_cpu.REG_FILE.rf[4][29] ),
    .B1_N(\u_cpu.REG_FILE._01380_ ),
    .Y(\u_cpu.REG_FILE._02617_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07313_  (.A1(\u_cpu.REG_FILE._02616_ ),
    .A2(\u_cpu.REG_FILE._01284_ ),
    .B1(\u_cpu.REG_FILE._02617_ ),
    .Y(\u_cpu.REG_FILE._02618_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07314_  (.A1(\u_cpu.REG_FILE._01774_ ),
    .A2(\u_cpu.REG_FILE.rf[6][29] ),
    .B1(\u_cpu.REG_FILE._01400_ ),
    .Y(\u_cpu.REG_FILE._02619_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07315_  (.A_N(\u_cpu.REG_FILE.rf[7][29] ),
    .B(\u_cpu.REG_FILE._01091_ ),
    .X(\u_cpu.REG_FILE._02620_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07316_  (.A1(\u_cpu.REG_FILE._02619_ ),
    .A2(\u_cpu.REG_FILE._02620_ ),
    .B1(\u_cpu.REG_FILE._02122_ ),
    .Y(\u_cpu.REG_FILE._02621_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07317_  (.A_N(\u_cpu.REG_FILE.rf[1][29] ),
    .B(\u_cpu.REG_FILE._01161_ ),
    .X(\u_cpu.REG_FILE._02622_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07318_  (.A1(\u_cpu.REG_FILE._02105_ ),
    .A2(\u_cpu.REG_FILE.rf[0][29] ),
    .B1_N(\u_cpu.REG_FILE._01078_ ),
    .Y(\u_cpu.REG_FILE._02623_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07319_  (.A(\u_cpu.REG_FILE.rf[3][29] ),
    .B_N(\u_cpu.REG_FILE._02057_ ),
    .X(\u_cpu.REG_FILE._02624_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07320_  (.A1(\u_cpu.REG_FILE._01053_ ),
    .A2(\u_cpu.REG_FILE.rf[2][29] ),
    .B1(\u_cpu.REG_FILE._02056_ ),
    .C1(\u_cpu.REG_FILE._02624_ ),
    .Y(\u_cpu.REG_FILE._02625_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07321_  (.A1(\u_cpu.REG_FILE._02622_ ),
    .A2(\u_cpu.REG_FILE._02623_ ),
    .B1(\u_cpu.REG_FILE._01139_ ),
    .C1(\u_cpu.REG_FILE._02625_ ),
    .Y(\u_cpu.REG_FILE._02626_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07322_  (.A1(\u_cpu.REG_FILE._02618_ ),
    .A2(\u_cpu.REG_FILE._02621_ ),
    .B1(\u_cpu.REG_FILE._01414_ ),
    .C1(\u_cpu.REG_FILE._02626_ ),
    .Y(\u_cpu.REG_FILE._02627_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._07323_  (.A(\u_cpu.REG_FILE._02615_ ),
    .B(\u_cpu.REG_FILE._02627_ ),
    .Y(\u_cpu.REG_FILE._02628_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07324_  (.A(\u_cpu.REG_FILE.rf[27][29] ),
    .B_N(\u_cpu.REG_FILE._01528_ ),
    .X(\u_cpu.REG_FILE._02629_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07325_  (.A1(\u_cpu.REG_FILE._01308_ ),
    .A2(\u_cpu.REG_FILE.rf[26][29] ),
    .B1(\u_cpu.REG_FILE._01660_ ),
    .C1(\u_cpu.REG_FILE._02629_ ),
    .X(\u_cpu.REG_FILE._02630_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07326_  (.A1(\u_cpu.REG_FILE._01447_ ),
    .A2(\u_cpu.REG_FILE.rf[24][29] ),
    .B1_N(\u_cpu.REG_FILE._01062_ ),
    .X(\u_cpu.REG_FILE._02631_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07327_  (.A(\u_cpu.REG_FILE.rf[25][29] ),
    .B_N(\u_cpu.REG_FILE._01125_ ),
    .X(\u_cpu.REG_FILE._02632_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._07328_  (.A1(\u_cpu.REG_FILE._02631_ ),
    .A2(\u_cpu.REG_FILE._02632_ ),
    .B1(\u_cpu.REG_FILE._01046_ ),
    .X(\u_cpu.REG_FILE._02633_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07329_  (.A(\u_cpu.REG_FILE._02010_ ),
    .B(\u_cpu.REG_FILE.rf[30][29] ),
    .Y(\u_cpu.REG_FILE._02634_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07330_  (.A1(\u_cpu.REG_FILE.rf[31][29] ),
    .A2(\u_cpu.REG_FILE._01969_ ),
    .B1(\u_cpu.REG_FILE._01107_ ),
    .Y(\u_cpu.REG_FILE._02635_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07331_  (.A1(\u_cpu.REG_FILE._02013_ ),
    .A2(\u_cpu.REG_FILE.rf[28][29] ),
    .B1_N(\u_cpu.REG_FILE._01098_ ),
    .X(\u_cpu.REG_FILE._02636_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07332_  (.A1(\u_cpu.REG_FILE._01668_ ),
    .A2(\u_cpu.REG_FILE.rf[29][29] ),
    .B1(\u_cpu.REG_FILE._02636_ ),
    .Y(\u_cpu.REG_FILE._02637_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07333_  (.A1(\u_cpu.REG_FILE._02634_ ),
    .A2(\u_cpu.REG_FILE._02635_ ),
    .B1(\u_cpu.REG_FILE._02637_ ),
    .C1(\u_cpu.REG_FILE._02016_ ),
    .Y(\u_cpu.REG_FILE._02638_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07334_  (.A1(\u_cpu.REG_FILE._02630_ ),
    .A2(\u_cpu.REG_FILE._02633_ ),
    .B1(\u_cpu.REG_FILE._01869_ ),
    .C1(\u_cpu.REG_FILE._02638_ ),
    .Y(\u_cpu.REG_FILE._02639_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07335_  (.A1(\u_cpu.REG_FILE._01206_ ),
    .A2(\u_cpu.REG_FILE.rf[18][29] ),
    .B1(\u_cpu.REG_FILE._01407_ ),
    .Y(\u_cpu.REG_FILE._02640_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07336_  (.A(\u_cpu.REG_FILE.rf[19][29] ),
    .B(\u_cpu.REG_FILE._01509_ ),
    .Y(\u_cpu.REG_FILE._02641_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07337_  (.A1(\u_cpu.REG_FILE._01152_ ),
    .A2(\u_cpu.REG_FILE.rf[16][29] ),
    .B1_N(\u_cpu.REG_FILE._01153_ ),
    .X(\u_cpu.REG_FILE._02642_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07338_  (.A1(\u_cpu.REG_FILE._01726_ ),
    .A2(\u_cpu.REG_FILE.rf[17][29] ),
    .B1(\u_cpu.REG_FILE._02642_ ),
    .Y(\u_cpu.REG_FILE._02643_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07339_  (.A1(\u_cpu.REG_FILE._02640_ ),
    .A2(\u_cpu.REG_FILE._02641_ ),
    .B1(\u_cpu.REG_FILE._01264_ ),
    .C1(\u_cpu.REG_FILE._02643_ ),
    .Y(\u_cpu.REG_FILE._02644_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._07340_  (.A(\u_cpu.REG_FILE._01324_ ),
    .B(\u_cpu.REG_FILE.rf[22][29] ),
    .X(\u_cpu.REG_FILE._02645_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07341_  (.A1(\u_cpu.REG_FILE._01321_ ),
    .A2(\u_cpu.REG_FILE.rf[23][29] ),
    .B1(\u_cpu.REG_FILE._01063_ ),
    .C1(\u_cpu.REG_FILE._02645_ ),
    .Y(\u_cpu.REG_FILE._02646_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07342_  (.A1(\u_cpu.REG_FILE._01632_ ),
    .A2(\u_cpu.REG_FILE.rf[20][29] ),
    .B1_N(\u_cpu.REG_FILE._01134_ ),
    .X(\u_cpu.REG_FILE._02647_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07343_  (.A1(\u_cpu.REG_FILE._01120_ ),
    .A2(\u_cpu.REG_FILE.rf[21][29] ),
    .B1(\u_cpu.REG_FILE._02647_ ),
    .Y(\u_cpu.REG_FILE._02648_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07344_  (.A(\u_cpu.REG_FILE._02646_ ),
    .B(\u_cpu.REG_FILE._02648_ ),
    .C(\u_cpu.REG_FILE._01552_ ),
    .Y(\u_cpu.REG_FILE._02649_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07345_  (.A(\u_cpu.REG_FILE._01541_ ),
    .B(\u_cpu.REG_FILE._02644_ ),
    .C(\u_cpu.REG_FILE._02649_ ),
    .Y(\u_cpu.REG_FILE._02650_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07346_  (.A(\u_cpu.REG_FILE._02639_ ),
    .B(\u_cpu.REG_FILE._02650_ ),
    .C(\u_cpu.REG_FILE._01025_ ),
    .Y(\u_cpu.REG_FILE._02651_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07347_  (.A1(\u_cpu.REG_FILE._01159_ ),
    .A2(\u_cpu.REG_FILE._02628_ ),
    .B1(\u_cpu.REG_FILE._02651_ ),
    .C1(\u_cpu.REG_FILE._02227_ ),
    .X(\u_cpu.ALU.SrcA[29] ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07348_  (.A1(\u_cpu.REG_FILE._01184_ ),
    .A2(\u_cpu.REG_FILE.rf[8][30] ),
    .B1_N(\u_cpu.REG_FILE._01094_ ),
    .Y(\u_cpu.REG_FILE._02652_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07349_  (.A_N(\u_cpu.REG_FILE.rf[9][30] ),
    .B(\u_cpu.REG_FILE._01074_ ),
    .X(\u_cpu.REG_FILE._02653_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07350_  (.A1(\u_cpu.REG_FILE._02652_ ),
    .A2(\u_cpu.REG_FILE._02653_ ),
    .B1(\u_cpu.REG_FILE._01525_ ),
    .Y(\u_cpu.REG_FILE._02654_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._07351_  (.A(\u_cpu.REG_FILE._01528_ ),
    .B(\u_cpu.REG_FILE.rf[10][30] ),
    .X(\u_cpu.REG_FILE._02655_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07352_  (.A1(\u_cpu.REG_FILE._01137_ ),
    .A2(\u_cpu.REG_FILE.rf[11][30] ),
    .B1(\u_cpu.REG_FILE._01387_ ),
    .C1(\u_cpu.REG_FILE._02655_ ),
    .X(\u_cpu.REG_FILE._02656_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07353_  (.A(\u_cpu.REG_FILE._01118_ ),
    .B(\u_cpu.REG_FILE.rf[12][30] ),
    .Y(\u_cpu.REG_FILE._02657_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07354_  (.A1(\u_cpu.REG_FILE.rf[13][30] ),
    .A2(\u_cpu.REG_FILE._01535_ ),
    .B1_N(\u_cpu.REG_FILE._01305_ ),
    .Y(\u_cpu.REG_FILE._02658_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._07355_  (.A(\u_cpu.REG_FILE._01536_ ),
    .B(\u_cpu.REG_FILE.rf[14][30] ),
    .X(\u_cpu.REG_FILE._02659_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07356_  (.A1(\u_cpu.REG_FILE._01535_ ),
    .A2(\u_cpu.REG_FILE.rf[15][30] ),
    .B1(\u_cpu.REG_FILE._01527_ ),
    .C1(\u_cpu.REG_FILE._02659_ ),
    .Y(\u_cpu.REG_FILE._02660_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07357_  (.A1(\u_cpu.REG_FILE._02657_ ),
    .A2(\u_cpu.REG_FILE._02658_ ),
    .B1(\u_cpu.REG_FILE._01129_ ),
    .C1(\u_cpu.REG_FILE._02660_ ),
    .Y(\u_cpu.REG_FILE._02661_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07358_  (.A1(\u_cpu.REG_FILE._02654_ ),
    .A2(\u_cpu.REG_FILE._02656_ ),
    .B1(\u_cpu.REG_FILE._01117_ ),
    .C1(\u_cpu.REG_FILE._02661_ ),
    .X(\u_cpu.REG_FILE._02662_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07359_  (.A_N(\u_cpu.REG_FILE.rf[1][30] ),
    .B(\u_cpu.REG_FILE._01547_ ),
    .X(\u_cpu.REG_FILE._02663_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07360_  (.A1(\u_cpu.REG_FILE._01549_ ),
    .A2(\u_cpu.REG_FILE.rf[0][30] ),
    .B1_N(\u_cpu.REG_FILE._01550_ ),
    .Y(\u_cpu.REG_FILE._02664_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07361_  (.A(\u_cpu.REG_FILE.rf[3][30] ),
    .B_N(\u_cpu.REG_FILE._01065_ ),
    .X(\u_cpu.REG_FILE._02665_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07362_  (.A1(\u_cpu.REG_FILE._01061_ ),
    .A2(\u_cpu.REG_FILE.rf[2][30] ),
    .B1(\u_cpu.REG_FILE._01147_ ),
    .C1(\u_cpu.REG_FILE._02665_ ),
    .Y(\u_cpu.REG_FILE._02666_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07363_  (.A1(\u_cpu.REG_FILE._02663_ ),
    .A2(\u_cpu.REG_FILE._02664_ ),
    .B1(\u_cpu.REG_FILE._01059_ ),
    .C1(\u_cpu.REG_FILE._02666_ ),
    .Y(\u_cpu.REG_FILE._02667_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07364_  (.A_N(\u_cpu.REG_FILE.rf[5][30] ),
    .B(\u_cpu.REG_FILE._01547_ ),
    .X(\u_cpu.REG_FILE._02668_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07365_  (.A1(\u_cpu.REG_FILE._01549_ ),
    .A2(\u_cpu.REG_FILE.rf[4][30] ),
    .B1_N(\u_cpu.REG_FILE._01055_ ),
    .Y(\u_cpu.REG_FILE._02669_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.REG_FILE._07366_  (.A1(\u_cpu.REG_FILE._01262_ ),
    .A2(\u_cpu.REG_FILE.rf[6][30] ),
    .B1(\u_cpu.REG_FILE._01553_ ),
    .X(\u_cpu.REG_FILE._02670_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07367_  (.A1(\u_cpu.REG_FILE.rf[7][30] ),
    .A2(\u_cpu.REG_FILE._01287_ ),
    .B1(\u_cpu.REG_FILE._02670_ ),
    .Y(\u_cpu.REG_FILE._02671_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07368_  (.A1(\u_cpu.REG_FILE._02668_ ),
    .A2(\u_cpu.REG_FILE._02669_ ),
    .B1(\u_cpu.REG_FILE._01087_ ),
    .C1(\u_cpu.REG_FILE._02671_ ),
    .Y(\u_cpu.REG_FILE._02672_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._07369_  (.A1(\u_cpu.REG_FILE._01541_ ),
    .A2(\u_cpu.REG_FILE._02667_ ),
    .A3(\u_cpu.REG_FILE._02672_ ),
    .B1(\u_cpu.REG_FILE._01024_ ),
    .X(\u_cpu.REG_FILE._02673_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07370_  (.A1(\u_cpu.REG_FILE._01081_ ),
    .A2(\u_cpu.REG_FILE.rf[24][30] ),
    .B1_N(\u_cpu.REG_FILE._01611_ ),
    .Y(\u_cpu.REG_FILE._02674_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07371_  (.A_N(\u_cpu.REG_FILE.rf[25][30] ),
    .B(\u_cpu.REG_FILE._01750_ ),
    .X(\u_cpu.REG_FILE._02675_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07372_  (.A1(\u_cpu.REG_FILE._02674_ ),
    .A2(\u_cpu.REG_FILE._02675_ ),
    .B1(\u_cpu.REG_FILE._01814_ ),
    .Y(\u_cpu.REG_FILE._02676_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._07373_  (.A(\u_cpu.REG_FILE._01310_ ),
    .B(\u_cpu.REG_FILE.rf[26][30] ),
    .X(\u_cpu.REG_FILE._02677_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07374_  (.A1(\u_cpu.REG_FILE._01124_ ),
    .A2(\u_cpu.REG_FILE.rf[27][30] ),
    .B1(\u_cpu.REG_FILE._01121_ ),
    .C1(\u_cpu.REG_FILE._02677_ ),
    .X(\u_cpu.REG_FILE._02678_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07375_  (.A(\u_cpu.REG_FILE._02010_ ),
    .B(\u_cpu.REG_FILE.rf[30][30] ),
    .Y(\u_cpu.REG_FILE._02679_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07376_  (.A1(\u_cpu.REG_FILE.rf[31][30] ),
    .A2(\u_cpu.REG_FILE._01969_ ),
    .B1(\u_cpu.REG_FILE._01107_ ),
    .Y(\u_cpu.REG_FILE._02680_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07377_  (.A1(\u_cpu.REG_FILE._02013_ ),
    .A2(\u_cpu.REG_FILE.rf[28][30] ),
    .B1_N(\u_cpu.REG_FILE._01098_ ),
    .X(\u_cpu.REG_FILE._02681_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07378_  (.A1(\u_cpu.REG_FILE._01140_ ),
    .A2(\u_cpu.REG_FILE.rf[29][30] ),
    .B1(\u_cpu.REG_FILE._02681_ ),
    .Y(\u_cpu.REG_FILE._02682_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07379_  (.A1(\u_cpu.REG_FILE._02679_ ),
    .A2(\u_cpu.REG_FILE._02680_ ),
    .B1(\u_cpu.REG_FILE._02682_ ),
    .C1(\u_cpu.REG_FILE._02016_ ),
    .Y(\u_cpu.REG_FILE._02683_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07380_  (.A1(\u_cpu.REG_FILE._02676_ ),
    .A2(\u_cpu.REG_FILE._02678_ ),
    .B1(\u_cpu.REG_FILE._01314_ ),
    .C1(\u_cpu.REG_FILE._02683_ ),
    .Y(\u_cpu.REG_FILE._02684_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07381_  (.A(\u_cpu.REG_FILE.rf[19][30] ),
    .Y(\u_cpu.REG_FILE._02685_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07382_  (.A1(\u_cpu.REG_FILE._01523_ ),
    .A2(\u_cpu.REG_FILE.rf[18][30] ),
    .B1(\u_cpu.REG_FILE._01533_ ),
    .Y(\u_cpu.REG_FILE._02686_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07383_  (.A1(\u_cpu.REG_FILE._02685_ ),
    .A2(\u_cpu.REG_FILE._01399_ ),
    .B1(\u_cpu.REG_FILE._02686_ ),
    .Y(\u_cpu.REG_FILE._02687_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07384_  (.A(\u_cpu.REG_FILE.rf[17][30] ),
    .Y(\u_cpu.REG_FILE._02688_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07385_  (.A1(\u_cpu.REG_FILE._01317_ ),
    .A2(\u_cpu.REG_FILE.rf[16][30] ),
    .B1_N(\u_cpu.REG_FILE._01258_ ),
    .Y(\u_cpu.REG_FILE._02689_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07386_  (.A1(\u_cpu.REG_FILE._02688_ ),
    .A2(\u_cpu.REG_FILE._01399_ ),
    .B1(\u_cpu.REG_FILE._02689_ ),
    .Y(\u_cpu.REG_FILE._02690_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07387_  (.A(\u_cpu.REG_FILE.rf[23][30] ),
    .B_N(\u_cpu.REG_FILE._01408_ ),
    .X(\u_cpu.REG_FILE._02691_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07388_  (.A1(\u_cpu.REG_FILE._01077_ ),
    .A2(\u_cpu.REG_FILE.rf[22][30] ),
    .B1(\u_cpu.REG_FILE._01083_ ),
    .C1(\u_cpu.REG_FILE._02691_ ),
    .Y(\u_cpu.REG_FILE._02692_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07389_  (.A1(\u_cpu.REG_FILE._01324_ ),
    .A2(\u_cpu.REG_FILE.rf[20][30] ),
    .B1_N(\u_cpu.REG_FILE._01304_ ),
    .X(\u_cpu.REG_FILE._02693_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07390_  (.A1(\u_cpu.REG_FILE._01038_ ),
    .A2(\u_cpu.REG_FILE.rf[21][30] ),
    .B1(\u_cpu.REG_FILE._02693_ ),
    .Y(\u_cpu.REG_FILE._02694_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07391_  (.A(\u_cpu.REG_FILE._02692_ ),
    .B(\u_cpu.REG_FILE._02694_ ),
    .C(\u_cpu.REG_FILE._01115_ ),
    .Y(\u_cpu.REG_FILE._02695_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._07392_  (.A1(\u_cpu.REG_FILE._01047_ ),
    .A2(\u_cpu.REG_FILE._02687_ ),
    .A3(\u_cpu.REG_FILE._02690_ ),
    .B1(\u_cpu.REG_FILE._02695_ ),
    .C1(\u_cpu.REG_FILE._01089_ ),
    .Y(\u_cpu.REG_FILE._02696_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07393_  (.A(\u_cpu.REG_FILE._02684_ ),
    .B(\u_cpu.REG_FILE._02696_ ),
    .C(\u_cpu.REG_FILE._01025_ ),
    .Y(\u_cpu.REG_FILE._02697_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07394_  (.A1(\u_cpu.REG_FILE._02662_ ),
    .A2(\u_cpu.REG_FILE._02673_ ),
    .B1(\u_cpu.REG_FILE._02697_ ),
    .C1(\u_cpu.REG_FILE._01164_ ),
    .X(\u_cpu.ALU.SrcA[30] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07395_  (.A(\u_cpu.REG_FILE.rf[15][31] ),
    .B_N(\u_cpu.REG_FILE._01262_ ),
    .X(\u_cpu.REG_FILE._02698_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07396_  (.A1(\u_cpu.REG_FILE._01531_ ),
    .A2(\u_cpu.REG_FILE.rf[14][31] ),
    .B1(\u_cpu.REG_FILE._01288_ ),
    .C1(\u_cpu.REG_FILE._02698_ ),
    .Y(\u_cpu.REG_FILE._02699_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07397_  (.A1(\u_cpu.REG_FILE._01299_ ),
    .A2(\u_cpu.REG_FILE.rf[12][31] ),
    .B1_N(\u_cpu.REG_FILE._01106_ ),
    .X(\u_cpu.REG_FILE._02700_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07398_  (.A1(\u_cpu.REG_FILE._01298_ ),
    .A2(\u_cpu.REG_FILE.rf[13][31] ),
    .B1(\u_cpu.REG_FILE._02700_ ),
    .Y(\u_cpu.REG_FILE._02701_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07399_  (.A(\u_cpu.REG_FILE._02699_ ),
    .B(\u_cpu.REG_FILE._02701_ ),
    .C(\u_cpu.REG_FILE._01293_ ),
    .Y(\u_cpu.REG_FILE._02702_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07400_  (.A_N(\u_cpu.REG_FILE.rf[9][31] ),
    .B(\u_cpu.REG_FILE._01382_ ),
    .X(\u_cpu.REG_FILE._02703_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07401_  (.A1(\u_cpu.REG_FILE._02018_ ),
    .A2(\u_cpu.REG_FILE.rf[8][31] ),
    .B1_N(\u_cpu.REG_FILE._01521_ ),
    .Y(\u_cpu.REG_FILE._02704_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07402_  (.A(\u_cpu.REG_FILE.rf[11][31] ),
    .B_N(\u_cpu.REG_FILE._01345_ ),
    .X(\u_cpu.REG_FILE._02705_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07403_  (.A1(\u_cpu.REG_FILE._01620_ ),
    .A2(\u_cpu.REG_FILE.rf[10][31] ),
    .B1(\u_cpu.REG_FILE._01339_ ),
    .C1(\u_cpu.REG_FILE._02705_ ),
    .Y(\u_cpu.REG_FILE._02706_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07404_  (.A1(\u_cpu.REG_FILE._02703_ ),
    .A2(\u_cpu.REG_FILE._02704_ ),
    .B1(\u_cpu.REG_FILE._01384_ ),
    .C1(\u_cpu.REG_FILE._02706_ ),
    .Y(\u_cpu.REG_FILE._02707_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07405_  (.A(\u_cpu.REG_FILE._02702_ ),
    .B(\u_cpu.REG_FILE._02707_ ),
    .C(\u_cpu.REG_FILE._01117_ ),
    .Y(\u_cpu.REG_FILE._02708_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07406_  (.A(\u_cpu.REG_FILE.rf[5][31] ),
    .Y(\u_cpu.REG_FILE._02709_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07407_  (.A1(\u_cpu.REG_FILE._01133_ ),
    .A2(\u_cpu.REG_FILE.rf[4][31] ),
    .B1_N(\u_cpu.REG_FILE._01380_ ),
    .Y(\u_cpu.REG_FILE._02710_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07408_  (.A1(\u_cpu.REG_FILE._02709_ ),
    .A2(\u_cpu.REG_FILE._01284_ ),
    .B1(\u_cpu.REG_FILE._02710_ ),
    .Y(\u_cpu.REG_FILE._02711_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07409_  (.A1(\u_cpu.REG_FILE._01774_ ),
    .A2(\u_cpu.REG_FILE.rf[6][31] ),
    .B1(\u_cpu.REG_FILE._01400_ ),
    .Y(\u_cpu.REG_FILE._02712_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07410_  (.A_N(\u_cpu.REG_FILE.rf[7][31] ),
    .B(\u_cpu.REG_FILE._01091_ ),
    .X(\u_cpu.REG_FILE._02713_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07411_  (.A1(\u_cpu.REG_FILE._02712_ ),
    .A2(\u_cpu.REG_FILE._02713_ ),
    .B1(\u_cpu.REG_FILE._02122_ ),
    .Y(\u_cpu.REG_FILE._02714_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07412_  (.A_N(\u_cpu.REG_FILE.rf[1][31] ),
    .B(\u_cpu.REG_FILE._01161_ ),
    .X(\u_cpu.REG_FILE._02715_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07413_  (.A1(\u_cpu.REG_FILE._02105_ ),
    .A2(\u_cpu.REG_FILE.rf[0][31] ),
    .B1_N(\u_cpu.REG_FILE._01078_ ),
    .Y(\u_cpu.REG_FILE._02716_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07414_  (.A(\u_cpu.REG_FILE.rf[3][31] ),
    .B_N(\u_cpu.REG_FILE._02057_ ),
    .X(\u_cpu.REG_FILE._02717_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07415_  (.A1(\u_cpu.REG_FILE._01053_ ),
    .A2(\u_cpu.REG_FILE.rf[2][31] ),
    .B1(\u_cpu.REG_FILE._02056_ ),
    .C1(\u_cpu.REG_FILE._02717_ ),
    .Y(\u_cpu.REG_FILE._02718_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07416_  (.A1(\u_cpu.REG_FILE._02715_ ),
    .A2(\u_cpu.REG_FILE._02716_ ),
    .B1(\u_cpu.REG_FILE._01139_ ),
    .C1(\u_cpu.REG_FILE._02718_ ),
    .Y(\u_cpu.REG_FILE._02719_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07417_  (.A1(\u_cpu.REG_FILE._02711_ ),
    .A2(\u_cpu.REG_FILE._02714_ ),
    .B1(\u_cpu.REG_FILE._01414_ ),
    .C1(\u_cpu.REG_FILE._02719_ ),
    .Y(\u_cpu.REG_FILE._02720_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._07418_  (.A(\u_cpu.REG_FILE._02708_ ),
    .B(\u_cpu.REG_FILE._02720_ ),
    .Y(\u_cpu.REG_FILE._02721_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07419_  (.A(\u_cpu.REG_FILE.rf[27][31] ),
    .B_N(\u_cpu.REG_FILE._01528_ ),
    .X(\u_cpu.REG_FILE._02722_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07420_  (.A1(\u_cpu.REG_FILE._01308_ ),
    .A2(\u_cpu.REG_FILE.rf[26][31] ),
    .B1(\u_cpu.REG_FILE._01660_ ),
    .C1(\u_cpu.REG_FILE._02722_ ),
    .X(\u_cpu.REG_FILE._02723_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07421_  (.A1(\u_cpu.REG_FILE._01447_ ),
    .A2(\u_cpu.REG_FILE.rf[24][31] ),
    .B1_N(\u_cpu.REG_FILE._01062_ ),
    .X(\u_cpu.REG_FILE._02724_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07422_  (.A(\u_cpu.REG_FILE.rf[25][31] ),
    .B_N(\u_cpu.REG_FILE._01125_ ),
    .X(\u_cpu.REG_FILE._02725_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._07423_  (.A1(\u_cpu.REG_FILE._02724_ ),
    .A2(\u_cpu.REG_FILE._02725_ ),
    .B1(\u_cpu.REG_FILE._01046_ ),
    .X(\u_cpu.REG_FILE._02726_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07424_  (.A(\u_cpu.REG_FILE._02010_ ),
    .B(\u_cpu.REG_FILE.rf[30][31] ),
    .Y(\u_cpu.REG_FILE._02727_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07425_  (.A1(\u_cpu.REG_FILE.rf[31][31] ),
    .A2(\u_cpu.REG_FILE._01969_ ),
    .B1(\u_cpu.REG_FILE._01107_ ),
    .Y(\u_cpu.REG_FILE._02728_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07426_  (.A1(\u_cpu.REG_FILE._02013_ ),
    .A2(\u_cpu.REG_FILE.rf[28][31] ),
    .B1_N(\u_cpu.REG_FILE._01098_ ),
    .X(\u_cpu.REG_FILE._02729_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07427_  (.A1(\u_cpu.REG_FILE._01140_ ),
    .A2(\u_cpu.REG_FILE.rf[29][31] ),
    .B1(\u_cpu.REG_FILE._02729_ ),
    .Y(\u_cpu.REG_FILE._02730_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07428_  (.A1(\u_cpu.REG_FILE._02727_ ),
    .A2(\u_cpu.REG_FILE._02728_ ),
    .B1(\u_cpu.REG_FILE._02730_ ),
    .C1(\u_cpu.REG_FILE._02016_ ),
    .Y(\u_cpu.REG_FILE._02731_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07429_  (.A1(\u_cpu.REG_FILE._02723_ ),
    .A2(\u_cpu.REG_FILE._02726_ ),
    .B1(\u_cpu.REG_FILE._01314_ ),
    .C1(\u_cpu.REG_FILE._02731_ ),
    .Y(\u_cpu.REG_FILE._02732_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07430_  (.A1(\u_cpu.REG_FILE._01260_ ),
    .A2(\u_cpu.REG_FILE.rf[18][31] ),
    .B1(\u_cpu.REG_FILE._01407_ ),
    .Y(\u_cpu.REG_FILE._02733_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07431_  (.A(\u_cpu.REG_FILE.rf[19][31] ),
    .B(\u_cpu.REG_FILE._01509_ ),
    .Y(\u_cpu.REG_FILE._02734_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07432_  (.A1(\u_cpu.REG_FILE._01152_ ),
    .A2(\u_cpu.REG_FILE.rf[16][31] ),
    .B1_N(\u_cpu.REG_FILE._01153_ ),
    .X(\u_cpu.REG_FILE._02735_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07433_  (.A1(\u_cpu.REG_FILE._01726_ ),
    .A2(\u_cpu.REG_FILE.rf[17][31] ),
    .B1(\u_cpu.REG_FILE._02735_ ),
    .Y(\u_cpu.REG_FILE._02736_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07434_  (.A1(\u_cpu.REG_FILE._02733_ ),
    .A2(\u_cpu.REG_FILE._02734_ ),
    .B1(\u_cpu.REG_FILE._01264_ ),
    .C1(\u_cpu.REG_FILE._02736_ ),
    .Y(\u_cpu.REG_FILE._02737_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._07435_  (.A(\u_cpu.REG_FILE._01324_ ),
    .B(\u_cpu.REG_FILE.rf[22][31] ),
    .X(\u_cpu.REG_FILE._02738_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07436_  (.A1(\u_cpu.REG_FILE._01321_ ),
    .A2(\u_cpu.REG_FILE.rf[23][31] ),
    .B1(\u_cpu.REG_FILE._01063_ ),
    .C1(\u_cpu.REG_FILE._02738_ ),
    .Y(\u_cpu.REG_FILE._02739_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07437_  (.A1(\u_cpu.REG_FILE._01632_ ),
    .A2(\u_cpu.REG_FILE.rf[20][31] ),
    .B1_N(\u_cpu.REG_FILE._01134_ ),
    .X(\u_cpu.REG_FILE._02740_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07438_  (.A1(\u_cpu.REG_FILE._01120_ ),
    .A2(\u_cpu.REG_FILE.rf[21][31] ),
    .B1(\u_cpu.REG_FILE._02740_ ),
    .Y(\u_cpu.REG_FILE._02741_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07439_  (.A(\u_cpu.REG_FILE._02739_ ),
    .B(\u_cpu.REG_FILE._02741_ ),
    .C(\u_cpu.REG_FILE._01552_ ),
    .Y(\u_cpu.REG_FILE._02742_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07440_  (.A(\u_cpu.REG_FILE._01541_ ),
    .B(\u_cpu.REG_FILE._02737_ ),
    .C(\u_cpu.REG_FILE._02742_ ),
    .Y(\u_cpu.REG_FILE._02743_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07441_  (.A(\u_cpu.REG_FILE._02732_ ),
    .B(\u_cpu.REG_FILE._02743_ ),
    .C(\u_cpu.REG_FILE._01025_ ),
    .Y(\u_cpu.REG_FILE._02744_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07442_  (.A1(\u_cpu.REG_FILE._01159_ ),
    .A2(\u_cpu.REG_FILE._02721_ ),
    .B1(\u_cpu.REG_FILE._02744_ ),
    .C1(\u_cpu.REG_FILE._01164_ ),
    .X(\u_cpu.ALU.SrcA[31] ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07443_  (.A(\u_cpu.M_AXI_WDATA[24] ),
    .X(\u_cpu.REG_FILE._02745_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07444_  (.A(\u_cpu.REG_FILE._02745_ ),
    .X(\u_cpu.REG_FILE._02746_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07445_  (.A(\u_cpu.M_AXI_WDATA[20] ),
    .X(\u_cpu.REG_FILE._02747_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07446_  (.A(\u_cpu.REG_FILE._02747_ ),
    .X(\u_cpu.REG_FILE._02748_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07447_  (.A(\u_cpu.REG_FILE._02748_ ),
    .X(\u_cpu.REG_FILE._02749_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07448_  (.A(\u_cpu.M_AXI_WDATA[21] ),
    .X(\u_cpu.REG_FILE._02750_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07449_  (.A(\u_cpu.REG_FILE._02750_ ),
    .X(\u_cpu.REG_FILE._02751_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07450_  (.A(\u_cpu.REG_FILE._02751_ ),
    .X(\u_cpu.REG_FILE._02752_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07451_  (.A(\u_cpu.M_AXI_WDATA[20] ),
    .X(\u_cpu.REG_FILE._02753_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07452_  (.A(\u_cpu.REG_FILE._02753_ ),
    .X(\u_cpu.REG_FILE._02754_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07453_  (.A(\u_cpu.REG_FILE.rf[15][0] ),
    .B_N(\u_cpu.REG_FILE._02754_ ),
    .X(\u_cpu.REG_FILE._02755_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07454_  (.A1(\u_cpu.REG_FILE.rf[14][0] ),
    .A2(\u_cpu.REG_FILE._02749_ ),
    .B1(\u_cpu.REG_FILE._02752_ ),
    .C1(\u_cpu.REG_FILE._02755_ ),
    .Y(\u_cpu.REG_FILE._02756_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07455_  (.A(\u_cpu.M_AXI_WDATA[20] ),
    .Y(\u_cpu.REG_FILE._02757_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07456_  (.A(\u_cpu.REG_FILE._02757_ ),
    .X(\u_cpu.REG_FILE._02758_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07457_  (.A(\u_cpu.REG_FILE._02758_ ),
    .X(\u_cpu.REG_FILE._02759_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07458_  (.A(\u_cpu.REG_FILE._02753_ ),
    .X(\u_cpu.REG_FILE._02760_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07459_  (.A(\u_cpu.REG_FILE._02750_ ),
    .X(\u_cpu.REG_FILE._02761_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07460_  (.A1(\u_cpu.REG_FILE.rf[12][0] ),
    .A2(\u_cpu.REG_FILE._02760_ ),
    .B1_N(\u_cpu.REG_FILE._02761_ ),
    .X(\u_cpu.REG_FILE._02762_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07461_  (.A1(\u_cpu.REG_FILE.rf[13][0] ),
    .A2(\u_cpu.REG_FILE._02759_ ),
    .B1(\u_cpu.REG_FILE._02762_ ),
    .Y(\u_cpu.REG_FILE._02763_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07462_  (.A(\u_cpu.M_AXI_WDATA[22] ),
    .X(\u_cpu.REG_FILE._02764_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07463_  (.A(\u_cpu.REG_FILE._02764_ ),
    .X(\u_cpu.REG_FILE._02765_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07464_  (.A(\u_cpu.REG_FILE._02756_ ),
    .B(\u_cpu.REG_FILE._02763_ ),
    .C(\u_cpu.REG_FILE._02765_ ),
    .Y(\u_cpu.REG_FILE._02766_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07465_  (.A(\u_cpu.M_AXI_WDATA[20] ),
    .X(\u_cpu.REG_FILE._02767_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07466_  (.A(\u_cpu.REG_FILE._02767_ ),
    .X(\u_cpu.REG_FILE._02768_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07467_  (.A_N(\u_cpu.REG_FILE.rf[9][0] ),
    .B(\u_cpu.REG_FILE._02768_ ),
    .X(\u_cpu.REG_FILE._02769_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07468_  (.A(\u_cpu.M_AXI_WDATA[20] ),
    .X(\u_cpu.REG_FILE._02770_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07469_  (.A(\u_cpu.REG_FILE._02770_ ),
    .X(\u_cpu.REG_FILE._02771_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07470_  (.A(\u_cpu.REG_FILE._02771_ ),
    .X(\u_cpu.REG_FILE._02772_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07471_  (.A(\u_cpu.M_AXI_WDATA[21] ),
    .X(\u_cpu.REG_FILE._02773_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07472_  (.A(\u_cpu.REG_FILE._02773_ ),
    .X(\u_cpu.REG_FILE._02774_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07473_  (.A1(\u_cpu.REG_FILE.rf[8][0] ),
    .A2(\u_cpu.REG_FILE._02772_ ),
    .B1_N(\u_cpu.REG_FILE._02774_ ),
    .Y(\u_cpu.REG_FILE._02775_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07474_  (.A(\u_cpu.M_AXI_WDATA[22] ),
    .Y(\u_cpu.REG_FILE._02776_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07475_  (.A(\u_cpu.REG_FILE._02776_ ),
    .X(\u_cpu.REG_FILE._02777_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07476_  (.A(\u_cpu.M_AXI_WDATA[20] ),
    .X(\u_cpu.REG_FILE._02778_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07477_  (.A(\u_cpu.REG_FILE._02778_ ),
    .X(\u_cpu.REG_FILE._02779_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07478_  (.A(\u_cpu.REG_FILE._02779_ ),
    .X(\u_cpu.REG_FILE._02780_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07479_  (.A(\u_cpu.REG_FILE._02750_ ),
    .X(\u_cpu.REG_FILE._02781_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07480_  (.A(\u_cpu.REG_FILE._02781_ ),
    .X(\u_cpu.REG_FILE._02782_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07481_  (.A(\u_cpu.REG_FILE._02778_ ),
    .X(\u_cpu.REG_FILE._02783_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07482_  (.A(\u_cpu.REG_FILE.rf[11][0] ),
    .B_N(\u_cpu.REG_FILE._02783_ ),
    .X(\u_cpu.REG_FILE._02784_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07483_  (.A1(\u_cpu.REG_FILE.rf[10][0] ),
    .A2(\u_cpu.REG_FILE._02780_ ),
    .B1(\u_cpu.REG_FILE._02782_ ),
    .C1(\u_cpu.REG_FILE._02784_ ),
    .Y(\u_cpu.REG_FILE._02785_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07484_  (.A1(\u_cpu.REG_FILE._02769_ ),
    .A2(\u_cpu.REG_FILE._02775_ ),
    .B1(\u_cpu.REG_FILE._02777_ ),
    .C1(\u_cpu.REG_FILE._02785_ ),
    .Y(\u_cpu.REG_FILE._02786_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07485_  (.A(\u_cpu.M_AXI_WDATA[23] ),
    .X(\u_cpu.REG_FILE._02787_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07486_  (.A(\u_cpu.REG_FILE._02787_ ),
    .X(\u_cpu.REG_FILE._02788_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07487_  (.A(\u_cpu.REG_FILE._02766_ ),
    .B(\u_cpu.REG_FILE._02786_ ),
    .C(\u_cpu.REG_FILE._02788_ ),
    .Y(\u_cpu.REG_FILE._02789_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07488_  (.A(\u_cpu.REG_FILE._02747_ ),
    .X(\u_cpu.REG_FILE._02790_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07489_  (.A(\u_cpu.REG_FILE._02790_ ),
    .X(\u_cpu.REG_FILE._02791_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07490_  (.A(\u_cpu.REG_FILE._02770_ ),
    .X(\u_cpu.REG_FILE._02792_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07491_  (.A(\u_cpu.REG_FILE._02792_ ),
    .X(\u_cpu.REG_FILE._02793_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07492_  (.A(\u_cpu.REG_FILE._02773_ ),
    .X(\u_cpu.REG_FILE._02794_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07493_  (.A1(\u_cpu.REG_FILE.rf[4][0] ),
    .A2(\u_cpu.REG_FILE._02793_ ),
    .B1_N(\u_cpu.REG_FILE._02794_ ),
    .Y(\u_cpu.REG_FILE._02795_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07494_  (.A1(\u_cpu.REG_FILE._01072_ ),
    .A2(\u_cpu.REG_FILE._02791_ ),
    .B1(\u_cpu.REG_FILE._02795_ ),
    .Y(\u_cpu.REG_FILE._02796_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07495_  (.A(\u_cpu.REG_FILE._02767_ ),
    .X(\u_cpu.REG_FILE._02797_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07496_  (.A(\u_cpu.M_AXI_WDATA[21] ),
    .X(\u_cpu.REG_FILE._02798_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07497_  (.A(\u_cpu.REG_FILE._02798_ ),
    .X(\u_cpu.REG_FILE._02799_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07498_  (.A1(\u_cpu.REG_FILE.rf[6][0] ),
    .A2(\u_cpu.REG_FILE._02797_ ),
    .B1(\u_cpu.REG_FILE._02799_ ),
    .Y(\u_cpu.REG_FILE._02800_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07499_  (.A(\u_cpu.REG_FILE._02747_ ),
    .X(\u_cpu.REG_FILE._02801_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07500_  (.A_N(\u_cpu.REG_FILE.rf[7][0] ),
    .B(\u_cpu.REG_FILE._02801_ ),
    .X(\u_cpu.REG_FILE._02802_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07501_  (.A(\u_cpu.M_AXI_WDATA[22] ),
    .X(\u_cpu.REG_FILE._02803_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07502_  (.A(\u_cpu.REG_FILE._02803_ ),
    .X(\u_cpu.REG_FILE._02804_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07503_  (.A1(\u_cpu.REG_FILE._02800_ ),
    .A2(\u_cpu.REG_FILE._02802_ ),
    .B1(\u_cpu.REG_FILE._02804_ ),
    .Y(\u_cpu.REG_FILE._02805_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07504_  (.A(\u_cpu.REG_FILE._02787_ ),
    .Y(\u_cpu.REG_FILE._02806_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07505_  (.A(\u_cpu.REG_FILE._02806_ ),
    .X(\u_cpu.REG_FILE._02807_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07506_  (.A(\u_cpu.REG_FILE._02747_ ),
    .X(\u_cpu.REG_FILE._02808_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07507_  (.A_N(\u_cpu.REG_FILE.rf[1][0] ),
    .B(\u_cpu.REG_FILE._02808_ ),
    .X(\u_cpu.REG_FILE._02809_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07508_  (.A(\u_cpu.REG_FILE._02770_ ),
    .X(\u_cpu.REG_FILE._02810_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07509_  (.A(\u_cpu.REG_FILE._02810_ ),
    .X(\u_cpu.REG_FILE._02811_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07510_  (.A(\u_cpu.REG_FILE._02750_ ),
    .X(\u_cpu.REG_FILE._02812_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07511_  (.A1(\u_cpu.REG_FILE.rf[0][0] ),
    .A2(\u_cpu.REG_FILE._02811_ ),
    .B1_N(\u_cpu.REG_FILE._02812_ ),
    .Y(\u_cpu.REG_FILE._02813_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07512_  (.A(\u_cpu.REG_FILE._02776_ ),
    .X(\u_cpu.REG_FILE._02814_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07513_  (.A(\u_cpu.REG_FILE._02778_ ),
    .X(\u_cpu.REG_FILE._02815_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07514_  (.A(\u_cpu.REG_FILE._02815_ ),
    .X(\u_cpu.REG_FILE._02816_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07515_  (.A(\u_cpu.REG_FILE._02750_ ),
    .X(\u_cpu.REG_FILE._02817_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07516_  (.A(\u_cpu.REG_FILE._02817_ ),
    .X(\u_cpu.REG_FILE._02818_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07517_  (.A(\u_cpu.REG_FILE.rf[3][0] ),
    .B_N(\u_cpu.REG_FILE._02771_ ),
    .X(\u_cpu.REG_FILE._02819_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07518_  (.A1(\u_cpu.REG_FILE.rf[2][0] ),
    .A2(\u_cpu.REG_FILE._02816_ ),
    .B1(\u_cpu.REG_FILE._02818_ ),
    .C1(\u_cpu.REG_FILE._02819_ ),
    .Y(\u_cpu.REG_FILE._02820_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07519_  (.A1(\u_cpu.REG_FILE._02809_ ),
    .A2(\u_cpu.REG_FILE._02813_ ),
    .B1(\u_cpu.REG_FILE._02814_ ),
    .C1(\u_cpu.REG_FILE._02820_ ),
    .Y(\u_cpu.REG_FILE._02821_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07520_  (.A1(\u_cpu.REG_FILE._02796_ ),
    .A2(\u_cpu.REG_FILE._02805_ ),
    .B1(\u_cpu.REG_FILE._02807_ ),
    .C1(\u_cpu.REG_FILE._02821_ ),
    .Y(\u_cpu.REG_FILE._02822_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._07521_  (.A(\u_cpu.REG_FILE._02789_ ),
    .B(\u_cpu.REG_FILE._02822_ ),
    .Y(\u_cpu.REG_FILE._02823_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07522_  (.A(\u_cpu.REG_FILE._02783_ ),
    .X(\u_cpu.REG_FILE._02824_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07523_  (.A(\u_cpu.REG_FILE._02750_ ),
    .X(\u_cpu.REG_FILE._02825_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07524_  (.A(\u_cpu.REG_FILE._02825_ ),
    .X(\u_cpu.REG_FILE._02826_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07525_  (.A(\u_cpu.REG_FILE._02753_ ),
    .X(\u_cpu.REG_FILE._02827_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07526_  (.A(\u_cpu.REG_FILE.rf[27][0] ),
    .B_N(\u_cpu.REG_FILE._02827_ ),
    .X(\u_cpu.REG_FILE._02828_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07527_  (.A1(\u_cpu.REG_FILE.rf[26][0] ),
    .A2(\u_cpu.REG_FILE._02824_ ),
    .B1(\u_cpu.REG_FILE._02826_ ),
    .C1(\u_cpu.REG_FILE._02828_ ),
    .X(\u_cpu.REG_FILE._02829_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07528_  (.A(\u_cpu.REG_FILE._02747_ ),
    .X(\u_cpu.REG_FILE._02830_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07529_  (.A1(\u_cpu.REG_FILE.rf[24][0] ),
    .A2(\u_cpu.REG_FILE._02830_ ),
    .B1_N(\u_cpu.REG_FILE._02825_ ),
    .X(\u_cpu.REG_FILE._02831_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07530_  (.A(\u_cpu.REG_FILE._02778_ ),
    .X(\u_cpu.REG_FILE._02832_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07531_  (.A(\u_cpu.REG_FILE.rf[25][0] ),
    .B_N(\u_cpu.REG_FILE._02832_ ),
    .X(\u_cpu.REG_FILE._02833_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07532_  (.A(\u_cpu.M_AXI_WDATA[22] ),
    .X(\u_cpu.REG_FILE._02834_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._07533_  (.A1(\u_cpu.REG_FILE._02831_ ),
    .A2(\u_cpu.REG_FILE._02833_ ),
    .B1(\u_cpu.REG_FILE._02834_ ),
    .X(\u_cpu.REG_FILE._02835_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07534_  (.A(\u_cpu.REG_FILE._02787_ ),
    .X(\u_cpu.REG_FILE._02836_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07535_  (.A(\u_cpu.REG_FILE._02767_ ),
    .X(\u_cpu.REG_FILE._02837_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07536_  (.A(\u_cpu.REG_FILE._02773_ ),
    .X(\u_cpu.REG_FILE._02838_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07537_  (.A1(\u_cpu.REG_FILE.rf[28][0] ),
    .A2(\u_cpu.REG_FILE._02837_ ),
    .B1_N(\u_cpu.REG_FILE._02838_ ),
    .Y(\u_cpu.REG_FILE._02839_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07538_  (.A(\u_cpu.REG_FILE._02757_ ),
    .X(\u_cpu.REG_FILE._02840_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07539_  (.A(\u_cpu.REG_FILE._02840_ ),
    .X(\u_cpu.REG_FILE._02841_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07540_  (.A(\u_cpu.REG_FILE.rf[29][0] ),
    .B(\u_cpu.REG_FILE._02841_ ),
    .Y(\u_cpu.REG_FILE._02842_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07541_  (.A(\u_cpu.REG_FILE._02779_ ),
    .X(\u_cpu.REG_FILE._02843_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07542_  (.A(\u_cpu.REG_FILE.rf[30][0] ),
    .B(\u_cpu.REG_FILE._02843_ ),
    .Y(\u_cpu.REG_FILE._02844_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07543_  (.A(\u_cpu.REG_FILE._02840_ ),
    .X(\u_cpu.REG_FILE._02845_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07544_  (.A(\u_cpu.REG_FILE._02781_ ),
    .X(\u_cpu.REG_FILE._02846_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07545_  (.A1(\u_cpu.REG_FILE.rf[31][0] ),
    .A2(\u_cpu.REG_FILE._02845_ ),
    .B1(\u_cpu.REG_FILE._02846_ ),
    .Y(\u_cpu.REG_FILE._02847_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07546_  (.A(\u_cpu.REG_FILE._02803_ ),
    .X(\u_cpu.REG_FILE._02848_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._07547_  (.A1(\u_cpu.REG_FILE._02839_ ),
    .A2(\u_cpu.REG_FILE._02842_ ),
    .B1(\u_cpu.REG_FILE._02844_ ),
    .B2(\u_cpu.REG_FILE._02847_ ),
    .C1(\u_cpu.REG_FILE._02848_ ),
    .Y(\u_cpu.REG_FILE._02849_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07548_  (.A1(\u_cpu.REG_FILE._02829_ ),
    .A2(\u_cpu.REG_FILE._02835_ ),
    .B1(\u_cpu.REG_FILE._02836_ ),
    .C1(\u_cpu.REG_FILE._02849_ ),
    .Y(\u_cpu.REG_FILE._02850_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07549_  (.A(\u_cpu.REG_FILE._02806_ ),
    .X(\u_cpu.REG_FILE._02851_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07550_  (.A(\u_cpu.REG_FILE._02770_ ),
    .X(\u_cpu.REG_FILE._02852_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07551_  (.A(\u_cpu.REG_FILE._02852_ ),
    .X(\u_cpu.REG_FILE._02853_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07552_  (.A(\u_cpu.REG_FILE._02798_ ),
    .X(\u_cpu.REG_FILE._02854_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07553_  (.A1(\u_cpu.REG_FILE.rf[18][0] ),
    .A2(\u_cpu.REG_FILE._02853_ ),
    .B1(\u_cpu.REG_FILE._02854_ ),
    .Y(\u_cpu.REG_FILE._02855_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07554_  (.A(\u_cpu.REG_FILE._02758_ ),
    .X(\u_cpu.REG_FILE._02856_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07555_  (.A(\u_cpu.REG_FILE.rf[19][0] ),
    .B(\u_cpu.REG_FILE._02856_ ),
    .Y(\u_cpu.REG_FILE._02857_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07556_  (.A(\u_cpu.REG_FILE._02776_ ),
    .X(\u_cpu.REG_FILE._02858_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07557_  (.A(\u_cpu.REG_FILE._02758_ ),
    .X(\u_cpu.REG_FILE._02859_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07558_  (.A(\u_cpu.REG_FILE._02753_ ),
    .X(\u_cpu.REG_FILE._02860_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07559_  (.A(\u_cpu.M_AXI_WDATA[21] ),
    .X(\u_cpu.REG_FILE._02861_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07560_  (.A1(\u_cpu.REG_FILE.rf[16][0] ),
    .A2(\u_cpu.REG_FILE._02860_ ),
    .B1_N(\u_cpu.REG_FILE._02861_ ),
    .X(\u_cpu.REG_FILE._02862_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07561_  (.A1(\u_cpu.REG_FILE.rf[17][0] ),
    .A2(\u_cpu.REG_FILE._02859_ ),
    .B1(\u_cpu.REG_FILE._02862_ ),
    .Y(\u_cpu.REG_FILE._02863_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07562_  (.A1(\u_cpu.REG_FILE._02855_ ),
    .A2(\u_cpu.REG_FILE._02857_ ),
    .B1(\u_cpu.REG_FILE._02858_ ),
    .C1(\u_cpu.REG_FILE._02863_ ),
    .Y(\u_cpu.REG_FILE._02864_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07563_  (.A(\u_cpu.REG_FILE._02750_ ),
    .X(\u_cpu.REG_FILE._02865_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07564_  (.A(\u_cpu.REG_FILE._02865_ ),
    .X(\u_cpu.REG_FILE._02866_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07565_  (.A(\u_cpu.REG_FILE._02770_ ),
    .X(\u_cpu.REG_FILE._02867_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._07566_  (.A(\u_cpu.REG_FILE.rf[22][0] ),
    .B(\u_cpu.REG_FILE._02867_ ),
    .X(\u_cpu.REG_FILE._02868_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07567_  (.A1(\u_cpu.REG_FILE.rf[23][0] ),
    .A2(\u_cpu.REG_FILE._02841_ ),
    .B1(\u_cpu.REG_FILE._02866_ ),
    .C1(\u_cpu.REG_FILE._02868_ ),
    .Y(\u_cpu.REG_FILE._02869_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07568_  (.A(\u_cpu.REG_FILE._02840_ ),
    .X(\u_cpu.REG_FILE._02870_ ));
 sky130_fd_sc_hd__buf_2 \u_cpu.REG_FILE._07569_  (.A(\u_cpu.REG_FILE._02770_ ),
    .X(\u_cpu.REG_FILE._02871_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07570_  (.A(\u_cpu.M_AXI_WDATA[21] ),
    .X(\u_cpu.REG_FILE._02872_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07571_  (.A1(\u_cpu.REG_FILE.rf[20][0] ),
    .A2(\u_cpu.REG_FILE._02871_ ),
    .B1_N(\u_cpu.REG_FILE._02872_ ),
    .X(\u_cpu.REG_FILE._02873_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07572_  (.A1(\u_cpu.REG_FILE.rf[21][0] ),
    .A2(\u_cpu.REG_FILE._02870_ ),
    .B1(\u_cpu.REG_FILE._02873_ ),
    .Y(\u_cpu.REG_FILE._02874_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07573_  (.A(\u_cpu.REG_FILE._02803_ ),
    .X(\u_cpu.REG_FILE._02875_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07574_  (.A(\u_cpu.REG_FILE._02869_ ),
    .B(\u_cpu.REG_FILE._02874_ ),
    .C(\u_cpu.REG_FILE._02875_ ),
    .Y(\u_cpu.REG_FILE._02876_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07575_  (.A(\u_cpu.REG_FILE._02851_ ),
    .B(\u_cpu.REG_FILE._02864_ ),
    .C(\u_cpu.REG_FILE._02876_ ),
    .Y(\u_cpu.REG_FILE._02877_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07576_  (.A(\u_cpu.REG_FILE._02745_ ),
    .X(\u_cpu.REG_FILE._02878_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07577_  (.A(\u_cpu.REG_FILE._02850_ ),
    .B(\u_cpu.REG_FILE._02877_ ),
    .C(\u_cpu.REG_FILE._02878_ ),
    .Y(\u_cpu.REG_FILE._02879_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07578_  (.A(\u_cpu.REG_FILE._02747_ ),
    .X(\u_cpu.REG_FILE._02880_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.REG_FILE._07579_  (.A(\u_cpu.M_AXI_WDATA[21] ),
    .B(\u_cpu.M_AXI_WDATA[22] ),
    .C(\u_cpu.REG_FILE._02787_ ),
    .X(\u_cpu.REG_FILE._02881_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu.REG_FILE._07580_  (.A(\u_cpu.REG_FILE._02745_ ),
    .B(\u_cpu.REG_FILE._02880_ ),
    .C(\u_cpu.REG_FILE._02881_ ),
    .X(\u_cpu.REG_FILE._02882_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07581_  (.A(\u_cpu.REG_FILE._02882_ ),
    .X(\u_cpu.REG_FILE._02883_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07582_  (.A(\u_cpu.REG_FILE._02883_ ),
    .X(\u_cpu.REG_FILE._02884_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07583_  (.A1(\u_cpu.REG_FILE._02746_ ),
    .A2(\u_cpu.REG_FILE._02823_ ),
    .B1(\u_cpu.REG_FILE._02879_ ),
    .C1(\u_cpu.REG_FILE._02884_ ),
    .X(\u_cpu.ALU.SrcB[0] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07584_  (.A(\u_cpu.REG_FILE.rf[15][1] ),
    .B_N(\u_cpu.REG_FILE._02754_ ),
    .X(\u_cpu.REG_FILE._02885_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07585_  (.A1(\u_cpu.REG_FILE.rf[14][1] ),
    .A2(\u_cpu.REG_FILE._02749_ ),
    .B1(\u_cpu.REG_FILE._02752_ ),
    .C1(\u_cpu.REG_FILE._02885_ ),
    .Y(\u_cpu.REG_FILE._02886_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07586_  (.A1(\u_cpu.REG_FILE.rf[12][1] ),
    .A2(\u_cpu.REG_FILE._02760_ ),
    .B1_N(\u_cpu.REG_FILE._02761_ ),
    .X(\u_cpu.REG_FILE._02887_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07587_  (.A1(\u_cpu.REG_FILE.rf[13][1] ),
    .A2(\u_cpu.REG_FILE._02759_ ),
    .B1(\u_cpu.REG_FILE._02887_ ),
    .Y(\u_cpu.REG_FILE._02888_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07588_  (.A(\u_cpu.REG_FILE._02886_ ),
    .B(\u_cpu.REG_FILE._02888_ ),
    .C(\u_cpu.REG_FILE._02765_ ),
    .Y(\u_cpu.REG_FILE._02889_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07589_  (.A_N(\u_cpu.REG_FILE.rf[9][1] ),
    .B(\u_cpu.REG_FILE._02768_ ),
    .X(\u_cpu.REG_FILE._02890_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07590_  (.A1(\u_cpu.REG_FILE.rf[8][1] ),
    .A2(\u_cpu.REG_FILE._02772_ ),
    .B1_N(\u_cpu.REG_FILE._02774_ ),
    .Y(\u_cpu.REG_FILE._02891_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07591_  (.A(\u_cpu.REG_FILE.rf[11][1] ),
    .B_N(\u_cpu.REG_FILE._02783_ ),
    .X(\u_cpu.REG_FILE._02892_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07592_  (.A1(\u_cpu.REG_FILE.rf[10][1] ),
    .A2(\u_cpu.REG_FILE._02780_ ),
    .B1(\u_cpu.REG_FILE._02782_ ),
    .C1(\u_cpu.REG_FILE._02892_ ),
    .Y(\u_cpu.REG_FILE._02893_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07593_  (.A1(\u_cpu.REG_FILE._02890_ ),
    .A2(\u_cpu.REG_FILE._02891_ ),
    .B1(\u_cpu.REG_FILE._02777_ ),
    .C1(\u_cpu.REG_FILE._02893_ ),
    .Y(\u_cpu.REG_FILE._02894_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07594_  (.A(\u_cpu.REG_FILE._02889_ ),
    .B(\u_cpu.REG_FILE._02894_ ),
    .C(\u_cpu.REG_FILE._02788_ ),
    .Y(\u_cpu.REG_FILE._02895_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07595_  (.A1(\u_cpu.REG_FILE.rf[4][1] ),
    .A2(\u_cpu.REG_FILE._02793_ ),
    .B1_N(\u_cpu.REG_FILE._02794_ ),
    .Y(\u_cpu.REG_FILE._02896_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07596_  (.A1(\u_cpu.REG_FILE._01177_ ),
    .A2(\u_cpu.REG_FILE._02791_ ),
    .B1(\u_cpu.REG_FILE._02896_ ),
    .Y(\u_cpu.REG_FILE._02897_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07597_  (.A1(\u_cpu.REG_FILE.rf[6][1] ),
    .A2(\u_cpu.REG_FILE._02797_ ),
    .B1(\u_cpu.REG_FILE._02799_ ),
    .Y(\u_cpu.REG_FILE._02898_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07598_  (.A_N(\u_cpu.REG_FILE.rf[7][1] ),
    .B(\u_cpu.REG_FILE._02801_ ),
    .X(\u_cpu.REG_FILE._02899_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07599_  (.A1(\u_cpu.REG_FILE._02898_ ),
    .A2(\u_cpu.REG_FILE._02899_ ),
    .B1(\u_cpu.REG_FILE._02804_ ),
    .Y(\u_cpu.REG_FILE._02900_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07600_  (.A_N(\u_cpu.REG_FILE.rf[1][1] ),
    .B(\u_cpu.REG_FILE._02808_ ),
    .X(\u_cpu.REG_FILE._02901_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07601_  (.A1(\u_cpu.REG_FILE.rf[0][1] ),
    .A2(\u_cpu.REG_FILE._02811_ ),
    .B1_N(\u_cpu.REG_FILE._02812_ ),
    .Y(\u_cpu.REG_FILE._02902_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07602_  (.A(\u_cpu.REG_FILE._02815_ ),
    .X(\u_cpu.REG_FILE._02903_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07603_  (.A(\u_cpu.REG_FILE.rf[3][1] ),
    .B_N(\u_cpu.REG_FILE._02771_ ),
    .X(\u_cpu.REG_FILE._02904_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07604_  (.A1(\u_cpu.REG_FILE.rf[2][1] ),
    .A2(\u_cpu.REG_FILE._02903_ ),
    .B1(\u_cpu.REG_FILE._02818_ ),
    .C1(\u_cpu.REG_FILE._02904_ ),
    .Y(\u_cpu.REG_FILE._02905_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07605_  (.A1(\u_cpu.REG_FILE._02901_ ),
    .A2(\u_cpu.REG_FILE._02902_ ),
    .B1(\u_cpu.REG_FILE._02814_ ),
    .C1(\u_cpu.REG_FILE._02905_ ),
    .Y(\u_cpu.REG_FILE._02906_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07606_  (.A1(\u_cpu.REG_FILE._02897_ ),
    .A2(\u_cpu.REG_FILE._02900_ ),
    .B1(\u_cpu.REG_FILE._02807_ ),
    .C1(\u_cpu.REG_FILE._02906_ ),
    .Y(\u_cpu.REG_FILE._02907_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._07607_  (.A(\u_cpu.REG_FILE._02895_ ),
    .B(\u_cpu.REG_FILE._02907_ ),
    .Y(\u_cpu.REG_FILE._02908_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07608_  (.A(\u_cpu.REG_FILE.rf[27][1] ),
    .B_N(\u_cpu.REG_FILE._02827_ ),
    .X(\u_cpu.REG_FILE._02909_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07609_  (.A1(\u_cpu.REG_FILE.rf[26][1] ),
    .A2(\u_cpu.REG_FILE._02824_ ),
    .B1(\u_cpu.REG_FILE._02826_ ),
    .C1(\u_cpu.REG_FILE._02909_ ),
    .X(\u_cpu.REG_FILE._02910_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07610_  (.A1(\u_cpu.REG_FILE.rf[24][1] ),
    .A2(\u_cpu.REG_FILE._02830_ ),
    .B1_N(\u_cpu.REG_FILE._02825_ ),
    .X(\u_cpu.REG_FILE._02911_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07611_  (.A(\u_cpu.REG_FILE.rf[25][1] ),
    .B_N(\u_cpu.REG_FILE._02832_ ),
    .X(\u_cpu.REG_FILE._02912_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._07612_  (.A1(\u_cpu.REG_FILE._02911_ ),
    .A2(\u_cpu.REG_FILE._02912_ ),
    .B1(\u_cpu.REG_FILE._02834_ ),
    .X(\u_cpu.REG_FILE._02913_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07613_  (.A1(\u_cpu.REG_FILE.rf[28][1] ),
    .A2(\u_cpu.REG_FILE._02837_ ),
    .B1_N(\u_cpu.REG_FILE._02838_ ),
    .Y(\u_cpu.REG_FILE._02914_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07614_  (.A(\u_cpu.REG_FILE.rf[29][1] ),
    .B(\u_cpu.REG_FILE._02841_ ),
    .Y(\u_cpu.REG_FILE._02915_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07615_  (.A(\u_cpu.REG_FILE._02779_ ),
    .X(\u_cpu.REG_FILE._02916_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07616_  (.A(\u_cpu.REG_FILE.rf[30][1] ),
    .B(\u_cpu.REG_FILE._02916_ ),
    .Y(\u_cpu.REG_FILE._02917_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07617_  (.A1(\u_cpu.REG_FILE.rf[31][1] ),
    .A2(\u_cpu.REG_FILE._02845_ ),
    .B1(\u_cpu.REG_FILE._02846_ ),
    .Y(\u_cpu.REG_FILE._02918_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07618_  (.A(\u_cpu.REG_FILE._02803_ ),
    .X(\u_cpu.REG_FILE._02919_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._07619_  (.A1(\u_cpu.REG_FILE._02914_ ),
    .A2(\u_cpu.REG_FILE._02915_ ),
    .B1(\u_cpu.REG_FILE._02917_ ),
    .B2(\u_cpu.REG_FILE._02918_ ),
    .C1(\u_cpu.REG_FILE._02919_ ),
    .Y(\u_cpu.REG_FILE._02920_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07620_  (.A1(\u_cpu.REG_FILE._02910_ ),
    .A2(\u_cpu.REG_FILE._02913_ ),
    .B1(\u_cpu.REG_FILE._02836_ ),
    .C1(\u_cpu.REG_FILE._02920_ ),
    .Y(\u_cpu.REG_FILE._02921_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07621_  (.A(\u_cpu.REG_FILE._02806_ ),
    .X(\u_cpu.REG_FILE._02922_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07622_  (.A(\u_cpu.REG_FILE._02792_ ),
    .X(\u_cpu.REG_FILE._02923_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07623_  (.A1(\u_cpu.REG_FILE.rf[18][1] ),
    .A2(\u_cpu.REG_FILE._02923_ ),
    .B1(\u_cpu.REG_FILE._02854_ ),
    .Y(\u_cpu.REG_FILE._02924_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07624_  (.A(\u_cpu.REG_FILE.rf[19][1] ),
    .B(\u_cpu.REG_FILE._02856_ ),
    .Y(\u_cpu.REG_FILE._02925_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07625_  (.A1(\u_cpu.REG_FILE.rf[16][1] ),
    .A2(\u_cpu.REG_FILE._02860_ ),
    .B1_N(\u_cpu.REG_FILE._02861_ ),
    .X(\u_cpu.REG_FILE._02926_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07626_  (.A1(\u_cpu.REG_FILE.rf[17][1] ),
    .A2(\u_cpu.REG_FILE._02859_ ),
    .B1(\u_cpu.REG_FILE._02926_ ),
    .Y(\u_cpu.REG_FILE._02927_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07627_  (.A1(\u_cpu.REG_FILE._02924_ ),
    .A2(\u_cpu.REG_FILE._02925_ ),
    .B1(\u_cpu.REG_FILE._02858_ ),
    .C1(\u_cpu.REG_FILE._02927_ ),
    .Y(\u_cpu.REG_FILE._02928_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._07628_  (.A(\u_cpu.REG_FILE.rf[22][1] ),
    .B(\u_cpu.REG_FILE._02867_ ),
    .X(\u_cpu.REG_FILE._02929_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07629_  (.A1(\u_cpu.REG_FILE.rf[23][1] ),
    .A2(\u_cpu.REG_FILE._02841_ ),
    .B1(\u_cpu.REG_FILE._02866_ ),
    .C1(\u_cpu.REG_FILE._02929_ ),
    .Y(\u_cpu.REG_FILE._02930_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07630_  (.A(\u_cpu.M_AXI_WDATA[21] ),
    .X(\u_cpu.REG_FILE._02931_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07631_  (.A1(\u_cpu.REG_FILE.rf[20][1] ),
    .A2(\u_cpu.REG_FILE._02871_ ),
    .B1_N(\u_cpu.REG_FILE._02931_ ),
    .X(\u_cpu.REG_FILE._02932_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07632_  (.A1(\u_cpu.REG_FILE.rf[21][1] ),
    .A2(\u_cpu.REG_FILE._02870_ ),
    .B1(\u_cpu.REG_FILE._02932_ ),
    .Y(\u_cpu.REG_FILE._02933_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07633_  (.A(\u_cpu.REG_FILE._02930_ ),
    .B(\u_cpu.REG_FILE._02933_ ),
    .C(\u_cpu.REG_FILE._02875_ ),
    .Y(\u_cpu.REG_FILE._02934_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07634_  (.A(\u_cpu.REG_FILE._02922_ ),
    .B(\u_cpu.REG_FILE._02928_ ),
    .C(\u_cpu.REG_FILE._02934_ ),
    .Y(\u_cpu.REG_FILE._02935_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07635_  (.A(\u_cpu.REG_FILE._02921_ ),
    .B(\u_cpu.REG_FILE._02935_ ),
    .C(\u_cpu.REG_FILE._02878_ ),
    .Y(\u_cpu.REG_FILE._02936_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07636_  (.A1(\u_cpu.REG_FILE._02746_ ),
    .A2(\u_cpu.REG_FILE._02908_ ),
    .B1(\u_cpu.REG_FILE._02936_ ),
    .C1(\u_cpu.REG_FILE._02884_ ),
    .X(\u_cpu.ALU.SrcB[1] ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07637_  (.A(\u_cpu.REG_FILE._02764_ ),
    .X(\u_cpu.REG_FILE._02937_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07638_  (.A(\u_cpu.REG_FILE.rf[19][2] ),
    .Y(\u_cpu.REG_FILE._02938_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07639_  (.A(\u_cpu.REG_FILE._02790_ ),
    .X(\u_cpu.REG_FILE._02939_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07640_  (.A(\u_cpu.REG_FILE._02810_ ),
    .X(\u_cpu.REG_FILE._02940_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07641_  (.A(\u_cpu.REG_FILE._02781_ ),
    .X(\u_cpu.REG_FILE._02941_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07642_  (.A1(\u_cpu.REG_FILE.rf[18][2] ),
    .A2(\u_cpu.REG_FILE._02940_ ),
    .B1(\u_cpu.REG_FILE._02941_ ),
    .Y(\u_cpu.REG_FILE._02942_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07643_  (.A1(\u_cpu.REG_FILE._02938_ ),
    .A2(\u_cpu.REG_FILE._02939_ ),
    .B1(\u_cpu.REG_FILE._02942_ ),
    .Y(\u_cpu.REG_FILE._02943_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07644_  (.A(\u_cpu.REG_FILE.rf[17][2] ),
    .Y(\u_cpu.REG_FILE._02944_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07645_  (.A(\u_cpu.REG_FILE._02747_ ),
    .X(\u_cpu.REG_FILE._02945_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07646_  (.A(\u_cpu.REG_FILE._02945_ ),
    .X(\u_cpu.REG_FILE._02946_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07647_  (.A(\u_cpu.REG_FILE._02750_ ),
    .X(\u_cpu.REG_FILE._02947_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07648_  (.A(\u_cpu.REG_FILE._02947_ ),
    .X(\u_cpu.REG_FILE._02948_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07649_  (.A(\u_cpu.REG_FILE._02778_ ),
    .X(\u_cpu.REG_FILE._02949_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07650_  (.A(\u_cpu.REG_FILE._02949_ ),
    .X(\u_cpu.REG_FILE._02950_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07651_  (.A(\u_cpu.REG_FILE.rf[16][2] ),
    .B(\u_cpu.REG_FILE._02950_ ),
    .Y(\u_cpu.REG_FILE._02951_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._07652_  (.A1(\u_cpu.REG_FILE._02944_ ),
    .A2(\u_cpu.REG_FILE._02946_ ),
    .B1(\u_cpu.REG_FILE._02948_ ),
    .C1(\u_cpu.REG_FILE._02951_ ),
    .Y(\u_cpu.REG_FILE._02952_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07653_  (.A(\u_cpu.REG_FILE._02792_ ),
    .X(\u_cpu.REG_FILE._02953_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07654_  (.A(\u_cpu.REG_FILE._02773_ ),
    .X(\u_cpu.REG_FILE._02954_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07655_  (.A1(\u_cpu.REG_FILE.rf[20][2] ),
    .A2(\u_cpu.REG_FILE._02953_ ),
    .B1_N(\u_cpu.REG_FILE._02954_ ),
    .Y(\u_cpu.REG_FILE._02955_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07656_  (.A(\u_cpu.REG_FILE._02758_ ),
    .X(\u_cpu.REG_FILE._02956_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07657_  (.A(\u_cpu.REG_FILE.rf[21][2] ),
    .B(\u_cpu.REG_FILE._02956_ ),
    .Y(\u_cpu.REG_FILE._02957_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07658_  (.A(\u_cpu.REG_FILE._02949_ ),
    .X(\u_cpu.REG_FILE._02958_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07659_  (.A(\u_cpu.REG_FILE.rf[22][2] ),
    .B(\u_cpu.REG_FILE._02958_ ),
    .Y(\u_cpu.REG_FILE._02959_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07660_  (.A(\u_cpu.REG_FILE._02840_ ),
    .X(\u_cpu.REG_FILE._02960_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07661_  (.A(\u_cpu.REG_FILE._02825_ ),
    .X(\u_cpu.REG_FILE._02961_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07662_  (.A1(\u_cpu.REG_FILE.rf[23][2] ),
    .A2(\u_cpu.REG_FILE._02960_ ),
    .B1(\u_cpu.REG_FILE._02961_ ),
    .Y(\u_cpu.REG_FILE._02962_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07663_  (.A(\u_cpu.REG_FILE._02803_ ),
    .X(\u_cpu.REG_FILE._02963_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._07664_  (.A1(\u_cpu.REG_FILE._02955_ ),
    .A2(\u_cpu.REG_FILE._02957_ ),
    .B1(\u_cpu.REG_FILE._02959_ ),
    .B2(\u_cpu.REG_FILE._02962_ ),
    .C1(\u_cpu.REG_FILE._02963_ ),
    .Y(\u_cpu.REG_FILE._02964_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07665_  (.A(\u_cpu.REG_FILE._02806_ ),
    .X(\u_cpu.REG_FILE._02965_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07666_  (.A(\u_cpu.REG_FILE._02965_ ),
    .X(\u_cpu.REG_FILE._02966_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.REG_FILE._07667_  (.A1(\u_cpu.REG_FILE._02937_ ),
    .A2(\u_cpu.REG_FILE._02943_ ),
    .A3(\u_cpu.REG_FILE._02952_ ),
    .B1(\u_cpu.REG_FILE._02964_ ),
    .C1(\u_cpu.REG_FILE._02966_ ),
    .X(\u_cpu.REG_FILE._02967_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07668_  (.A(\u_cpu.REG_FILE._02748_ ),
    .X(\u_cpu.REG_FILE._02968_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07669_  (.A(\u_cpu.REG_FILE._02751_ ),
    .X(\u_cpu.REG_FILE._02969_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07670_  (.A(\u_cpu.REG_FILE._02753_ ),
    .X(\u_cpu.REG_FILE._02970_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07671_  (.A(\u_cpu.REG_FILE.rf[31][2] ),
    .B_N(\u_cpu.REG_FILE._02970_ ),
    .X(\u_cpu.REG_FILE._02971_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07672_  (.A1(\u_cpu.REG_FILE.rf[30][2] ),
    .A2(\u_cpu.REG_FILE._02968_ ),
    .B1(\u_cpu.REG_FILE._02969_ ),
    .C1(\u_cpu.REG_FILE._02971_ ),
    .Y(\u_cpu.REG_FILE._02972_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07673_  (.A(\u_cpu.REG_FILE._02758_ ),
    .X(\u_cpu.REG_FILE._02973_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07674_  (.A(\u_cpu.REG_FILE._02747_ ),
    .X(\u_cpu.REG_FILE._02974_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07675_  (.A(\u_cpu.REG_FILE._02750_ ),
    .X(\u_cpu.REG_FILE._02975_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07676_  (.A1(\u_cpu.REG_FILE.rf[28][2] ),
    .A2(\u_cpu.REG_FILE._02974_ ),
    .B1_N(\u_cpu.REG_FILE._02975_ ),
    .X(\u_cpu.REG_FILE._02976_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07677_  (.A1(\u_cpu.REG_FILE.rf[29][2] ),
    .A2(\u_cpu.REG_FILE._02973_ ),
    .B1(\u_cpu.REG_FILE._02976_ ),
    .Y(\u_cpu.REG_FILE._02977_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07678_  (.A(\u_cpu.REG_FILE._02764_ ),
    .X(\u_cpu.REG_FILE._02978_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07679_  (.A(\u_cpu.REG_FILE._02972_ ),
    .B(\u_cpu.REG_FILE._02977_ ),
    .C(\u_cpu.REG_FILE._02978_ ),
    .Y(\u_cpu.REG_FILE._02979_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07680_  (.A(\u_cpu.REG_FILE._02767_ ),
    .X(\u_cpu.REG_FILE._02980_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07681_  (.A_N(\u_cpu.REG_FILE.rf[25][2] ),
    .B(\u_cpu.REG_FILE._02980_ ),
    .X(\u_cpu.REG_FILE._02981_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07682_  (.A(\u_cpu.REG_FILE._02779_ ),
    .X(\u_cpu.REG_FILE._02982_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07683_  (.A(\u_cpu.REG_FILE._02773_ ),
    .X(\u_cpu.REG_FILE._02983_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07684_  (.A1(\u_cpu.REG_FILE.rf[24][2] ),
    .A2(\u_cpu.REG_FILE._02982_ ),
    .B1_N(\u_cpu.REG_FILE._02983_ ),
    .Y(\u_cpu.REG_FILE._02984_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07685_  (.A(\u_cpu.REG_FILE._02776_ ),
    .X(\u_cpu.REG_FILE._02985_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07686_  (.A(\u_cpu.REG_FILE._02778_ ),
    .X(\u_cpu.REG_FILE._02986_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07687_  (.A(\u_cpu.REG_FILE._02986_ ),
    .X(\u_cpu.REG_FILE._02987_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07688_  (.A(\u_cpu.REG_FILE._02825_ ),
    .X(\u_cpu.REG_FILE._02988_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07689_  (.A(\u_cpu.REG_FILE.rf[27][2] ),
    .B_N(\u_cpu.REG_FILE._02949_ ),
    .X(\u_cpu.REG_FILE._02989_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07690_  (.A1(\u_cpu.REG_FILE.rf[26][2] ),
    .A2(\u_cpu.REG_FILE._02987_ ),
    .B1(\u_cpu.REG_FILE._02988_ ),
    .C1(\u_cpu.REG_FILE._02989_ ),
    .Y(\u_cpu.REG_FILE._02990_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07691_  (.A1(\u_cpu.REG_FILE._02981_ ),
    .A2(\u_cpu.REG_FILE._02984_ ),
    .B1(\u_cpu.REG_FILE._02985_ ),
    .C1(\u_cpu.REG_FILE._02990_ ),
    .Y(\u_cpu.REG_FILE._02991_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07692_  (.A(\u_cpu.REG_FILE._02787_ ),
    .X(\u_cpu.REG_FILE._02992_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07693_  (.A(\u_cpu.REG_FILE._02745_ ),
    .Y(\u_cpu.REG_FILE._02993_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07694_  (.A(\u_cpu.REG_FILE._02993_ ),
    .X(\u_cpu.REG_FILE._02994_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._07695_  (.A1(\u_cpu.REG_FILE._02979_ ),
    .A2(\u_cpu.REG_FILE._02991_ ),
    .A3(\u_cpu.REG_FILE._02992_ ),
    .B1(\u_cpu.REG_FILE._02994_ ),
    .X(\u_cpu.REG_FILE._02995_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07696_  (.A(\u_cpu.REG_FILE._02993_ ),
    .X(\u_cpu.REG_FILE._02996_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07697_  (.A(\u_cpu.REG_FILE._02996_ ),
    .X(\u_cpu.REG_FILE._02997_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07698_  (.A(\u_cpu.REG_FILE._02827_ ),
    .X(\u_cpu.REG_FILE._02998_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07699_  (.A(\u_cpu.REG_FILE.rf[14][2] ),
    .B(\u_cpu.REG_FILE._02998_ ),
    .Y(\u_cpu.REG_FILE._02999_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07700_  (.A(\u_cpu.REG_FILE._02825_ ),
    .X(\u_cpu.REG_FILE._03000_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07701_  (.A1(\u_cpu.REG_FILE.rf[15][2] ),
    .A2(\u_cpu.REG_FILE._02960_ ),
    .B1(\u_cpu.REG_FILE._03000_ ),
    .Y(\u_cpu.REG_FILE._03001_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07702_  (.A(\u_cpu.REG_FILE._02758_ ),
    .X(\u_cpu.REG_FILE._03002_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07703_  (.A(\u_cpu.REG_FILE._02770_ ),
    .X(\u_cpu.REG_FILE._03003_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07704_  (.A1(\u_cpu.REG_FILE.rf[12][2] ),
    .A2(\u_cpu.REG_FILE._03003_ ),
    .B1_N(\u_cpu.REG_FILE._02817_ ),
    .X(\u_cpu.REG_FILE._03004_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07705_  (.A1(\u_cpu.REG_FILE.rf[13][2] ),
    .A2(\u_cpu.REG_FILE._03002_ ),
    .B1(\u_cpu.REG_FILE._03004_ ),
    .Y(\u_cpu.REG_FILE._03005_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07706_  (.A(\u_cpu.REG_FILE._02803_ ),
    .X(\u_cpu.REG_FILE._03006_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07707_  (.A1(\u_cpu.REG_FILE._02999_ ),
    .A2(\u_cpu.REG_FILE._03001_ ),
    .B1(\u_cpu.REG_FILE._03005_ ),
    .C1(\u_cpu.REG_FILE._03006_ ),
    .Y(\u_cpu.REG_FILE._03007_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07708_  (.A(\u_cpu.REG_FILE._02776_ ),
    .X(\u_cpu.REG_FILE._03008_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07709_  (.A(\u_cpu.REG_FILE._03008_ ),
    .X(\u_cpu.REG_FILE._03009_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07710_  (.A(\u_cpu.REG_FILE._02867_ ),
    .X(\u_cpu.REG_FILE._03010_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07711_  (.A(\u_cpu.REG_FILE._02817_ ),
    .X(\u_cpu.REG_FILE._03011_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07712_  (.A(\u_cpu.REG_FILE._02770_ ),
    .X(\u_cpu.REG_FILE._03012_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07713_  (.A(\u_cpu.REG_FILE.rf[11][2] ),
    .B_N(\u_cpu.REG_FILE._03012_ ),
    .X(\u_cpu.REG_FILE._03013_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07714_  (.A1(\u_cpu.REG_FILE.rf[10][2] ),
    .A2(\u_cpu.REG_FILE._03010_ ),
    .B1(\u_cpu.REG_FILE._03011_ ),
    .C1(\u_cpu.REG_FILE._03013_ ),
    .Y(\u_cpu.REG_FILE._03014_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07715_  (.A(\u_cpu.REG_FILE._02840_ ),
    .X(\u_cpu.REG_FILE._03015_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07716_  (.A(\u_cpu.REG_FILE._02753_ ),
    .X(\u_cpu.REG_FILE._03016_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07717_  (.A(\u_cpu.M_AXI_WDATA[21] ),
    .X(\u_cpu.REG_FILE._03017_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07718_  (.A1(\u_cpu.REG_FILE.rf[8][2] ),
    .A2(\u_cpu.REG_FILE._03016_ ),
    .B1_N(\u_cpu.REG_FILE._03017_ ),
    .X(\u_cpu.REG_FILE._03018_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07719_  (.A1(\u_cpu.REG_FILE.rf[9][2] ),
    .A2(\u_cpu.REG_FILE._03015_ ),
    .B1(\u_cpu.REG_FILE._03018_ ),
    .Y(\u_cpu.REG_FILE._03019_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07720_  (.A(\u_cpu.REG_FILE._03009_ ),
    .B(\u_cpu.REG_FILE._03014_ ),
    .C(\u_cpu.REG_FILE._03019_ ),
    .Y(\u_cpu.REG_FILE._03020_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07721_  (.A(\u_cpu.REG_FILE._02787_ ),
    .X(\u_cpu.REG_FILE._03021_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07722_  (.A(\u_cpu.REG_FILE._03007_ ),
    .B(\u_cpu.REG_FILE._03020_ ),
    .C(\u_cpu.REG_FILE._03021_ ),
    .Y(\u_cpu.REG_FILE._03022_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07723_  (.A(\u_cpu.REG_FILE._02965_ ),
    .X(\u_cpu.REG_FILE._03023_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07724_  (.A(\u_cpu.REG_FILE._02776_ ),
    .X(\u_cpu.REG_FILE._03024_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07725_  (.A(\u_cpu.REG_FILE._02867_ ),
    .X(\u_cpu.REG_FILE._03025_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07726_  (.A(\u_cpu.REG_FILE._02817_ ),
    .X(\u_cpu.REG_FILE._03026_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07727_  (.A(\u_cpu.REG_FILE.rf[3][2] ),
    .B_N(\u_cpu.REG_FILE._02815_ ),
    .X(\u_cpu.REG_FILE._03027_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07728_  (.A1(\u_cpu.REG_FILE.rf[2][2] ),
    .A2(\u_cpu.REG_FILE._03025_ ),
    .B1(\u_cpu.REG_FILE._03026_ ),
    .C1(\u_cpu.REG_FILE._03027_ ),
    .Y(\u_cpu.REG_FILE._03028_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07729_  (.A(\u_cpu.REG_FILE._02758_ ),
    .X(\u_cpu.REG_FILE._03029_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07730_  (.A(\u_cpu.REG_FILE._02753_ ),
    .X(\u_cpu.REG_FILE._03030_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07731_  (.A1(\u_cpu.REG_FILE.rf[0][2] ),
    .A2(\u_cpu.REG_FILE._03030_ ),
    .B1_N(\u_cpu.REG_FILE._02872_ ),
    .X(\u_cpu.REG_FILE._03031_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07732_  (.A1(\u_cpu.REG_FILE.rf[1][2] ),
    .A2(\u_cpu.REG_FILE._03029_ ),
    .B1(\u_cpu.REG_FILE._03031_ ),
    .Y(\u_cpu.REG_FILE._03032_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07733_  (.A(\u_cpu.REG_FILE._03024_ ),
    .B(\u_cpu.REG_FILE._03028_ ),
    .C(\u_cpu.REG_FILE._03032_ ),
    .Y(\u_cpu.REG_FILE._03033_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07734_  (.A(\u_cpu.REG_FILE._02778_ ),
    .X(\u_cpu.REG_FILE._03034_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07735_  (.A(\u_cpu.REG_FILE.rf[7][2] ),
    .B_N(\u_cpu.REG_FILE._03034_ ),
    .X(\u_cpu.REG_FILE._03035_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07736_  (.A1(\u_cpu.REG_FILE.rf[6][2] ),
    .A2(\u_cpu.REG_FILE._02843_ ),
    .B1(\u_cpu.REG_FILE._02866_ ),
    .C1(\u_cpu.REG_FILE._03035_ ),
    .Y(\u_cpu.REG_FILE._03036_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07737_  (.A(\u_cpu.REG_FILE._02758_ ),
    .X(\u_cpu.REG_FILE._03037_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07738_  (.A(\u_cpu.REG_FILE._02753_ ),
    .X(\u_cpu.REG_FILE._03038_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07739_  (.A(\u_cpu.M_AXI_WDATA[21] ),
    .X(\u_cpu.REG_FILE._03039_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07740_  (.A1(\u_cpu.REG_FILE.rf[4][2] ),
    .A2(\u_cpu.REG_FILE._03038_ ),
    .B1_N(\u_cpu.REG_FILE._03039_ ),
    .X(\u_cpu.REG_FILE._03040_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07741_  (.A1(\u_cpu.REG_FILE.rf[5][2] ),
    .A2(\u_cpu.REG_FILE._03037_ ),
    .B1(\u_cpu.REG_FILE._03040_ ),
    .Y(\u_cpu.REG_FILE._03041_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07742_  (.A(\u_cpu.REG_FILE._02803_ ),
    .X(\u_cpu.REG_FILE._03042_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07743_  (.A(\u_cpu.REG_FILE._03036_ ),
    .B(\u_cpu.REG_FILE._03041_ ),
    .C(\u_cpu.REG_FILE._03042_ ),
    .Y(\u_cpu.REG_FILE._03043_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07744_  (.A(\u_cpu.REG_FILE._03023_ ),
    .B(\u_cpu.REG_FILE._03033_ ),
    .C(\u_cpu.REG_FILE._03043_ ),
    .Y(\u_cpu.REG_FILE._03044_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07745_  (.A(\u_cpu.REG_FILE._02997_ ),
    .B(\u_cpu.REG_FILE._03022_ ),
    .C(\u_cpu.REG_FILE._03044_ ),
    .Y(\u_cpu.REG_FILE._03045_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07746_  (.A1(\u_cpu.REG_FILE._02967_ ),
    .A2(\u_cpu.REG_FILE._02995_ ),
    .B1(\u_cpu.REG_FILE._03045_ ),
    .C1(\u_cpu.REG_FILE._02884_ ),
    .X(\u_cpu.ALU.SrcB[2] ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07747_  (.A1(\u_cpu.REG_FILE.rf[18][3] ),
    .A2(\u_cpu.REG_FILE._02940_ ),
    .B1(\u_cpu.REG_FILE._02941_ ),
    .Y(\u_cpu.REG_FILE._03046_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07748_  (.A1(\u_cpu.REG_FILE._01278_ ),
    .A2(\u_cpu.REG_FILE._02939_ ),
    .B1(\u_cpu.REG_FILE._03046_ ),
    .Y(\u_cpu.REG_FILE._03047_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07749_  (.A(\u_cpu.REG_FILE.rf[16][3] ),
    .B(\u_cpu.REG_FILE._02950_ ),
    .Y(\u_cpu.REG_FILE._03048_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._07750_  (.A1(\u_cpu.REG_FILE._01283_ ),
    .A2(\u_cpu.REG_FILE._02946_ ),
    .B1(\u_cpu.REG_FILE._02948_ ),
    .C1(\u_cpu.REG_FILE._03048_ ),
    .Y(\u_cpu.REG_FILE._03049_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07751_  (.A(\u_cpu.REG_FILE._02773_ ),
    .X(\u_cpu.REG_FILE._03050_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07752_  (.A1(\u_cpu.REG_FILE.rf[20][3] ),
    .A2(\u_cpu.REG_FILE._02953_ ),
    .B1_N(\u_cpu.REG_FILE._03050_ ),
    .Y(\u_cpu.REG_FILE._03051_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07753_  (.A(\u_cpu.REG_FILE.rf[21][3] ),
    .B(\u_cpu.REG_FILE._02956_ ),
    .Y(\u_cpu.REG_FILE._03052_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07754_  (.A(\u_cpu.REG_FILE.rf[22][3] ),
    .B(\u_cpu.REG_FILE._02958_ ),
    .Y(\u_cpu.REG_FILE._03053_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07755_  (.A1(\u_cpu.REG_FILE.rf[23][3] ),
    .A2(\u_cpu.REG_FILE._02960_ ),
    .B1(\u_cpu.REG_FILE._02961_ ),
    .Y(\u_cpu.REG_FILE._03054_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._07756_  (.A1(\u_cpu.REG_FILE._03051_ ),
    .A2(\u_cpu.REG_FILE._03052_ ),
    .B1(\u_cpu.REG_FILE._03053_ ),
    .B2(\u_cpu.REG_FILE._03054_ ),
    .C1(\u_cpu.REG_FILE._02963_ ),
    .Y(\u_cpu.REG_FILE._03055_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.REG_FILE._07757_  (.A1(\u_cpu.REG_FILE._02937_ ),
    .A2(\u_cpu.REG_FILE._03047_ ),
    .A3(\u_cpu.REG_FILE._03049_ ),
    .B1(\u_cpu.REG_FILE._03055_ ),
    .C1(\u_cpu.REG_FILE._02966_ ),
    .X(\u_cpu.REG_FILE._03056_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07758_  (.A(\u_cpu.REG_FILE._02812_ ),
    .X(\u_cpu.REG_FILE._03057_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07759_  (.A(\u_cpu.REG_FILE._02771_ ),
    .X(\u_cpu.REG_FILE._03058_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07760_  (.A(\u_cpu.REG_FILE.rf[24][3] ),
    .B(\u_cpu.REG_FILE._03058_ ),
    .Y(\u_cpu.REG_FILE._03059_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07761_  (.A(\u_cpu.REG_FILE._02747_ ),
    .X(\u_cpu.REG_FILE._03060_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07762_  (.A_N(\u_cpu.REG_FILE.rf[25][3] ),
    .B(\u_cpu.REG_FILE._03060_ ),
    .X(\u_cpu.REG_FILE._03061_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07763_  (.A(\u_cpu.REG_FILE._02776_ ),
    .X(\u_cpu.REG_FILE._03062_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07764_  (.A(\u_cpu.REG_FILE._02771_ ),
    .X(\u_cpu.REG_FILE._03063_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07765_  (.A(\u_cpu.REG_FILE._02781_ ),
    .X(\u_cpu.REG_FILE._03064_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07766_  (.A(\u_cpu.REG_FILE._02770_ ),
    .X(\u_cpu.REG_FILE._03065_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07767_  (.A(\u_cpu.REG_FILE.rf[27][3] ),
    .B_N(\u_cpu.REG_FILE._03065_ ),
    .X(\u_cpu.REG_FILE._03066_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07768_  (.A1(\u_cpu.REG_FILE.rf[26][3] ),
    .A2(\u_cpu.REG_FILE._03063_ ),
    .B1(\u_cpu.REG_FILE._03064_ ),
    .C1(\u_cpu.REG_FILE._03066_ ),
    .Y(\u_cpu.REG_FILE._03067_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._07769_  (.A1(\u_cpu.REG_FILE._03057_ ),
    .A2(\u_cpu.REG_FILE._03059_ ),
    .A3(\u_cpu.REG_FILE._03061_ ),
    .B1(\u_cpu.REG_FILE._03062_ ),
    .C1(\u_cpu.REG_FILE._03067_ ),
    .Y(\u_cpu.REG_FILE._03068_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07770_  (.A(\u_cpu.REG_FILE._02767_ ),
    .X(\u_cpu.REG_FILE._03069_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07771_  (.A_N(\u_cpu.REG_FILE.rf[29][3] ),
    .B(\u_cpu.REG_FILE._03069_ ),
    .X(\u_cpu.REG_FILE._03070_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07772_  (.A(\u_cpu.REG_FILE._03065_ ),
    .X(\u_cpu.REG_FILE._03071_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07773_  (.A(\u_cpu.REG_FILE._02773_ ),
    .X(\u_cpu.REG_FILE._03072_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07774_  (.A1(\u_cpu.REG_FILE.rf[28][3] ),
    .A2(\u_cpu.REG_FILE._03071_ ),
    .B1_N(\u_cpu.REG_FILE._03072_ ),
    .Y(\u_cpu.REG_FILE._03073_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07775_  (.A(\u_cpu.REG_FILE._02803_ ),
    .X(\u_cpu.REG_FILE._03074_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07776_  (.A(\u_cpu.REG_FILE._02783_ ),
    .X(\u_cpu.REG_FILE._03075_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07777_  (.A(\u_cpu.REG_FILE._02865_ ),
    .X(\u_cpu.REG_FILE._03076_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07778_  (.A(\u_cpu.REG_FILE._02778_ ),
    .X(\u_cpu.REG_FILE._03077_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07779_  (.A(\u_cpu.REG_FILE.rf[31][3] ),
    .B_N(\u_cpu.REG_FILE._03077_ ),
    .X(\u_cpu.REG_FILE._03078_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07780_  (.A1(\u_cpu.REG_FILE.rf[30][3] ),
    .A2(\u_cpu.REG_FILE._03075_ ),
    .B1(\u_cpu.REG_FILE._03076_ ),
    .C1(\u_cpu.REG_FILE._03078_ ),
    .Y(\u_cpu.REG_FILE._03079_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07781_  (.A1(\u_cpu.REG_FILE._03070_ ),
    .A2(\u_cpu.REG_FILE._03073_ ),
    .B1(\u_cpu.REG_FILE._03074_ ),
    .C1(\u_cpu.REG_FILE._03079_ ),
    .Y(\u_cpu.REG_FILE._03080_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07782_  (.A(\u_cpu.REG_FILE._02996_ ),
    .X(\u_cpu.REG_FILE._03081_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._07783_  (.A1(\u_cpu.REG_FILE._03068_ ),
    .A2(\u_cpu.REG_FILE._02992_ ),
    .A3(\u_cpu.REG_FILE._03080_ ),
    .B1(\u_cpu.REG_FILE._03081_ ),
    .X(\u_cpu.REG_FILE._03082_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07784_  (.A(\u_cpu.REG_FILE.rf[14][3] ),
    .B(\u_cpu.REG_FILE._02998_ ),
    .Y(\u_cpu.REG_FILE._03083_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07785_  (.A1(\u_cpu.REG_FILE.rf[15][3] ),
    .A2(\u_cpu.REG_FILE._02960_ ),
    .B1(\u_cpu.REG_FILE._03000_ ),
    .Y(\u_cpu.REG_FILE._03084_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07786_  (.A1(\u_cpu.REG_FILE.rf[12][3] ),
    .A2(\u_cpu.REG_FILE._03003_ ),
    .B1_N(\u_cpu.REG_FILE._02817_ ),
    .X(\u_cpu.REG_FILE._03085_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07787_  (.A1(\u_cpu.REG_FILE.rf[13][3] ),
    .A2(\u_cpu.REG_FILE._03002_ ),
    .B1(\u_cpu.REG_FILE._03085_ ),
    .Y(\u_cpu.REG_FILE._03086_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07788_  (.A1(\u_cpu.REG_FILE._03083_ ),
    .A2(\u_cpu.REG_FILE._03084_ ),
    .B1(\u_cpu.REG_FILE._03086_ ),
    .C1(\u_cpu.REG_FILE._03006_ ),
    .Y(\u_cpu.REG_FILE._03087_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07789_  (.A(\u_cpu.REG_FILE.rf[11][3] ),
    .B_N(\u_cpu.REG_FILE._03012_ ),
    .X(\u_cpu.REG_FILE._03088_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07790_  (.A1(\u_cpu.REG_FILE.rf[10][3] ),
    .A2(\u_cpu.REG_FILE._03010_ ),
    .B1(\u_cpu.REG_FILE._03011_ ),
    .C1(\u_cpu.REG_FILE._03088_ ),
    .Y(\u_cpu.REG_FILE._03089_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07791_  (.A(\u_cpu.REG_FILE._02753_ ),
    .X(\u_cpu.REG_FILE._03090_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07792_  (.A1(\u_cpu.REG_FILE.rf[8][3] ),
    .A2(\u_cpu.REG_FILE._03090_ ),
    .B1_N(\u_cpu.REG_FILE._03017_ ),
    .X(\u_cpu.REG_FILE._03091_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07793_  (.A1(\u_cpu.REG_FILE.rf[9][3] ),
    .A2(\u_cpu.REG_FILE._03015_ ),
    .B1(\u_cpu.REG_FILE._03091_ ),
    .Y(\u_cpu.REG_FILE._03092_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07794_  (.A(\u_cpu.REG_FILE._03009_ ),
    .B(\u_cpu.REG_FILE._03089_ ),
    .C(\u_cpu.REG_FILE._03092_ ),
    .Y(\u_cpu.REG_FILE._03093_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07795_  (.A(\u_cpu.REG_FILE._03087_ ),
    .B(\u_cpu.REG_FILE._03093_ ),
    .C(\u_cpu.REG_FILE._03021_ ),
    .Y(\u_cpu.REG_FILE._03094_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07796_  (.A(\u_cpu.REG_FILE.rf[3][3] ),
    .B_N(\u_cpu.REG_FILE._02815_ ),
    .X(\u_cpu.REG_FILE._03095_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07797_  (.A1(\u_cpu.REG_FILE.rf[2][3] ),
    .A2(\u_cpu.REG_FILE._03025_ ),
    .B1(\u_cpu.REG_FILE._03026_ ),
    .C1(\u_cpu.REG_FILE._03095_ ),
    .Y(\u_cpu.REG_FILE._03096_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07798_  (.A1(\u_cpu.REG_FILE.rf[0][3] ),
    .A2(\u_cpu.REG_FILE._03030_ ),
    .B1_N(\u_cpu.REG_FILE._02872_ ),
    .X(\u_cpu.REG_FILE._03097_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07799_  (.A1(\u_cpu.REG_FILE.rf[1][3] ),
    .A2(\u_cpu.REG_FILE._03029_ ),
    .B1(\u_cpu.REG_FILE._03097_ ),
    .Y(\u_cpu.REG_FILE._03098_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07800_  (.A(\u_cpu.REG_FILE._03009_ ),
    .B(\u_cpu.REG_FILE._03096_ ),
    .C(\u_cpu.REG_FILE._03098_ ),
    .Y(\u_cpu.REG_FILE._03099_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07801_  (.A(\u_cpu.REG_FILE.rf[7][3] ),
    .B_N(\u_cpu.REG_FILE._03034_ ),
    .X(\u_cpu.REG_FILE._03100_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07802_  (.A1(\u_cpu.REG_FILE.rf[6][3] ),
    .A2(\u_cpu.REG_FILE._02843_ ),
    .B1(\u_cpu.REG_FILE._02866_ ),
    .C1(\u_cpu.REG_FILE._03100_ ),
    .Y(\u_cpu.REG_FILE._03101_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07803_  (.A1(\u_cpu.REG_FILE.rf[4][3] ),
    .A2(\u_cpu.REG_FILE._03038_ ),
    .B1_N(\u_cpu.REG_FILE._03039_ ),
    .X(\u_cpu.REG_FILE._03102_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07804_  (.A1(\u_cpu.REG_FILE.rf[5][3] ),
    .A2(\u_cpu.REG_FILE._03037_ ),
    .B1(\u_cpu.REG_FILE._03102_ ),
    .Y(\u_cpu.REG_FILE._03103_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07805_  (.A(\u_cpu.REG_FILE._03101_ ),
    .B(\u_cpu.REG_FILE._03103_ ),
    .C(\u_cpu.REG_FILE._03042_ ),
    .Y(\u_cpu.REG_FILE._03104_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07806_  (.A(\u_cpu.REG_FILE._03023_ ),
    .B(\u_cpu.REG_FILE._03099_ ),
    .C(\u_cpu.REG_FILE._03104_ ),
    .Y(\u_cpu.REG_FILE._03105_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07807_  (.A(\u_cpu.REG_FILE._02997_ ),
    .B(\u_cpu.REG_FILE._03094_ ),
    .C(\u_cpu.REG_FILE._03105_ ),
    .Y(\u_cpu.REG_FILE._03106_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07808_  (.A1(\u_cpu.REG_FILE._03056_ ),
    .A2(\u_cpu.REG_FILE._03082_ ),
    .B1(\u_cpu.REG_FILE._03106_ ),
    .C1(\u_cpu.REG_FILE._02884_ ),
    .X(\u_cpu.ALU.SrcB[3] ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07809_  (.A1(\u_cpu.REG_FILE.rf[18][4] ),
    .A2(\u_cpu.REG_FILE._02940_ ),
    .B1(\u_cpu.REG_FILE._02941_ ),
    .Y(\u_cpu.REG_FILE._03107_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07810_  (.A1(\u_cpu.REG_FILE._01398_ ),
    .A2(\u_cpu.REG_FILE._02939_ ),
    .B1(\u_cpu.REG_FILE._03107_ ),
    .Y(\u_cpu.REG_FILE._03108_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07811_  (.A(\u_cpu.REG_FILE.rf[16][4] ),
    .B(\u_cpu.REG_FILE._02950_ ),
    .Y(\u_cpu.REG_FILE._03109_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._07812_  (.A1(\u_cpu.REG_FILE._01403_ ),
    .A2(\u_cpu.REG_FILE._02946_ ),
    .B1(\u_cpu.REG_FILE._02948_ ),
    .C1(\u_cpu.REG_FILE._03109_ ),
    .Y(\u_cpu.REG_FILE._03110_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07813_  (.A1(\u_cpu.REG_FILE.rf[20][4] ),
    .A2(\u_cpu.REG_FILE._02953_ ),
    .B1_N(\u_cpu.REG_FILE._03050_ ),
    .Y(\u_cpu.REG_FILE._03111_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07814_  (.A(\u_cpu.REG_FILE.rf[21][4] ),
    .B(\u_cpu.REG_FILE._02956_ ),
    .Y(\u_cpu.REG_FILE._03112_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07815_  (.A(\u_cpu.REG_FILE.rf[22][4] ),
    .B(\u_cpu.REG_FILE._02958_ ),
    .Y(\u_cpu.REG_FILE._03113_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07816_  (.A(\u_cpu.REG_FILE._02840_ ),
    .X(\u_cpu.REG_FILE._03114_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07817_  (.A1(\u_cpu.REG_FILE.rf[23][4] ),
    .A2(\u_cpu.REG_FILE._03114_ ),
    .B1(\u_cpu.REG_FILE._02961_ ),
    .Y(\u_cpu.REG_FILE._03115_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._07818_  (.A1(\u_cpu.REG_FILE._03111_ ),
    .A2(\u_cpu.REG_FILE._03112_ ),
    .B1(\u_cpu.REG_FILE._03113_ ),
    .B2(\u_cpu.REG_FILE._03115_ ),
    .C1(\u_cpu.REG_FILE._02963_ ),
    .Y(\u_cpu.REG_FILE._03116_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.REG_FILE._07819_  (.A1(\u_cpu.REG_FILE._02937_ ),
    .A2(\u_cpu.REG_FILE._03108_ ),
    .A3(\u_cpu.REG_FILE._03110_ ),
    .B1(\u_cpu.REG_FILE._03116_ ),
    .C1(\u_cpu.REG_FILE._02966_ ),
    .X(\u_cpu.REG_FILE._03117_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07820_  (.A(\u_cpu.REG_FILE.rf[31][4] ),
    .B_N(\u_cpu.REG_FILE._02970_ ),
    .X(\u_cpu.REG_FILE._03118_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07821_  (.A1(\u_cpu.REG_FILE.rf[30][4] ),
    .A2(\u_cpu.REG_FILE._02968_ ),
    .B1(\u_cpu.REG_FILE._02969_ ),
    .C1(\u_cpu.REG_FILE._03118_ ),
    .Y(\u_cpu.REG_FILE._03119_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07822_  (.A1(\u_cpu.REG_FILE.rf[28][4] ),
    .A2(\u_cpu.REG_FILE._02974_ ),
    .B1_N(\u_cpu.REG_FILE._02975_ ),
    .X(\u_cpu.REG_FILE._03120_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07823_  (.A1(\u_cpu.REG_FILE.rf[29][4] ),
    .A2(\u_cpu.REG_FILE._02973_ ),
    .B1(\u_cpu.REG_FILE._03120_ ),
    .Y(\u_cpu.REG_FILE._03121_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07824_  (.A(\u_cpu.REG_FILE._03119_ ),
    .B(\u_cpu.REG_FILE._03121_ ),
    .C(\u_cpu.REG_FILE._02978_ ),
    .Y(\u_cpu.REG_FILE._03122_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07825_  (.A_N(\u_cpu.REG_FILE.rf[25][4] ),
    .B(\u_cpu.REG_FILE._02980_ ),
    .X(\u_cpu.REG_FILE._03123_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07826_  (.A1(\u_cpu.REG_FILE.rf[24][4] ),
    .A2(\u_cpu.REG_FILE._02982_ ),
    .B1_N(\u_cpu.REG_FILE._02983_ ),
    .Y(\u_cpu.REG_FILE._03124_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07827_  (.A(\u_cpu.REG_FILE._02783_ ),
    .X(\u_cpu.REG_FILE._03125_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07828_  (.A(\u_cpu.REG_FILE.rf[27][4] ),
    .B_N(\u_cpu.REG_FILE._02949_ ),
    .X(\u_cpu.REG_FILE._03126_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07829_  (.A1(\u_cpu.REG_FILE.rf[26][4] ),
    .A2(\u_cpu.REG_FILE._03125_ ),
    .B1(\u_cpu.REG_FILE._02988_ ),
    .C1(\u_cpu.REG_FILE._03126_ ),
    .Y(\u_cpu.REG_FILE._03127_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07830_  (.A1(\u_cpu.REG_FILE._03123_ ),
    .A2(\u_cpu.REG_FILE._03124_ ),
    .B1(\u_cpu.REG_FILE._02985_ ),
    .C1(\u_cpu.REG_FILE._03127_ ),
    .Y(\u_cpu.REG_FILE._03128_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07831_  (.A(\u_cpu.REG_FILE._02787_ ),
    .X(\u_cpu.REG_FILE._03129_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._07832_  (.A1(\u_cpu.REG_FILE._03122_ ),
    .A2(\u_cpu.REG_FILE._03128_ ),
    .A3(\u_cpu.REG_FILE._03129_ ),
    .B1(\u_cpu.REG_FILE._03081_ ),
    .X(\u_cpu.REG_FILE._03130_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07833_  (.A(\u_cpu.REG_FILE.rf[8][4] ),
    .B(\u_cpu.REG_FILE._02998_ ),
    .Y(\u_cpu.REG_FILE._03131_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07834_  (.A(\u_cpu.REG_FILE._02840_ ),
    .X(\u_cpu.REG_FILE._03132_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07835_  (.A(\u_cpu.REG_FILE._02750_ ),
    .X(\u_cpu.REG_FILE._03133_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07836_  (.A1(\u_cpu.REG_FILE.rf[9][4] ),
    .A2(\u_cpu.REG_FILE._03132_ ),
    .B1_N(\u_cpu.REG_FILE._03133_ ),
    .Y(\u_cpu.REG_FILE._03134_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07837_  (.A(\u_cpu.REG_FILE._02776_ ),
    .X(\u_cpu.REG_FILE._03135_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07838_  (.A(\u_cpu.REG_FILE._02840_ ),
    .X(\u_cpu.REG_FILE._03136_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07839_  (.A(\u_cpu.REG_FILE._02825_ ),
    .X(\u_cpu.REG_FILE._03137_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._07840_  (.A(\u_cpu.REG_FILE.rf[10][4] ),
    .B(\u_cpu.REG_FILE._03012_ ),
    .X(\u_cpu.REG_FILE._03138_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07841_  (.A1(\u_cpu.REG_FILE.rf[11][4] ),
    .A2(\u_cpu.REG_FILE._03136_ ),
    .B1(\u_cpu.REG_FILE._03137_ ),
    .C1(\u_cpu.REG_FILE._03138_ ),
    .Y(\u_cpu.REG_FILE._03139_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07842_  (.A1(\u_cpu.REG_FILE._03131_ ),
    .A2(\u_cpu.REG_FILE._03134_ ),
    .B1(\u_cpu.REG_FILE._03135_ ),
    .C1(\u_cpu.REG_FILE._03139_ ),
    .Y(\u_cpu.REG_FILE._03140_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07843_  (.A(\u_cpu.REG_FILE._02787_ ),
    .X(\u_cpu.REG_FILE._03141_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07844_  (.A(\u_cpu.REG_FILE._02840_ ),
    .X(\u_cpu.REG_FILE._03142_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07845_  (.A(\u_cpu.REG_FILE._02770_ ),
    .X(\u_cpu.REG_FILE._03143_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._07846_  (.A(\u_cpu.REG_FILE.rf[14][4] ),
    .B(\u_cpu.REG_FILE._03143_ ),
    .X(\u_cpu.REG_FILE._03144_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07847_  (.A1(\u_cpu.REG_FILE.rf[15][4] ),
    .A2(\u_cpu.REG_FILE._03142_ ),
    .B1(\u_cpu.REG_FILE._02866_ ),
    .C1(\u_cpu.REG_FILE._03144_ ),
    .Y(\u_cpu.REG_FILE._03145_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07848_  (.A1(\u_cpu.REG_FILE.rf[12][4] ),
    .A2(\u_cpu.REG_FILE._02871_ ),
    .B1_N(\u_cpu.REG_FILE._02931_ ),
    .X(\u_cpu.REG_FILE._03146_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07849_  (.A1(\u_cpu.REG_FILE.rf[13][4] ),
    .A2(\u_cpu.REG_FILE._02870_ ),
    .B1(\u_cpu.REG_FILE._03146_ ),
    .Y(\u_cpu.REG_FILE._03147_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07850_  (.A(\u_cpu.REG_FILE._03145_ ),
    .B(\u_cpu.REG_FILE._03147_ ),
    .C(\u_cpu.REG_FILE._02875_ ),
    .Y(\u_cpu.REG_FILE._03148_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07851_  (.A(\u_cpu.REG_FILE._03140_ ),
    .B(\u_cpu.REG_FILE._03141_ ),
    .C(\u_cpu.REG_FILE._03148_ ),
    .Y(\u_cpu.REG_FILE._03149_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07852_  (.A(\u_cpu.REG_FILE.rf[3][4] ),
    .B_N(\u_cpu.REG_FILE._02815_ ),
    .X(\u_cpu.REG_FILE._03150_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07853_  (.A1(\u_cpu.REG_FILE.rf[2][4] ),
    .A2(\u_cpu.REG_FILE._03025_ ),
    .B1(\u_cpu.REG_FILE._03026_ ),
    .C1(\u_cpu.REG_FILE._03150_ ),
    .Y(\u_cpu.REG_FILE._03151_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07854_  (.A1(\u_cpu.REG_FILE.rf[0][4] ),
    .A2(\u_cpu.REG_FILE._03030_ ),
    .B1_N(\u_cpu.REG_FILE._02872_ ),
    .X(\u_cpu.REG_FILE._03152_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07855_  (.A1(\u_cpu.REG_FILE.rf[1][4] ),
    .A2(\u_cpu.REG_FILE._03029_ ),
    .B1(\u_cpu.REG_FILE._03152_ ),
    .Y(\u_cpu.REG_FILE._03153_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07856_  (.A(\u_cpu.REG_FILE._03009_ ),
    .B(\u_cpu.REG_FILE._03151_ ),
    .C(\u_cpu.REG_FILE._03153_ ),
    .Y(\u_cpu.REG_FILE._03154_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07857_  (.A(\u_cpu.REG_FILE.rf[7][4] ),
    .B_N(\u_cpu.REG_FILE._03034_ ),
    .X(\u_cpu.REG_FILE._03155_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07858_  (.A1(\u_cpu.REG_FILE.rf[6][4] ),
    .A2(\u_cpu.REG_FILE._02843_ ),
    .B1(\u_cpu.REG_FILE._02866_ ),
    .C1(\u_cpu.REG_FILE._03155_ ),
    .Y(\u_cpu.REG_FILE._03156_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07859_  (.A1(\u_cpu.REG_FILE.rf[4][4] ),
    .A2(\u_cpu.REG_FILE._03038_ ),
    .B1_N(\u_cpu.REG_FILE._03039_ ),
    .X(\u_cpu.REG_FILE._03157_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07860_  (.A1(\u_cpu.REG_FILE.rf[5][4] ),
    .A2(\u_cpu.REG_FILE._03037_ ),
    .B1(\u_cpu.REG_FILE._03157_ ),
    .Y(\u_cpu.REG_FILE._03158_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07861_  (.A(\u_cpu.REG_FILE._03156_ ),
    .B(\u_cpu.REG_FILE._03158_ ),
    .C(\u_cpu.REG_FILE._03042_ ),
    .Y(\u_cpu.REG_FILE._03159_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07862_  (.A(\u_cpu.REG_FILE._03023_ ),
    .B(\u_cpu.REG_FILE._03154_ ),
    .C(\u_cpu.REG_FILE._03159_ ),
    .Y(\u_cpu.REG_FILE._03160_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07863_  (.A(\u_cpu.REG_FILE._02997_ ),
    .B(\u_cpu.REG_FILE._03149_ ),
    .C(\u_cpu.REG_FILE._03160_ ),
    .Y(\u_cpu.REG_FILE._03161_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07864_  (.A1(\u_cpu.REG_FILE._03117_ ),
    .A2(\u_cpu.REG_FILE._03130_ ),
    .B1(\u_cpu.REG_FILE._03161_ ),
    .C1(\u_cpu.REG_FILE._02884_ ),
    .X(\u_cpu.ALU.SrcB[4] ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07865_  (.A(\u_cpu.REG_FILE.rf[19][5] ),
    .Y(\u_cpu.REG_FILE._03162_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07866_  (.A1(\u_cpu.REG_FILE.rf[18][5] ),
    .A2(\u_cpu.REG_FILE._02940_ ),
    .B1(\u_cpu.REG_FILE._02941_ ),
    .Y(\u_cpu.REG_FILE._03163_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07867_  (.A1(\u_cpu.REG_FILE._03162_ ),
    .A2(\u_cpu.REG_FILE._02939_ ),
    .B1(\u_cpu.REG_FILE._03163_ ),
    .Y(\u_cpu.REG_FILE._03164_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07868_  (.A(\u_cpu.REG_FILE.rf[17][5] ),
    .Y(\u_cpu.REG_FILE._03165_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07869_  (.A(\u_cpu.REG_FILE._02945_ ),
    .X(\u_cpu.REG_FILE._03166_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07870_  (.A(\u_cpu.REG_FILE.rf[16][5] ),
    .B(\u_cpu.REG_FILE._02950_ ),
    .Y(\u_cpu.REG_FILE._03167_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._07871_  (.A1(\u_cpu.REG_FILE._03165_ ),
    .A2(\u_cpu.REG_FILE._03166_ ),
    .B1(\u_cpu.REG_FILE._02948_ ),
    .C1(\u_cpu.REG_FILE._03167_ ),
    .Y(\u_cpu.REG_FILE._03168_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07872_  (.A1(\u_cpu.REG_FILE.rf[20][5] ),
    .A2(\u_cpu.REG_FILE._02953_ ),
    .B1_N(\u_cpu.REG_FILE._03050_ ),
    .Y(\u_cpu.REG_FILE._03169_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07873_  (.A(\u_cpu.REG_FILE.rf[21][5] ),
    .B(\u_cpu.REG_FILE._02956_ ),
    .Y(\u_cpu.REG_FILE._03170_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07874_  (.A(\u_cpu.REG_FILE.rf[22][5] ),
    .B(\u_cpu.REG_FILE._02958_ ),
    .Y(\u_cpu.REG_FILE._03171_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07875_  (.A1(\u_cpu.REG_FILE.rf[23][5] ),
    .A2(\u_cpu.REG_FILE._03114_ ),
    .B1(\u_cpu.REG_FILE._02961_ ),
    .Y(\u_cpu.REG_FILE._03172_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._07876_  (.A1(\u_cpu.REG_FILE._03169_ ),
    .A2(\u_cpu.REG_FILE._03170_ ),
    .B1(\u_cpu.REG_FILE._03171_ ),
    .B2(\u_cpu.REG_FILE._03172_ ),
    .C1(\u_cpu.REG_FILE._02963_ ),
    .Y(\u_cpu.REG_FILE._03173_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.REG_FILE._07877_  (.A1(\u_cpu.REG_FILE._02937_ ),
    .A2(\u_cpu.REG_FILE._03164_ ),
    .A3(\u_cpu.REG_FILE._03168_ ),
    .B1(\u_cpu.REG_FILE._03173_ ),
    .C1(\u_cpu.REG_FILE._02966_ ),
    .X(\u_cpu.REG_FILE._03174_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07878_  (.A(\u_cpu.REG_FILE.rf[31][5] ),
    .B_N(\u_cpu.REG_FILE._02970_ ),
    .X(\u_cpu.REG_FILE._03175_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07879_  (.A1(\u_cpu.REG_FILE.rf[30][5] ),
    .A2(\u_cpu.REG_FILE._02968_ ),
    .B1(\u_cpu.REG_FILE._02969_ ),
    .C1(\u_cpu.REG_FILE._03175_ ),
    .Y(\u_cpu.REG_FILE._03176_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07880_  (.A1(\u_cpu.REG_FILE.rf[28][5] ),
    .A2(\u_cpu.REG_FILE._02974_ ),
    .B1_N(\u_cpu.REG_FILE._02975_ ),
    .X(\u_cpu.REG_FILE._03177_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07881_  (.A1(\u_cpu.REG_FILE.rf[29][5] ),
    .A2(\u_cpu.REG_FILE._02973_ ),
    .B1(\u_cpu.REG_FILE._03177_ ),
    .Y(\u_cpu.REG_FILE._03178_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07882_  (.A(\u_cpu.REG_FILE._03176_ ),
    .B(\u_cpu.REG_FILE._03178_ ),
    .C(\u_cpu.REG_FILE._03006_ ),
    .Y(\u_cpu.REG_FILE._03179_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07883_  (.A_N(\u_cpu.REG_FILE.rf[25][5] ),
    .B(\u_cpu.REG_FILE._02980_ ),
    .X(\u_cpu.REG_FILE._03180_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07884_  (.A1(\u_cpu.REG_FILE.rf[24][5] ),
    .A2(\u_cpu.REG_FILE._02982_ ),
    .B1_N(\u_cpu.REG_FILE._02983_ ),
    .Y(\u_cpu.REG_FILE._03181_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07885_  (.A(\u_cpu.REG_FILE.rf[27][5] ),
    .B_N(\u_cpu.REG_FILE._02949_ ),
    .X(\u_cpu.REG_FILE._03182_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07886_  (.A1(\u_cpu.REG_FILE.rf[26][5] ),
    .A2(\u_cpu.REG_FILE._03125_ ),
    .B1(\u_cpu.REG_FILE._02988_ ),
    .C1(\u_cpu.REG_FILE._03182_ ),
    .Y(\u_cpu.REG_FILE._03183_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07887_  (.A1(\u_cpu.REG_FILE._03180_ ),
    .A2(\u_cpu.REG_FILE._03181_ ),
    .B1(\u_cpu.REG_FILE._02985_ ),
    .C1(\u_cpu.REG_FILE._03183_ ),
    .Y(\u_cpu.REG_FILE._03184_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._07888_  (.A1(\u_cpu.REG_FILE._03179_ ),
    .A2(\u_cpu.REG_FILE._03184_ ),
    .A3(\u_cpu.REG_FILE._03129_ ),
    .B1(\u_cpu.REG_FILE._03081_ ),
    .X(\u_cpu.REG_FILE._03185_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07889_  (.A(\u_cpu.REG_FILE.rf[14][5] ),
    .B(\u_cpu.REG_FILE._02998_ ),
    .Y(\u_cpu.REG_FILE._03186_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07890_  (.A1(\u_cpu.REG_FILE.rf[15][5] ),
    .A2(\u_cpu.REG_FILE._02960_ ),
    .B1(\u_cpu.REG_FILE._02961_ ),
    .Y(\u_cpu.REG_FILE._03187_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07891_  (.A1(\u_cpu.REG_FILE.rf[12][5] ),
    .A2(\u_cpu.REG_FILE._03003_ ),
    .B1_N(\u_cpu.REG_FILE._02817_ ),
    .X(\u_cpu.REG_FILE._03188_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07892_  (.A1(\u_cpu.REG_FILE.rf[13][5] ),
    .A2(\u_cpu.REG_FILE._03002_ ),
    .B1(\u_cpu.REG_FILE._03188_ ),
    .Y(\u_cpu.REG_FILE._03189_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07893_  (.A1(\u_cpu.REG_FILE._03186_ ),
    .A2(\u_cpu.REG_FILE._03187_ ),
    .B1(\u_cpu.REG_FILE._03189_ ),
    .C1(\u_cpu.REG_FILE._02963_ ),
    .Y(\u_cpu.REG_FILE._03190_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07894_  (.A(\u_cpu.REG_FILE.rf[11][5] ),
    .B_N(\u_cpu.REG_FILE._03012_ ),
    .X(\u_cpu.REG_FILE._03191_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07895_  (.A1(\u_cpu.REG_FILE.rf[10][5] ),
    .A2(\u_cpu.REG_FILE._03010_ ),
    .B1(\u_cpu.REG_FILE._03011_ ),
    .C1(\u_cpu.REG_FILE._03191_ ),
    .Y(\u_cpu.REG_FILE._03192_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07896_  (.A1(\u_cpu.REG_FILE.rf[8][5] ),
    .A2(\u_cpu.REG_FILE._03090_ ),
    .B1_N(\u_cpu.REG_FILE._03017_ ),
    .X(\u_cpu.REG_FILE._03193_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07897_  (.A1(\u_cpu.REG_FILE.rf[9][5] ),
    .A2(\u_cpu.REG_FILE._03015_ ),
    .B1(\u_cpu.REG_FILE._03193_ ),
    .Y(\u_cpu.REG_FILE._03194_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07898_  (.A(\u_cpu.REG_FILE._03009_ ),
    .B(\u_cpu.REG_FILE._03192_ ),
    .C(\u_cpu.REG_FILE._03194_ ),
    .Y(\u_cpu.REG_FILE._03195_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07899_  (.A(\u_cpu.REG_FILE._03190_ ),
    .B(\u_cpu.REG_FILE._03195_ ),
    .C(\u_cpu.REG_FILE._03021_ ),
    .Y(\u_cpu.REG_FILE._03196_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07900_  (.A(\u_cpu.REG_FILE.rf[7][5] ),
    .Y(\u_cpu.REG_FILE._03197_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07901_  (.A(\u_cpu.REG_FILE._02773_ ),
    .X(\u_cpu.REG_FILE._03198_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07902_  (.A1(\u_cpu.REG_FILE.rf[6][5] ),
    .A2(\u_cpu.REG_FILE._02790_ ),
    .B1(\u_cpu.REG_FILE._03198_ ),
    .Y(\u_cpu.REG_FILE._03199_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07903_  (.A1(\u_cpu.REG_FILE._03197_ ),
    .A2(\u_cpu.REG_FILE._02968_ ),
    .B1(\u_cpu.REG_FILE._03199_ ),
    .Y(\u_cpu.REG_FILE._03200_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07904_  (.A(\u_cpu.REG_FILE._02773_ ),
    .X(\u_cpu.REG_FILE._03201_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07905_  (.A1(\u_cpu.REG_FILE.rf[4][5] ),
    .A2(\u_cpu.REG_FILE._02797_ ),
    .B1_N(\u_cpu.REG_FILE._03201_ ),
    .Y(\u_cpu.REG_FILE._03202_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07906_  (.A1(\u_cpu.REG_FILE._01430_ ),
    .A2(\u_cpu.REG_FILE._02968_ ),
    .B1(\u_cpu.REG_FILE._03202_ ),
    .Y(\u_cpu.REG_FILE._03203_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07907_  (.A(\u_cpu.REG_FILE._02767_ ),
    .X(\u_cpu.REG_FILE._03204_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07908_  (.A(\u_cpu.REG_FILE.rf[0][5] ),
    .B(\u_cpu.REG_FILE._03204_ ),
    .Y(\u_cpu.REG_FILE._03205_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07909_  (.A_N(\u_cpu.REG_FILE.rf[1][5] ),
    .B(\u_cpu.REG_FILE._03090_ ),
    .X(\u_cpu.REG_FILE._03206_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07910_  (.A(\u_cpu.REG_FILE.rf[3][5] ),
    .B_N(\u_cpu.REG_FILE._02767_ ),
    .X(\u_cpu.REG_FILE._03207_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07911_  (.A1(\u_cpu.REG_FILE.rf[2][5] ),
    .A2(\u_cpu.REG_FILE._03204_ ),
    .B1(\u_cpu.REG_FILE._03133_ ),
    .C1(\u_cpu.REG_FILE._03207_ ),
    .Y(\u_cpu.REG_FILE._03208_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._07912_  (.A1(\u_cpu.REG_FILE._02826_ ),
    .A2(\u_cpu.REG_FILE._03205_ ),
    .A3(\u_cpu.REG_FILE._03206_ ),
    .B1(\u_cpu.REG_FILE._03008_ ),
    .C1(\u_cpu.REG_FILE._03208_ ),
    .Y(\u_cpu.REG_FILE._03209_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._07913_  (.A1(\u_cpu.REG_FILE._03024_ ),
    .A2(\u_cpu.REG_FILE._03200_ ),
    .A3(\u_cpu.REG_FILE._03203_ ),
    .B1(\u_cpu.REG_FILE._02965_ ),
    .C1(\u_cpu.REG_FILE._03209_ ),
    .Y(\u_cpu.REG_FILE._03210_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07914_  (.A(\u_cpu.REG_FILE._02997_ ),
    .B(\u_cpu.REG_FILE._03196_ ),
    .C(\u_cpu.REG_FILE._03210_ ),
    .Y(\u_cpu.REG_FILE._03211_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07915_  (.A1(\u_cpu.REG_FILE._03174_ ),
    .A2(\u_cpu.REG_FILE._03185_ ),
    .B1(\u_cpu.REG_FILE._03211_ ),
    .C1(\u_cpu.REG_FILE._02884_ ),
    .X(\u_cpu.ALU.SrcB[5] ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07916_  (.A(\u_cpu.REG_FILE._02779_ ),
    .X(\u_cpu.REG_FILE._03212_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07917_  (.A(\u_cpu.REG_FILE.rf[8][6] ),
    .B(\u_cpu.REG_FILE._03212_ ),
    .Y(\u_cpu.REG_FILE._03213_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07918_  (.A_N(\u_cpu.REG_FILE.rf[9][6] ),
    .B(\u_cpu.REG_FILE._02945_ ),
    .X(\u_cpu.REG_FILE._03214_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07919_  (.A(\u_cpu.REG_FILE.rf[11][6] ),
    .B_N(\u_cpu.REG_FILE._02779_ ),
    .X(\u_cpu.REG_FILE._03215_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07920_  (.A1(\u_cpu.REG_FILE.rf[10][6] ),
    .A2(\u_cpu.REG_FILE._03071_ ),
    .B1(\u_cpu.REG_FILE._02941_ ),
    .C1(\u_cpu.REG_FILE._03215_ ),
    .Y(\u_cpu.REG_FILE._03216_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._07921_  (.A1(\u_cpu.REG_FILE._03057_ ),
    .A2(\u_cpu.REG_FILE._03213_ ),
    .A3(\u_cpu.REG_FILE._03214_ ),
    .B1(\u_cpu.REG_FILE._03062_ ),
    .C1(\u_cpu.REG_FILE._03216_ ),
    .Y(\u_cpu.REG_FILE._03217_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07922_  (.A(\u_cpu.REG_FILE._02787_ ),
    .X(\u_cpu.REG_FILE._03218_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07923_  (.A_N(\u_cpu.REG_FILE.rf[13][6] ),
    .B(\u_cpu.REG_FILE._03069_ ),
    .X(\u_cpu.REG_FILE._03219_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07924_  (.A1(\u_cpu.REG_FILE.rf[12][6] ),
    .A2(\u_cpu.REG_FILE._03063_ ),
    .B1_N(\u_cpu.REG_FILE._02774_ ),
    .Y(\u_cpu.REG_FILE._03220_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07925_  (.A(\u_cpu.REG_FILE._02803_ ),
    .X(\u_cpu.REG_FILE._03221_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07926_  (.A(\u_cpu.REG_FILE.rf[15][6] ),
    .B_N(\u_cpu.REG_FILE._02783_ ),
    .X(\u_cpu.REG_FILE._03222_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07927_  (.A1(\u_cpu.REG_FILE.rf[14][6] ),
    .A2(\u_cpu.REG_FILE._02780_ ),
    .B1(\u_cpu.REG_FILE._02782_ ),
    .C1(\u_cpu.REG_FILE._03222_ ),
    .Y(\u_cpu.REG_FILE._03223_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07928_  (.A1(\u_cpu.REG_FILE._03219_ ),
    .A2(\u_cpu.REG_FILE._03220_ ),
    .B1(\u_cpu.REG_FILE._03221_ ),
    .C1(\u_cpu.REG_FILE._03223_ ),
    .Y(\u_cpu.REG_FILE._03224_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07929_  (.A(\u_cpu.REG_FILE._03217_ ),
    .B(\u_cpu.REG_FILE._03218_ ),
    .C(\u_cpu.REG_FILE._03224_ ),
    .Y(\u_cpu.REG_FILE._03225_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07930_  (.A1(\u_cpu.REG_FILE.rf[4][6] ),
    .A2(\u_cpu.REG_FILE._02793_ ),
    .B1_N(\u_cpu.REG_FILE._02794_ ),
    .Y(\u_cpu.REG_FILE._03226_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07931_  (.A1(\u_cpu.REG_FILE._01481_ ),
    .A2(\u_cpu.REG_FILE._02791_ ),
    .B1(\u_cpu.REG_FILE._03226_ ),
    .Y(\u_cpu.REG_FILE._03227_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07932_  (.A1(\u_cpu.REG_FILE.rf[6][6] ),
    .A2(\u_cpu.REG_FILE._02797_ ),
    .B1(\u_cpu.REG_FILE._02799_ ),
    .Y(\u_cpu.REG_FILE._03228_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07933_  (.A_N(\u_cpu.REG_FILE.rf[7][6] ),
    .B(\u_cpu.REG_FILE._02801_ ),
    .X(\u_cpu.REG_FILE._03229_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07934_  (.A1(\u_cpu.REG_FILE._03228_ ),
    .A2(\u_cpu.REG_FILE._03229_ ),
    .B1(\u_cpu.REG_FILE._02804_ ),
    .Y(\u_cpu.REG_FILE._03230_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07935_  (.A_N(\u_cpu.REG_FILE.rf[1][6] ),
    .B(\u_cpu.REG_FILE._02808_ ),
    .X(\u_cpu.REG_FILE._03231_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07936_  (.A1(\u_cpu.REG_FILE.rf[0][6] ),
    .A2(\u_cpu.REG_FILE._02811_ ),
    .B1_N(\u_cpu.REG_FILE._02812_ ),
    .Y(\u_cpu.REG_FILE._03232_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07937_  (.A(\u_cpu.REG_FILE.rf[3][6] ),
    .B_N(\u_cpu.REG_FILE._02771_ ),
    .X(\u_cpu.REG_FILE._03233_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07938_  (.A1(\u_cpu.REG_FILE.rf[2][6] ),
    .A2(\u_cpu.REG_FILE._02903_ ),
    .B1(\u_cpu.REG_FILE._02818_ ),
    .C1(\u_cpu.REG_FILE._03233_ ),
    .Y(\u_cpu.REG_FILE._03234_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07939_  (.A1(\u_cpu.REG_FILE._03231_ ),
    .A2(\u_cpu.REG_FILE._03232_ ),
    .B1(\u_cpu.REG_FILE._02814_ ),
    .C1(\u_cpu.REG_FILE._03234_ ),
    .Y(\u_cpu.REG_FILE._03235_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07940_  (.A1(\u_cpu.REG_FILE._03227_ ),
    .A2(\u_cpu.REG_FILE._03230_ ),
    .B1(\u_cpu.REG_FILE._02807_ ),
    .C1(\u_cpu.REG_FILE._03235_ ),
    .Y(\u_cpu.REG_FILE._03236_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._07941_  (.A(\u_cpu.REG_FILE._03225_ ),
    .B(\u_cpu.REG_FILE._03236_ ),
    .Y(\u_cpu.REG_FILE._03237_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07942_  (.A(\u_cpu.REG_FILE.rf[27][6] ),
    .B_N(\u_cpu.REG_FILE._02827_ ),
    .X(\u_cpu.REG_FILE._03238_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07943_  (.A1(\u_cpu.REG_FILE.rf[26][6] ),
    .A2(\u_cpu.REG_FILE._02824_ ),
    .B1(\u_cpu.REG_FILE._02826_ ),
    .C1(\u_cpu.REG_FILE._03238_ ),
    .X(\u_cpu.REG_FILE._03239_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07944_  (.A1(\u_cpu.REG_FILE.rf[24][6] ),
    .A2(\u_cpu.REG_FILE._02830_ ),
    .B1_N(\u_cpu.REG_FILE._02865_ ),
    .X(\u_cpu.REG_FILE._03240_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07945_  (.A(\u_cpu.REG_FILE.rf[25][6] ),
    .B_N(\u_cpu.REG_FILE._02832_ ),
    .X(\u_cpu.REG_FILE._03241_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._07946_  (.A1(\u_cpu.REG_FILE._03240_ ),
    .A2(\u_cpu.REG_FILE._03241_ ),
    .B1(\u_cpu.REG_FILE._02834_ ),
    .X(\u_cpu.REG_FILE._03242_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07947_  (.A1(\u_cpu.REG_FILE.rf[28][6] ),
    .A2(\u_cpu.REG_FILE._02837_ ),
    .B1_N(\u_cpu.REG_FILE._02838_ ),
    .Y(\u_cpu.REG_FILE._03243_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07948_  (.A(\u_cpu.REG_FILE.rf[29][6] ),
    .B(\u_cpu.REG_FILE._02841_ ),
    .Y(\u_cpu.REG_FILE._03244_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07949_  (.A(\u_cpu.REG_FILE.rf[30][6] ),
    .B(\u_cpu.REG_FILE._02916_ ),
    .Y(\u_cpu.REG_FILE._03245_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07950_  (.A1(\u_cpu.REG_FILE.rf[31][6] ),
    .A2(\u_cpu.REG_FILE._02845_ ),
    .B1(\u_cpu.REG_FILE._02846_ ),
    .Y(\u_cpu.REG_FILE._03246_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._07951_  (.A1(\u_cpu.REG_FILE._03243_ ),
    .A2(\u_cpu.REG_FILE._03244_ ),
    .B1(\u_cpu.REG_FILE._03245_ ),
    .B2(\u_cpu.REG_FILE._03246_ ),
    .C1(\u_cpu.REG_FILE._02919_ ),
    .Y(\u_cpu.REG_FILE._03247_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07952_  (.A1(\u_cpu.REG_FILE._03239_ ),
    .A2(\u_cpu.REG_FILE._03242_ ),
    .B1(\u_cpu.REG_FILE._02836_ ),
    .C1(\u_cpu.REG_FILE._03247_ ),
    .Y(\u_cpu.REG_FILE._03248_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07953_  (.A(\u_cpu.REG_FILE._02798_ ),
    .X(\u_cpu.REG_FILE._03249_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07954_  (.A1(\u_cpu.REG_FILE.rf[18][6] ),
    .A2(\u_cpu.REG_FILE._02923_ ),
    .B1(\u_cpu.REG_FILE._03249_ ),
    .Y(\u_cpu.REG_FILE._03250_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07955_  (.A(\u_cpu.REG_FILE.rf[19][6] ),
    .B(\u_cpu.REG_FILE._02856_ ),
    .Y(\u_cpu.REG_FILE._03251_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07956_  (.A1(\u_cpu.REG_FILE.rf[16][6] ),
    .A2(\u_cpu.REG_FILE._02860_ ),
    .B1_N(\u_cpu.REG_FILE._02861_ ),
    .X(\u_cpu.REG_FILE._03252_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07957_  (.A1(\u_cpu.REG_FILE.rf[17][6] ),
    .A2(\u_cpu.REG_FILE._02859_ ),
    .B1(\u_cpu.REG_FILE._03252_ ),
    .Y(\u_cpu.REG_FILE._03253_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07958_  (.A1(\u_cpu.REG_FILE._03250_ ),
    .A2(\u_cpu.REG_FILE._03251_ ),
    .B1(\u_cpu.REG_FILE._02858_ ),
    .C1(\u_cpu.REG_FILE._03253_ ),
    .Y(\u_cpu.REG_FILE._03254_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07959_  (.A(\u_cpu.REG_FILE._02781_ ),
    .X(\u_cpu.REG_FILE._03255_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._07960_  (.A(\u_cpu.REG_FILE.rf[22][6] ),
    .B(\u_cpu.REG_FILE._03143_ ),
    .X(\u_cpu.REG_FILE._03256_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07961_  (.A1(\u_cpu.REG_FILE.rf[23][6] ),
    .A2(\u_cpu.REG_FILE._03142_ ),
    .B1(\u_cpu.REG_FILE._03255_ ),
    .C1(\u_cpu.REG_FILE._03256_ ),
    .Y(\u_cpu.REG_FILE._03257_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._07962_  (.A1(\u_cpu.REG_FILE.rf[20][6] ),
    .A2(\u_cpu.REG_FILE._02871_ ),
    .B1_N(\u_cpu.REG_FILE._02931_ ),
    .X(\u_cpu.REG_FILE._03258_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07963_  (.A1(\u_cpu.REG_FILE.rf[21][6] ),
    .A2(\u_cpu.REG_FILE._02870_ ),
    .B1(\u_cpu.REG_FILE._03258_ ),
    .Y(\u_cpu.REG_FILE._03259_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07964_  (.A(\u_cpu.REG_FILE._03257_ ),
    .B(\u_cpu.REG_FILE._03259_ ),
    .C(\u_cpu.REG_FILE._02875_ ),
    .Y(\u_cpu.REG_FILE._03260_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07965_  (.A(\u_cpu.REG_FILE._02922_ ),
    .B(\u_cpu.REG_FILE._03254_ ),
    .C(\u_cpu.REG_FILE._03260_ ),
    .Y(\u_cpu.REG_FILE._03261_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07966_  (.A(\u_cpu.REG_FILE._03248_ ),
    .B(\u_cpu.REG_FILE._03261_ ),
    .C(\u_cpu.REG_FILE._02878_ ),
    .Y(\u_cpu.REG_FILE._03262_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07967_  (.A1(\u_cpu.REG_FILE._02746_ ),
    .A2(\u_cpu.REG_FILE._03237_ ),
    .B1(\u_cpu.REG_FILE._03262_ ),
    .C1(\u_cpu.REG_FILE._02884_ ),
    .X(\u_cpu.ALU.SrcB[6] ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._07968_  (.A(\u_cpu.REG_FILE.rf[12][7] ),
    .B(\u_cpu.REG_FILE._03212_ ),
    .Y(\u_cpu.REG_FILE._03263_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07969_  (.A_N(\u_cpu.REG_FILE.rf[13][7] ),
    .B(\u_cpu.REG_FILE._03060_ ),
    .X(\u_cpu.REG_FILE._03264_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07970_  (.A(\u_cpu.REG_FILE.rf[15][7] ),
    .B_N(\u_cpu.REG_FILE._02779_ ),
    .X(\u_cpu.REG_FILE._03265_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07971_  (.A1(\u_cpu.REG_FILE.rf[14][7] ),
    .A2(\u_cpu.REG_FILE._03058_ ),
    .B1(\u_cpu.REG_FILE._02941_ ),
    .C1(\u_cpu.REG_FILE._03265_ ),
    .Y(\u_cpu.REG_FILE._03266_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._07972_  (.A1(\u_cpu.REG_FILE._03057_ ),
    .A2(\u_cpu.REG_FILE._03263_ ),
    .A3(\u_cpu.REG_FILE._03264_ ),
    .B1(\u_cpu.REG_FILE._03221_ ),
    .C1(\u_cpu.REG_FILE._03266_ ),
    .Y(\u_cpu.REG_FILE._03267_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07973_  (.A_N(\u_cpu.REG_FILE.rf[9][7] ),
    .B(\u_cpu.REG_FILE._02768_ ),
    .X(\u_cpu.REG_FILE._03268_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07974_  (.A1(\u_cpu.REG_FILE.rf[8][7] ),
    .A2(\u_cpu.REG_FILE._02772_ ),
    .B1_N(\u_cpu.REG_FILE._02774_ ),
    .Y(\u_cpu.REG_FILE._03269_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07975_  (.A(\u_cpu.REG_FILE.rf[11][7] ),
    .B_N(\u_cpu.REG_FILE._02986_ ),
    .X(\u_cpu.REG_FILE._03270_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07976_  (.A1(\u_cpu.REG_FILE.rf[10][7] ),
    .A2(\u_cpu.REG_FILE._02780_ ),
    .B1(\u_cpu.REG_FILE._02782_ ),
    .C1(\u_cpu.REG_FILE._03270_ ),
    .Y(\u_cpu.REG_FILE._03271_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07977_  (.A1(\u_cpu.REG_FILE._03268_ ),
    .A2(\u_cpu.REG_FILE._03269_ ),
    .B1(\u_cpu.REG_FILE._02777_ ),
    .C1(\u_cpu.REG_FILE._03271_ ),
    .Y(\u_cpu.REG_FILE._03272_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._07978_  (.A(\u_cpu.REG_FILE._03267_ ),
    .B(\u_cpu.REG_FILE._03272_ ),
    .C(\u_cpu.REG_FILE._02788_ ),
    .Y(\u_cpu.REG_FILE._03273_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._07979_  (.A(\u_cpu.REG_FILE.rf[5][7] ),
    .Y(\u_cpu.REG_FILE._03274_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07980_  (.A1(\u_cpu.REG_FILE.rf[4][7] ),
    .A2(\u_cpu.REG_FILE._02793_ ),
    .B1_N(\u_cpu.REG_FILE._02794_ ),
    .Y(\u_cpu.REG_FILE._03275_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._07981_  (.A1(\u_cpu.REG_FILE._03274_ ),
    .A2(\u_cpu.REG_FILE._02791_ ),
    .B1(\u_cpu.REG_FILE._03275_ ),
    .Y(\u_cpu.REG_FILE._03276_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07982_  (.A1(\u_cpu.REG_FILE.rf[6][7] ),
    .A2(\u_cpu.REG_FILE._02797_ ),
    .B1(\u_cpu.REG_FILE._02799_ ),
    .Y(\u_cpu.REG_FILE._03277_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07983_  (.A_N(\u_cpu.REG_FILE.rf[7][7] ),
    .B(\u_cpu.REG_FILE._02801_ ),
    .X(\u_cpu.REG_FILE._03278_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07984_  (.A1(\u_cpu.REG_FILE._03277_ ),
    .A2(\u_cpu.REG_FILE._03278_ ),
    .B1(\u_cpu.REG_FILE._02804_ ),
    .Y(\u_cpu.REG_FILE._03279_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07985_  (.A_N(\u_cpu.REG_FILE.rf[1][7] ),
    .B(\u_cpu.REG_FILE._02808_ ),
    .X(\u_cpu.REG_FILE._03280_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07986_  (.A1(\u_cpu.REG_FILE.rf[0][7] ),
    .A2(\u_cpu.REG_FILE._02811_ ),
    .B1_N(\u_cpu.REG_FILE._02812_ ),
    .Y(\u_cpu.REG_FILE._03281_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07987_  (.A(\u_cpu.REG_FILE.rf[3][7] ),
    .B_N(\u_cpu.REG_FILE._02771_ ),
    .X(\u_cpu.REG_FILE._03282_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07988_  (.A1(\u_cpu.REG_FILE.rf[2][7] ),
    .A2(\u_cpu.REG_FILE._02903_ ),
    .B1(\u_cpu.REG_FILE._02818_ ),
    .C1(\u_cpu.REG_FILE._03282_ ),
    .Y(\u_cpu.REG_FILE._03283_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07989_  (.A1(\u_cpu.REG_FILE._03280_ ),
    .A2(\u_cpu.REG_FILE._03281_ ),
    .B1(\u_cpu.REG_FILE._02814_ ),
    .C1(\u_cpu.REG_FILE._03283_ ),
    .Y(\u_cpu.REG_FILE._03284_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._07990_  (.A1(\u_cpu.REG_FILE._03276_ ),
    .A2(\u_cpu.REG_FILE._03279_ ),
    .B1(\u_cpu.REG_FILE._02807_ ),
    .C1(\u_cpu.REG_FILE._03284_ ),
    .Y(\u_cpu.REG_FILE._03285_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._07991_  (.A(\u_cpu.REG_FILE._03273_ ),
    .B(\u_cpu.REG_FILE._03285_ ),
    .Y(\u_cpu.REG_FILE._03286_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07992_  (.A(\u_cpu.REG_FILE._02792_ ),
    .X(\u_cpu.REG_FILE._03287_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._07993_  (.A(\u_cpu.REG_FILE.rf[27][7] ),
    .B_N(\u_cpu.REG_FILE._02771_ ),
    .X(\u_cpu.REG_FILE._03288_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._07994_  (.A1(\u_cpu.REG_FILE.rf[26][7] ),
    .A2(\u_cpu.REG_FILE._03287_ ),
    .B1(\u_cpu.REG_FILE._02854_ ),
    .C1(\u_cpu.REG_FILE._03288_ ),
    .X(\u_cpu.REG_FILE._03289_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07995_  (.A1(\u_cpu.REG_FILE.rf[24][7] ),
    .A2(\u_cpu.REG_FILE._03204_ ),
    .B1_N(\u_cpu.REG_FILE._03201_ ),
    .Y(\u_cpu.REG_FILE._03290_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._07996_  (.A_N(\u_cpu.REG_FILE.rf[25][7] ),
    .B(\u_cpu.REG_FILE._02880_ ),
    .X(\u_cpu.REG_FILE._03291_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._07997_  (.A(\u_cpu.REG_FILE._02776_ ),
    .X(\u_cpu.REG_FILE._03292_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._07998_  (.A1(\u_cpu.REG_FILE._03290_ ),
    .A2(\u_cpu.REG_FILE._03291_ ),
    .B1(\u_cpu.REG_FILE._03292_ ),
    .Y(\u_cpu.REG_FILE._03293_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._07999_  (.A1(\u_cpu.REG_FILE.rf[28][7] ),
    .A2(\u_cpu.REG_FILE._02790_ ),
    .B1_N(\u_cpu.REG_FILE._02751_ ),
    .Y(\u_cpu.REG_FILE._03294_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08000_  (.A_N(\u_cpu.REG_FILE.rf[29][7] ),
    .B(\u_cpu.REG_FILE._02754_ ),
    .X(\u_cpu.REG_FILE._03295_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08001_  (.A(\u_cpu.REG_FILE.rf[30][7] ),
    .B(\u_cpu.REG_FILE._03212_ ),
    .Y(\u_cpu.REG_FILE._03296_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08002_  (.A(\u_cpu.REG_FILE._02757_ ),
    .X(\u_cpu.REG_FILE._03297_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08003_  (.A(\u_cpu.REG_FILE._02781_ ),
    .X(\u_cpu.REG_FILE._03298_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08004_  (.A1(\u_cpu.REG_FILE.rf[31][7] ),
    .A2(\u_cpu.REG_FILE._03297_ ),
    .B1(\u_cpu.REG_FILE._03298_ ),
    .Y(\u_cpu.REG_FILE._03299_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.REG_FILE._08005_  (.A1(\u_cpu.REG_FILE._03294_ ),
    .A2(\u_cpu.REG_FILE._03295_ ),
    .B1(\u_cpu.REG_FILE._03296_ ),
    .B2(\u_cpu.REG_FILE._03299_ ),
    .Y(\u_cpu.REG_FILE._03300_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._08006_  (.A1(\u_cpu.REG_FILE._03289_ ),
    .A2(\u_cpu.REG_FILE._03293_ ),
    .B1(\u_cpu.REG_FILE._03024_ ),
    .B2(\u_cpu.REG_FILE._03300_ ),
    .C1(\u_cpu.REG_FILE._03218_ ),
    .Y(\u_cpu.REG_FILE._03301_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08007_  (.A1(\u_cpu.REG_FILE.rf[18][7] ),
    .A2(\u_cpu.REG_FILE._02923_ ),
    .B1(\u_cpu.REG_FILE._03249_ ),
    .Y(\u_cpu.REG_FILE._03302_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08008_  (.A(\u_cpu.REG_FILE.rf[19][7] ),
    .B(\u_cpu.REG_FILE._02856_ ),
    .Y(\u_cpu.REG_FILE._03303_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08009_  (.A(\u_cpu.REG_FILE._02758_ ),
    .X(\u_cpu.REG_FILE._03304_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08010_  (.A1(\u_cpu.REG_FILE.rf[16][7] ),
    .A2(\u_cpu.REG_FILE._02860_ ),
    .B1_N(\u_cpu.REG_FILE._02861_ ),
    .X(\u_cpu.REG_FILE._03305_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08011_  (.A1(\u_cpu.REG_FILE.rf[17][7] ),
    .A2(\u_cpu.REG_FILE._03304_ ),
    .B1(\u_cpu.REG_FILE._03305_ ),
    .Y(\u_cpu.REG_FILE._03306_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08012_  (.A1(\u_cpu.REG_FILE._03302_ ),
    .A2(\u_cpu.REG_FILE._03303_ ),
    .B1(\u_cpu.REG_FILE._02858_ ),
    .C1(\u_cpu.REG_FILE._03306_ ),
    .Y(\u_cpu.REG_FILE._03307_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08013_  (.A(\u_cpu.REG_FILE._02751_ ),
    .X(\u_cpu.REG_FILE._03308_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08014_  (.A(\u_cpu.REG_FILE._02852_ ),
    .X(\u_cpu.REG_FILE._03309_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08015_  (.A(\u_cpu.REG_FILE.rf[20][7] ),
    .B(\u_cpu.REG_FILE._03309_ ),
    .Y(\u_cpu.REG_FILE._03310_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08016_  (.A(\u_cpu.REG_FILE._02778_ ),
    .X(\u_cpu.REG_FILE._03311_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08017_  (.A_N(\u_cpu.REG_FILE.rf[21][7] ),
    .B(\u_cpu.REG_FILE._03311_ ),
    .X(\u_cpu.REG_FILE._03312_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08018_  (.A(\u_cpu.REG_FILE.rf[23][7] ),
    .B_N(\u_cpu.REG_FILE._02852_ ),
    .X(\u_cpu.REG_FILE._03313_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08019_  (.A1(\u_cpu.REG_FILE.rf[22][7] ),
    .A2(\u_cpu.REG_FILE._02837_ ),
    .B1(\u_cpu.REG_FILE._03198_ ),
    .C1(\u_cpu.REG_FILE._03313_ ),
    .Y(\u_cpu.REG_FILE._03314_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._08020_  (.A1(\u_cpu.REG_FILE._03308_ ),
    .A2(\u_cpu.REG_FILE._03310_ ),
    .A3(\u_cpu.REG_FILE._03312_ ),
    .B1(\u_cpu.REG_FILE._02834_ ),
    .C1(\u_cpu.REG_FILE._03314_ ),
    .Y(\u_cpu.REG_FILE._03315_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08021_  (.A(\u_cpu.REG_FILE._02922_ ),
    .B(\u_cpu.REG_FILE._03307_ ),
    .C(\u_cpu.REG_FILE._03315_ ),
    .Y(\u_cpu.REG_FILE._03316_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08022_  (.A(\u_cpu.REG_FILE._03301_ ),
    .B(\u_cpu.REG_FILE._03316_ ),
    .C(\u_cpu.REG_FILE._02878_ ),
    .Y(\u_cpu.REG_FILE._03317_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08023_  (.A1(\u_cpu.REG_FILE._02746_ ),
    .A2(\u_cpu.REG_FILE._03286_ ),
    .B1(\u_cpu.REG_FILE._03317_ ),
    .C1(\u_cpu.REG_FILE._02884_ ),
    .X(\u_cpu.ALU.SrcB[7] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08024_  (.A(\u_cpu.REG_FILE.rf[15][8] ),
    .B_N(\u_cpu.REG_FILE._02754_ ),
    .X(\u_cpu.REG_FILE._03318_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08025_  (.A1(\u_cpu.REG_FILE.rf[14][8] ),
    .A2(\u_cpu.REG_FILE._02749_ ),
    .B1(\u_cpu.REG_FILE._02752_ ),
    .C1(\u_cpu.REG_FILE._03318_ ),
    .Y(\u_cpu.REG_FILE._03319_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08026_  (.A1(\u_cpu.REG_FILE.rf[12][8] ),
    .A2(\u_cpu.REG_FILE._02760_ ),
    .B1_N(\u_cpu.REG_FILE._02761_ ),
    .X(\u_cpu.REG_FILE._03320_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08027_  (.A1(\u_cpu.REG_FILE.rf[13][8] ),
    .A2(\u_cpu.REG_FILE._02759_ ),
    .B1(\u_cpu.REG_FILE._03320_ ),
    .Y(\u_cpu.REG_FILE._03321_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08028_  (.A(\u_cpu.REG_FILE._03319_ ),
    .B(\u_cpu.REG_FILE._03321_ ),
    .C(\u_cpu.REG_FILE._02978_ ),
    .Y(\u_cpu.REG_FILE._03322_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08029_  (.A_N(\u_cpu.REG_FILE.rf[9][8] ),
    .B(\u_cpu.REG_FILE._02768_ ),
    .X(\u_cpu.REG_FILE._03323_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08030_  (.A1(\u_cpu.REG_FILE.rf[8][8] ),
    .A2(\u_cpu.REG_FILE._02772_ ),
    .B1_N(\u_cpu.REG_FILE._02774_ ),
    .Y(\u_cpu.REG_FILE._03324_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08031_  (.A(\u_cpu.REG_FILE.rf[11][8] ),
    .B_N(\u_cpu.REG_FILE._02986_ ),
    .X(\u_cpu.REG_FILE._03325_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08032_  (.A1(\u_cpu.REG_FILE.rf[10][8] ),
    .A2(\u_cpu.REG_FILE._02780_ ),
    .B1(\u_cpu.REG_FILE._02782_ ),
    .C1(\u_cpu.REG_FILE._03325_ ),
    .Y(\u_cpu.REG_FILE._03326_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08033_  (.A1(\u_cpu.REG_FILE._03323_ ),
    .A2(\u_cpu.REG_FILE._03324_ ),
    .B1(\u_cpu.REG_FILE._02777_ ),
    .C1(\u_cpu.REG_FILE._03326_ ),
    .Y(\u_cpu.REG_FILE._03327_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08034_  (.A(\u_cpu.REG_FILE._03322_ ),
    .B(\u_cpu.REG_FILE._03327_ ),
    .C(\u_cpu.REG_FILE._02788_ ),
    .Y(\u_cpu.REG_FILE._03328_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08035_  (.A1(\u_cpu.REG_FILE.rf[4][8] ),
    .A2(\u_cpu.REG_FILE._02793_ ),
    .B1_N(\u_cpu.REG_FILE._02794_ ),
    .Y(\u_cpu.REG_FILE._03329_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._08036_  (.A1(\u_cpu.REG_FILE._01595_ ),
    .A2(\u_cpu.REG_FILE._02791_ ),
    .B1(\u_cpu.REG_FILE._03329_ ),
    .Y(\u_cpu.REG_FILE._03330_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08037_  (.A(\u_cpu.REG_FILE._02767_ ),
    .X(\u_cpu.REG_FILE._03331_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08038_  (.A1(\u_cpu.REG_FILE.rf[6][8] ),
    .A2(\u_cpu.REG_FILE._03331_ ),
    .B1(\u_cpu.REG_FILE._02799_ ),
    .Y(\u_cpu.REG_FILE._03332_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08039_  (.A_N(\u_cpu.REG_FILE.rf[7][8] ),
    .B(\u_cpu.REG_FILE._02801_ ),
    .X(\u_cpu.REG_FILE._03333_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08040_  (.A1(\u_cpu.REG_FILE._03332_ ),
    .A2(\u_cpu.REG_FILE._03333_ ),
    .B1(\u_cpu.REG_FILE._02804_ ),
    .Y(\u_cpu.REG_FILE._03334_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08041_  (.A_N(\u_cpu.REG_FILE.rf[1][8] ),
    .B(\u_cpu.REG_FILE._02808_ ),
    .X(\u_cpu.REG_FILE._03335_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08042_  (.A1(\u_cpu.REG_FILE.rf[0][8] ),
    .A2(\u_cpu.REG_FILE._02811_ ),
    .B1_N(\u_cpu.REG_FILE._02812_ ),
    .Y(\u_cpu.REG_FILE._03336_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08043_  (.A(\u_cpu.REG_FILE._02778_ ),
    .X(\u_cpu.REG_FILE._03337_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08044_  (.A(\u_cpu.REG_FILE.rf[3][8] ),
    .B_N(\u_cpu.REG_FILE._03337_ ),
    .X(\u_cpu.REG_FILE._03338_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08045_  (.A1(\u_cpu.REG_FILE.rf[2][8] ),
    .A2(\u_cpu.REG_FILE._02903_ ),
    .B1(\u_cpu.REG_FILE._02818_ ),
    .C1(\u_cpu.REG_FILE._03338_ ),
    .Y(\u_cpu.REG_FILE._03339_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08046_  (.A1(\u_cpu.REG_FILE._03335_ ),
    .A2(\u_cpu.REG_FILE._03336_ ),
    .B1(\u_cpu.REG_FILE._02814_ ),
    .C1(\u_cpu.REG_FILE._03339_ ),
    .Y(\u_cpu.REG_FILE._03340_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08047_  (.A1(\u_cpu.REG_FILE._03330_ ),
    .A2(\u_cpu.REG_FILE._03334_ ),
    .B1(\u_cpu.REG_FILE._02807_ ),
    .C1(\u_cpu.REG_FILE._03340_ ),
    .Y(\u_cpu.REG_FILE._03341_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._08048_  (.A(\u_cpu.REG_FILE._03328_ ),
    .B(\u_cpu.REG_FILE._03341_ ),
    .Y(\u_cpu.REG_FILE._03342_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08049_  (.A(\u_cpu.REG_FILE.rf[27][8] ),
    .B_N(\u_cpu.REG_FILE._02827_ ),
    .X(\u_cpu.REG_FILE._03343_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08050_  (.A1(\u_cpu.REG_FILE.rf[26][8] ),
    .A2(\u_cpu.REG_FILE._02824_ ),
    .B1(\u_cpu.REG_FILE._03000_ ),
    .C1(\u_cpu.REG_FILE._03343_ ),
    .X(\u_cpu.REG_FILE._03344_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08051_  (.A1(\u_cpu.REG_FILE.rf[24][8] ),
    .A2(\u_cpu.REG_FILE._02830_ ),
    .B1_N(\u_cpu.REG_FILE._02865_ ),
    .X(\u_cpu.REG_FILE._03345_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08052_  (.A(\u_cpu.REG_FILE.rf[25][8] ),
    .B_N(\u_cpu.REG_FILE._02832_ ),
    .X(\u_cpu.REG_FILE._03346_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._08053_  (.A1(\u_cpu.REG_FILE._03345_ ),
    .A2(\u_cpu.REG_FILE._03346_ ),
    .B1(\u_cpu.REG_FILE._02764_ ),
    .X(\u_cpu.REG_FILE._03347_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08054_  (.A(\u_cpu.REG_FILE.rf[30][8] ),
    .B(\u_cpu.REG_FILE._03063_ ),
    .Y(\u_cpu.REG_FILE._03348_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08055_  (.A1(\u_cpu.REG_FILE.rf[31][8] ),
    .A2(\u_cpu.REG_FILE._03297_ ),
    .B1(\u_cpu.REG_FILE._02854_ ),
    .Y(\u_cpu.REG_FILE._03349_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08056_  (.A(\u_cpu.REG_FILE.rf[28][8] ),
    .B(\u_cpu.REG_FILE._02916_ ),
    .Y(\u_cpu.REG_FILE._03350_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08057_  (.A(\u_cpu.REG_FILE._02840_ ),
    .X(\u_cpu.REG_FILE._03351_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08058_  (.A1(\u_cpu.REG_FILE.rf[29][8] ),
    .A2(\u_cpu.REG_FILE._03351_ ),
    .B1_N(\u_cpu.REG_FILE._02947_ ),
    .Y(\u_cpu.REG_FILE._03352_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._08059_  (.A1(\u_cpu.REG_FILE._03348_ ),
    .A2(\u_cpu.REG_FILE._03349_ ),
    .B1(\u_cpu.REG_FILE._03350_ ),
    .B2(\u_cpu.REG_FILE._03352_ ),
    .C1(\u_cpu.REG_FILE._02919_ ),
    .Y(\u_cpu.REG_FILE._03353_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08060_  (.A1(\u_cpu.REG_FILE._03344_ ),
    .A2(\u_cpu.REG_FILE._03347_ ),
    .B1(\u_cpu.REG_FILE._02836_ ),
    .C1(\u_cpu.REG_FILE._03353_ ),
    .Y(\u_cpu.REG_FILE._03354_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08061_  (.A1(\u_cpu.REG_FILE.rf[18][8] ),
    .A2(\u_cpu.REG_FILE._02923_ ),
    .B1(\u_cpu.REG_FILE._03249_ ),
    .Y(\u_cpu.REG_FILE._03355_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08062_  (.A(\u_cpu.REG_FILE.rf[19][8] ),
    .B(\u_cpu.REG_FILE._02856_ ),
    .Y(\u_cpu.REG_FILE._03356_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08063_  (.A1(\u_cpu.REG_FILE.rf[16][8] ),
    .A2(\u_cpu.REG_FILE._02860_ ),
    .B1_N(\u_cpu.REG_FILE._02861_ ),
    .X(\u_cpu.REG_FILE._03357_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08064_  (.A1(\u_cpu.REG_FILE.rf[17][8] ),
    .A2(\u_cpu.REG_FILE._03304_ ),
    .B1(\u_cpu.REG_FILE._03357_ ),
    .Y(\u_cpu.REG_FILE._03358_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08065_  (.A1(\u_cpu.REG_FILE._03355_ ),
    .A2(\u_cpu.REG_FILE._03356_ ),
    .B1(\u_cpu.REG_FILE._02858_ ),
    .C1(\u_cpu.REG_FILE._03358_ ),
    .Y(\u_cpu.REG_FILE._03359_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._08066_  (.A(\u_cpu.REG_FILE.rf[22][8] ),
    .B(\u_cpu.REG_FILE._03143_ ),
    .X(\u_cpu.REG_FILE._03360_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08067_  (.A1(\u_cpu.REG_FILE.rf[23][8] ),
    .A2(\u_cpu.REG_FILE._03142_ ),
    .B1(\u_cpu.REG_FILE._03255_ ),
    .C1(\u_cpu.REG_FILE._03360_ ),
    .Y(\u_cpu.REG_FILE._03361_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08068_  (.A1(\u_cpu.REG_FILE.rf[20][8] ),
    .A2(\u_cpu.REG_FILE._02871_ ),
    .B1_N(\u_cpu.REG_FILE._02931_ ),
    .X(\u_cpu.REG_FILE._03362_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08069_  (.A1(\u_cpu.REG_FILE.rf[21][8] ),
    .A2(\u_cpu.REG_FILE._02870_ ),
    .B1(\u_cpu.REG_FILE._03362_ ),
    .Y(\u_cpu.REG_FILE._03363_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08070_  (.A(\u_cpu.REG_FILE._03361_ ),
    .B(\u_cpu.REG_FILE._03363_ ),
    .C(\u_cpu.REG_FILE._02875_ ),
    .Y(\u_cpu.REG_FILE._03364_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08071_  (.A(\u_cpu.REG_FILE._02922_ ),
    .B(\u_cpu.REG_FILE._03359_ ),
    .C(\u_cpu.REG_FILE._03364_ ),
    .Y(\u_cpu.REG_FILE._03365_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08072_  (.A(\u_cpu.REG_FILE._03354_ ),
    .B(\u_cpu.REG_FILE._03365_ ),
    .C(\u_cpu.REG_FILE._02878_ ),
    .Y(\u_cpu.REG_FILE._03366_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08073_  (.A1(\u_cpu.REG_FILE._02746_ ),
    .A2(\u_cpu.REG_FILE._03342_ ),
    .B1(\u_cpu.REG_FILE._03366_ ),
    .C1(\u_cpu.REG_FILE._02884_ ),
    .X(\u_cpu.ALU.SrcB[8] ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._08074_  (.A(\u_cpu.REG_FILE.rf[19][9] ),
    .Y(\u_cpu.REG_FILE._03367_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08075_  (.A1(\u_cpu.REG_FILE.rf[18][9] ),
    .A2(\u_cpu.REG_FILE._02940_ ),
    .B1(\u_cpu.REG_FILE._02941_ ),
    .Y(\u_cpu.REG_FILE._03368_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._08076_  (.A1(\u_cpu.REG_FILE._03367_ ),
    .A2(\u_cpu.REG_FILE._02939_ ),
    .B1(\u_cpu.REG_FILE._03368_ ),
    .Y(\u_cpu.REG_FILE._03369_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._08077_  (.A(\u_cpu.REG_FILE.rf[17][9] ),
    .Y(\u_cpu.REG_FILE._03370_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08078_  (.A(\u_cpu.REG_FILE._02949_ ),
    .X(\u_cpu.REG_FILE._03371_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08079_  (.A(\u_cpu.REG_FILE.rf[16][9] ),
    .B(\u_cpu.REG_FILE._03371_ ),
    .Y(\u_cpu.REG_FILE._03372_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._08080_  (.A1(\u_cpu.REG_FILE._03370_ ),
    .A2(\u_cpu.REG_FILE._03166_ ),
    .B1(\u_cpu.REG_FILE._02948_ ),
    .C1(\u_cpu.REG_FILE._03372_ ),
    .Y(\u_cpu.REG_FILE._03373_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08081_  (.A1(\u_cpu.REG_FILE.rf[20][9] ),
    .A2(\u_cpu.REG_FILE._02953_ ),
    .B1_N(\u_cpu.REG_FILE._03050_ ),
    .Y(\u_cpu.REG_FILE._03374_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08082_  (.A(\u_cpu.REG_FILE.rf[21][9] ),
    .B(\u_cpu.REG_FILE._02956_ ),
    .Y(\u_cpu.REG_FILE._03375_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08083_  (.A(\u_cpu.REG_FILE.rf[22][9] ),
    .B(\u_cpu.REG_FILE._02958_ ),
    .Y(\u_cpu.REG_FILE._03376_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08084_  (.A(\u_cpu.REG_FILE._02825_ ),
    .X(\u_cpu.REG_FILE._03377_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08085_  (.A1(\u_cpu.REG_FILE.rf[23][9] ),
    .A2(\u_cpu.REG_FILE._03114_ ),
    .B1(\u_cpu.REG_FILE._03377_ ),
    .Y(\u_cpu.REG_FILE._03378_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._08086_  (.A1(\u_cpu.REG_FILE._03374_ ),
    .A2(\u_cpu.REG_FILE._03375_ ),
    .B1(\u_cpu.REG_FILE._03376_ ),
    .B2(\u_cpu.REG_FILE._03378_ ),
    .C1(\u_cpu.REG_FILE._02848_ ),
    .Y(\u_cpu.REG_FILE._03379_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.REG_FILE._08087_  (.A1(\u_cpu.REG_FILE._02937_ ),
    .A2(\u_cpu.REG_FILE._03369_ ),
    .A3(\u_cpu.REG_FILE._03373_ ),
    .B1(\u_cpu.REG_FILE._03379_ ),
    .C1(\u_cpu.REG_FILE._02966_ ),
    .X(\u_cpu.REG_FILE._03380_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08088_  (.A(\u_cpu.REG_FILE.rf[31][9] ),
    .B_N(\u_cpu.REG_FILE._02970_ ),
    .X(\u_cpu.REG_FILE._03381_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08089_  (.A1(\u_cpu.REG_FILE.rf[30][9] ),
    .A2(\u_cpu.REG_FILE._02749_ ),
    .B1(\u_cpu.REG_FILE._02969_ ),
    .C1(\u_cpu.REG_FILE._03381_ ),
    .Y(\u_cpu.REG_FILE._03382_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08090_  (.A1(\u_cpu.REG_FILE.rf[28][9] ),
    .A2(\u_cpu.REG_FILE._02974_ ),
    .B1_N(\u_cpu.REG_FILE._02975_ ),
    .X(\u_cpu.REG_FILE._03383_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08091_  (.A1(\u_cpu.REG_FILE.rf[29][9] ),
    .A2(\u_cpu.REG_FILE._02973_ ),
    .B1(\u_cpu.REG_FILE._03383_ ),
    .Y(\u_cpu.REG_FILE._03384_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08092_  (.A(\u_cpu.REG_FILE._03382_ ),
    .B(\u_cpu.REG_FILE._03384_ ),
    .C(\u_cpu.REG_FILE._03006_ ),
    .Y(\u_cpu.REG_FILE._03385_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08093_  (.A_N(\u_cpu.REG_FILE.rf[25][9] ),
    .B(\u_cpu.REG_FILE._02980_ ),
    .X(\u_cpu.REG_FILE._03386_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08094_  (.A1(\u_cpu.REG_FILE.rf[24][9] ),
    .A2(\u_cpu.REG_FILE._02982_ ),
    .B1_N(\u_cpu.REG_FILE._02983_ ),
    .Y(\u_cpu.REG_FILE._03387_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08095_  (.A(\u_cpu.REG_FILE.rf[27][9] ),
    .B_N(\u_cpu.REG_FILE._02949_ ),
    .X(\u_cpu.REG_FILE._03388_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08096_  (.A1(\u_cpu.REG_FILE.rf[26][9] ),
    .A2(\u_cpu.REG_FILE._03125_ ),
    .B1(\u_cpu.REG_FILE._02988_ ),
    .C1(\u_cpu.REG_FILE._03388_ ),
    .Y(\u_cpu.REG_FILE._03389_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08097_  (.A1(\u_cpu.REG_FILE._03386_ ),
    .A2(\u_cpu.REG_FILE._03387_ ),
    .B1(\u_cpu.REG_FILE._02985_ ),
    .C1(\u_cpu.REG_FILE._03389_ ),
    .Y(\u_cpu.REG_FILE._03390_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._08098_  (.A1(\u_cpu.REG_FILE._03385_ ),
    .A2(\u_cpu.REG_FILE._03390_ ),
    .A3(\u_cpu.REG_FILE._03129_ ),
    .B1(\u_cpu.REG_FILE._03081_ ),
    .X(\u_cpu.REG_FILE._03391_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08099_  (.A(\u_cpu.REG_FILE.rf[12][9] ),
    .B(\u_cpu.REG_FILE._02998_ ),
    .Y(\u_cpu.REG_FILE._03392_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08100_  (.A1(\u_cpu.REG_FILE.rf[13][9] ),
    .A2(\u_cpu.REG_FILE._03132_ ),
    .B1_N(\u_cpu.REG_FILE._03133_ ),
    .Y(\u_cpu.REG_FILE._03393_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._08101_  (.A(\u_cpu.REG_FILE.rf[14][9] ),
    .B(\u_cpu.REG_FILE._02867_ ),
    .X(\u_cpu.REG_FILE._03394_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08102_  (.A1(\u_cpu.REG_FILE.rf[15][9] ),
    .A2(\u_cpu.REG_FILE._03136_ ),
    .B1(\u_cpu.REG_FILE._03137_ ),
    .C1(\u_cpu.REG_FILE._03394_ ),
    .Y(\u_cpu.REG_FILE._03395_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08103_  (.A1(\u_cpu.REG_FILE._03392_ ),
    .A2(\u_cpu.REG_FILE._03393_ ),
    .B1(\u_cpu.REG_FILE._03042_ ),
    .C1(\u_cpu.REG_FILE._03395_ ),
    .Y(\u_cpu.REG_FILE._03396_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08104_  (.A(\u_cpu.REG_FILE.rf[8][9] ),
    .B(\u_cpu.REG_FILE._03309_ ),
    .Y(\u_cpu.REG_FILE._03397_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08105_  (.A_N(\u_cpu.REG_FILE.rf[9][9] ),
    .B(\u_cpu.REG_FILE._03311_ ),
    .X(\u_cpu.REG_FILE._03398_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08106_  (.A(\u_cpu.REG_FILE.rf[11][9] ),
    .B_N(\u_cpu.REG_FILE._02852_ ),
    .X(\u_cpu.REG_FILE._03399_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08107_  (.A1(\u_cpu.REG_FILE.rf[10][9] ),
    .A2(\u_cpu.REG_FILE._02797_ ),
    .B1(\u_cpu.REG_FILE._03198_ ),
    .C1(\u_cpu.REG_FILE._03399_ ),
    .Y(\u_cpu.REG_FILE._03400_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._08108_  (.A1(\u_cpu.REG_FILE._03308_ ),
    .A2(\u_cpu.REG_FILE._03397_ ),
    .A3(\u_cpu.REG_FILE._03398_ ),
    .B1(\u_cpu.REG_FILE._03008_ ),
    .C1(\u_cpu.REG_FILE._03400_ ),
    .Y(\u_cpu.REG_FILE._03401_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08109_  (.A(\u_cpu.REG_FILE._03396_ ),
    .B(\u_cpu.REG_FILE._03401_ ),
    .C(\u_cpu.REG_FILE._03021_ ),
    .Y(\u_cpu.REG_FILE._03402_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08110_  (.A(\u_cpu.REG_FILE._03201_ ),
    .X(\u_cpu.REG_FILE._03403_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08111_  (.A(\u_cpu.REG_FILE._02852_ ),
    .X(\u_cpu.REG_FILE._03404_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08112_  (.A(\u_cpu.REG_FILE.rf[0][9] ),
    .B(\u_cpu.REG_FILE._03404_ ),
    .Y(\u_cpu.REG_FILE._03405_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08113_  (.A_N(\u_cpu.REG_FILE.rf[1][9] ),
    .B(\u_cpu.REG_FILE._03311_ ),
    .X(\u_cpu.REG_FILE._03406_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08114_  (.A(\u_cpu.REG_FILE._02798_ ),
    .X(\u_cpu.REG_FILE._03407_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08115_  (.A(\u_cpu.REG_FILE.rf[3][9] ),
    .B_N(\u_cpu.REG_FILE._02792_ ),
    .X(\u_cpu.REG_FILE._03408_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08116_  (.A1(\u_cpu.REG_FILE.rf[2][9] ),
    .A2(\u_cpu.REG_FILE._03309_ ),
    .B1(\u_cpu.REG_FILE._03407_ ),
    .C1(\u_cpu.REG_FILE._03408_ ),
    .Y(\u_cpu.REG_FILE._03409_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._08117_  (.A1(\u_cpu.REG_FILE._03403_ ),
    .A2(\u_cpu.REG_FILE._03405_ ),
    .A3(\u_cpu.REG_FILE._03406_ ),
    .B1(\u_cpu.REG_FILE._03008_ ),
    .C1(\u_cpu.REG_FILE._03409_ ),
    .Y(\u_cpu.REG_FILE._03410_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08118_  (.A1(\u_cpu.REG_FILE.rf[4][9] ),
    .A2(\u_cpu.REG_FILE._02748_ ),
    .B1_N(\u_cpu.REG_FILE._02781_ ),
    .X(\u_cpu.REG_FILE._03411_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08119_  (.A1(\u_cpu.REG_FILE.rf[5][9] ),
    .A2(\u_cpu.REG_FILE._03002_ ),
    .B1(\u_cpu.REG_FILE._03411_ ),
    .Y(\u_cpu.REG_FILE._03412_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.REG_FILE._08120_  (.A1(\u_cpu.REG_FILE.rf[6][9] ),
    .A2(\u_cpu.REG_FILE._03003_ ),
    .B1(\u_cpu.REG_FILE._02751_ ),
    .X(\u_cpu.REG_FILE._03413_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08121_  (.A1(\u_cpu.REG_FILE.rf[7][9] ),
    .A2(\u_cpu.REG_FILE._03037_ ),
    .B1(\u_cpu.REG_FILE._03413_ ),
    .Y(\u_cpu.REG_FILE._03414_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08122_  (.A(\u_cpu.REG_FILE._03412_ ),
    .B(\u_cpu.REG_FILE._02875_ ),
    .C(\u_cpu.REG_FILE._03414_ ),
    .Y(\u_cpu.REG_FILE._03415_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08123_  (.A(\u_cpu.REG_FILE._02851_ ),
    .B(\u_cpu.REG_FILE._03410_ ),
    .C(\u_cpu.REG_FILE._03415_ ),
    .Y(\u_cpu.REG_FILE._03416_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08124_  (.A(\u_cpu.REG_FILE._02997_ ),
    .B(\u_cpu.REG_FILE._03402_ ),
    .C(\u_cpu.REG_FILE._03416_ ),
    .Y(\u_cpu.REG_FILE._03417_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08125_  (.A1(\u_cpu.REG_FILE._03380_ ),
    .A2(\u_cpu.REG_FILE._03391_ ),
    .B1(\u_cpu.REG_FILE._03417_ ),
    .C1(\u_cpu.REG_FILE._02884_ ),
    .X(\u_cpu.ALU.SrcB[9] ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08126_  (.A(\u_cpu.REG_FILE._03311_ ),
    .X(\u_cpu.REG_FILE._03418_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08127_  (.A(\u_cpu.REG_FILE.rf[15][10] ),
    .B_N(\u_cpu.REG_FILE._02754_ ),
    .X(\u_cpu.REG_FILE._03419_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08128_  (.A1(\u_cpu.REG_FILE.rf[14][10] ),
    .A2(\u_cpu.REG_FILE._03418_ ),
    .B1(\u_cpu.REG_FILE._02752_ ),
    .C1(\u_cpu.REG_FILE._03419_ ),
    .Y(\u_cpu.REG_FILE._03420_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08129_  (.A1(\u_cpu.REG_FILE.rf[12][10] ),
    .A2(\u_cpu.REG_FILE._02760_ ),
    .B1_N(\u_cpu.REG_FILE._02761_ ),
    .X(\u_cpu.REG_FILE._03421_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08130_  (.A1(\u_cpu.REG_FILE.rf[13][10] ),
    .A2(\u_cpu.REG_FILE._02759_ ),
    .B1(\u_cpu.REG_FILE._03421_ ),
    .Y(\u_cpu.REG_FILE._03422_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08131_  (.A(\u_cpu.REG_FILE._03420_ ),
    .B(\u_cpu.REG_FILE._03422_ ),
    .C(\u_cpu.REG_FILE._02978_ ),
    .Y(\u_cpu.REG_FILE._03423_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08132_  (.A_N(\u_cpu.REG_FILE.rf[9][10] ),
    .B(\u_cpu.REG_FILE._02768_ ),
    .X(\u_cpu.REG_FILE._03424_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08133_  (.A1(\u_cpu.REG_FILE.rf[8][10] ),
    .A2(\u_cpu.REG_FILE._02772_ ),
    .B1_N(\u_cpu.REG_FILE._02774_ ),
    .Y(\u_cpu.REG_FILE._03425_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08134_  (.A(\u_cpu.REG_FILE.rf[11][10] ),
    .B_N(\u_cpu.REG_FILE._02986_ ),
    .X(\u_cpu.REG_FILE._03426_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08135_  (.A1(\u_cpu.REG_FILE.rf[10][10] ),
    .A2(\u_cpu.REG_FILE._02780_ ),
    .B1(\u_cpu.REG_FILE._02782_ ),
    .C1(\u_cpu.REG_FILE._03426_ ),
    .Y(\u_cpu.REG_FILE._03427_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08136_  (.A1(\u_cpu.REG_FILE._03424_ ),
    .A2(\u_cpu.REG_FILE._03425_ ),
    .B1(\u_cpu.REG_FILE._03062_ ),
    .C1(\u_cpu.REG_FILE._03427_ ),
    .Y(\u_cpu.REG_FILE._03428_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08137_  (.A(\u_cpu.REG_FILE._03423_ ),
    .B(\u_cpu.REG_FILE._03428_ ),
    .C(\u_cpu.REG_FILE._02788_ ),
    .Y(\u_cpu.REG_FILE._03429_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08138_  (.A1(\u_cpu.REG_FILE.rf[4][10] ),
    .A2(\u_cpu.REG_FILE._02793_ ),
    .B1_N(\u_cpu.REG_FILE._02794_ ),
    .Y(\u_cpu.REG_FILE._03430_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._08139_  (.A1(\u_cpu.REG_FILE._01698_ ),
    .A2(\u_cpu.REG_FILE._02791_ ),
    .B1(\u_cpu.REG_FILE._03430_ ),
    .Y(\u_cpu.REG_FILE._03431_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08140_  (.A1(\u_cpu.REG_FILE.rf[6][10] ),
    .A2(\u_cpu.REG_FILE._03331_ ),
    .B1(\u_cpu.REG_FILE._02799_ ),
    .Y(\u_cpu.REG_FILE._03432_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08141_  (.A_N(\u_cpu.REG_FILE.rf[7][10] ),
    .B(\u_cpu.REG_FILE._02801_ ),
    .X(\u_cpu.REG_FILE._03433_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08142_  (.A(\u_cpu.REG_FILE._02803_ ),
    .X(\u_cpu.REG_FILE._03434_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08143_  (.A1(\u_cpu.REG_FILE._03432_ ),
    .A2(\u_cpu.REG_FILE._03433_ ),
    .B1(\u_cpu.REG_FILE._03434_ ),
    .Y(\u_cpu.REG_FILE._03435_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08144_  (.A_N(\u_cpu.REG_FILE.rf[1][10] ),
    .B(\u_cpu.REG_FILE._02808_ ),
    .X(\u_cpu.REG_FILE._03436_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08145_  (.A1(\u_cpu.REG_FILE.rf[0][10] ),
    .A2(\u_cpu.REG_FILE._02811_ ),
    .B1_N(\u_cpu.REG_FILE._02812_ ),
    .Y(\u_cpu.REG_FILE._03437_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08146_  (.A(\u_cpu.REG_FILE.rf[3][10] ),
    .B_N(\u_cpu.REG_FILE._03337_ ),
    .X(\u_cpu.REG_FILE._03438_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08147_  (.A1(\u_cpu.REG_FILE.rf[2][10] ),
    .A2(\u_cpu.REG_FILE._02903_ ),
    .B1(\u_cpu.REG_FILE._02818_ ),
    .C1(\u_cpu.REG_FILE._03438_ ),
    .Y(\u_cpu.REG_FILE._03439_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08148_  (.A1(\u_cpu.REG_FILE._03436_ ),
    .A2(\u_cpu.REG_FILE._03437_ ),
    .B1(\u_cpu.REG_FILE._02814_ ),
    .C1(\u_cpu.REG_FILE._03439_ ),
    .Y(\u_cpu.REG_FILE._03440_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08149_  (.A1(\u_cpu.REG_FILE._03431_ ),
    .A2(\u_cpu.REG_FILE._03435_ ),
    .B1(\u_cpu.REG_FILE._02807_ ),
    .C1(\u_cpu.REG_FILE._03440_ ),
    .Y(\u_cpu.REG_FILE._03441_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._08150_  (.A(\u_cpu.REG_FILE._03429_ ),
    .B(\u_cpu.REG_FILE._03441_ ),
    .Y(\u_cpu.REG_FILE._03442_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08151_  (.A(\u_cpu.REG_FILE.rf[27][10] ),
    .B_N(\u_cpu.REG_FILE._02827_ ),
    .X(\u_cpu.REG_FILE._03443_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08152_  (.A1(\u_cpu.REG_FILE.rf[26][10] ),
    .A2(\u_cpu.REG_FILE._02824_ ),
    .B1(\u_cpu.REG_FILE._03000_ ),
    .C1(\u_cpu.REG_FILE._03443_ ),
    .X(\u_cpu.REG_FILE._03444_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08153_  (.A(\u_cpu.REG_FILE._02753_ ),
    .X(\u_cpu.REG_FILE._03445_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08154_  (.A1(\u_cpu.REG_FILE.rf[24][10] ),
    .A2(\u_cpu.REG_FILE._03445_ ),
    .B1_N(\u_cpu.REG_FILE._02865_ ),
    .X(\u_cpu.REG_FILE._03446_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08155_  (.A(\u_cpu.REG_FILE.rf[25][10] ),
    .B_N(\u_cpu.REG_FILE._02832_ ),
    .X(\u_cpu.REG_FILE._03447_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._08156_  (.A1(\u_cpu.REG_FILE._03446_ ),
    .A2(\u_cpu.REG_FILE._03447_ ),
    .B1(\u_cpu.REG_FILE._02764_ ),
    .X(\u_cpu.REG_FILE._03448_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08157_  (.A1(\u_cpu.REG_FILE.rf[28][10] ),
    .A2(\u_cpu.REG_FILE._02837_ ),
    .B1_N(\u_cpu.REG_FILE._02838_ ),
    .Y(\u_cpu.REG_FILE._03449_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08158_  (.A(\u_cpu.REG_FILE.rf[29][10] ),
    .B(\u_cpu.REG_FILE._02841_ ),
    .Y(\u_cpu.REG_FILE._03450_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08159_  (.A(\u_cpu.REG_FILE.rf[30][10] ),
    .B(\u_cpu.REG_FILE._02916_ ),
    .Y(\u_cpu.REG_FILE._03451_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08160_  (.A1(\u_cpu.REG_FILE.rf[31][10] ),
    .A2(\u_cpu.REG_FILE._02845_ ),
    .B1(\u_cpu.REG_FILE._02846_ ),
    .Y(\u_cpu.REG_FILE._03452_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._08161_  (.A1(\u_cpu.REG_FILE._03449_ ),
    .A2(\u_cpu.REG_FILE._03450_ ),
    .B1(\u_cpu.REG_FILE._03451_ ),
    .B2(\u_cpu.REG_FILE._03452_ ),
    .C1(\u_cpu.REG_FILE._02919_ ),
    .Y(\u_cpu.REG_FILE._03453_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08162_  (.A1(\u_cpu.REG_FILE._03444_ ),
    .A2(\u_cpu.REG_FILE._03448_ ),
    .B1(\u_cpu.REG_FILE._02836_ ),
    .C1(\u_cpu.REG_FILE._03453_ ),
    .Y(\u_cpu.REG_FILE._03454_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08163_  (.A1(\u_cpu.REG_FILE.rf[18][10] ),
    .A2(\u_cpu.REG_FILE._02923_ ),
    .B1(\u_cpu.REG_FILE._03249_ ),
    .Y(\u_cpu.REG_FILE._03455_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08164_  (.A(\u_cpu.REG_FILE.rf[19][10] ),
    .B(\u_cpu.REG_FILE._02856_ ),
    .Y(\u_cpu.REG_FILE._03456_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08165_  (.A1(\u_cpu.REG_FILE.rf[16][10] ),
    .A2(\u_cpu.REG_FILE._02860_ ),
    .B1_N(\u_cpu.REG_FILE._02861_ ),
    .X(\u_cpu.REG_FILE._03457_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08166_  (.A1(\u_cpu.REG_FILE.rf[17][10] ),
    .A2(\u_cpu.REG_FILE._03304_ ),
    .B1(\u_cpu.REG_FILE._03457_ ),
    .Y(\u_cpu.REG_FILE._03458_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08167_  (.A1(\u_cpu.REG_FILE._03455_ ),
    .A2(\u_cpu.REG_FILE._03456_ ),
    .B1(\u_cpu.REG_FILE._02858_ ),
    .C1(\u_cpu.REG_FILE._03458_ ),
    .Y(\u_cpu.REG_FILE._03459_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._08168_  (.A(\u_cpu.REG_FILE.rf[22][10] ),
    .B(\u_cpu.REG_FILE._03143_ ),
    .X(\u_cpu.REG_FILE._03460_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08169_  (.A1(\u_cpu.REG_FILE.rf[23][10] ),
    .A2(\u_cpu.REG_FILE._03142_ ),
    .B1(\u_cpu.REG_FILE._03255_ ),
    .C1(\u_cpu.REG_FILE._03460_ ),
    .Y(\u_cpu.REG_FILE._03461_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08170_  (.A1(\u_cpu.REG_FILE.rf[20][10] ),
    .A2(\u_cpu.REG_FILE._02871_ ),
    .B1_N(\u_cpu.REG_FILE._02931_ ),
    .X(\u_cpu.REG_FILE._03462_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08171_  (.A1(\u_cpu.REG_FILE.rf[21][10] ),
    .A2(\u_cpu.REG_FILE._02870_ ),
    .B1(\u_cpu.REG_FILE._03462_ ),
    .Y(\u_cpu.REG_FILE._03463_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08172_  (.A(\u_cpu.REG_FILE._03461_ ),
    .B(\u_cpu.REG_FILE._03463_ ),
    .C(\u_cpu.REG_FILE._02875_ ),
    .Y(\u_cpu.REG_FILE._03464_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08173_  (.A(\u_cpu.REG_FILE._02922_ ),
    .B(\u_cpu.REG_FILE._03459_ ),
    .C(\u_cpu.REG_FILE._03464_ ),
    .Y(\u_cpu.REG_FILE._03465_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08174_  (.A(\u_cpu.REG_FILE._03454_ ),
    .B(\u_cpu.REG_FILE._03465_ ),
    .C(\u_cpu.REG_FILE._02878_ ),
    .Y(\u_cpu.REG_FILE._03466_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08175_  (.A(\u_cpu.REG_FILE._02883_ ),
    .X(\u_cpu.REG_FILE._03467_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08176_  (.A1(\u_cpu.REG_FILE._02746_ ),
    .A2(\u_cpu.REG_FILE._03442_ ),
    .B1(\u_cpu.REG_FILE._03466_ ),
    .C1(\u_cpu.REG_FILE._03467_ ),
    .X(\u_cpu.ALU.SrcB[10] ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08177_  (.A1(\u_cpu.REG_FILE.rf[16][11] ),
    .A2(\u_cpu.REG_FILE._02790_ ),
    .B1_N(\u_cpu.REG_FILE._02751_ ),
    .Y(\u_cpu.REG_FILE._03468_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08178_  (.A_N(\u_cpu.REG_FILE.rf[17][11] ),
    .B(\u_cpu.REG_FILE._03445_ ),
    .X(\u_cpu.REG_FILE._03469_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08179_  (.A(\u_cpu.REG_FILE._02798_ ),
    .X(\u_cpu.REG_FILE._03470_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08180_  (.A1(\u_cpu.REG_FILE.rf[18][11] ),
    .A2(\u_cpu.REG_FILE._03404_ ),
    .B1(\u_cpu.REG_FILE._03470_ ),
    .Y(\u_cpu.REG_FILE._03471_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08181_  (.A_N(\u_cpu.REG_FILE.rf[19][11] ),
    .B(\u_cpu.REG_FILE._02790_ ),
    .X(\u_cpu.REG_FILE._03472_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.REG_FILE._08182_  (.A1(\u_cpu.REG_FILE._03468_ ),
    .A2(\u_cpu.REG_FILE._03469_ ),
    .B1(\u_cpu.REG_FILE._03471_ ),
    .B2(\u_cpu.REG_FILE._03472_ ),
    .Y(\u_cpu.REG_FILE._03473_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08183_  (.A(\u_cpu.REG_FILE.rf[23][11] ),
    .B_N(\u_cpu.REG_FILE._03003_ ),
    .X(\u_cpu.REG_FILE._03474_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08184_  (.A1(\u_cpu.REG_FILE.rf[22][11] ),
    .A2(\u_cpu.REG_FILE._02987_ ),
    .B1(\u_cpu.REG_FILE._02826_ ),
    .C1(\u_cpu.REG_FILE._03474_ ),
    .X(\u_cpu.REG_FILE._03475_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08185_  (.A(\u_cpu.REG_FILE.rf[20][11] ),
    .B(\u_cpu.REG_FILE._02940_ ),
    .Y(\u_cpu.REG_FILE._03476_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08186_  (.A_N(\u_cpu.REG_FILE.rf[21][11] ),
    .B(\u_cpu.REG_FILE._02880_ ),
    .X(\u_cpu.REG_FILE._03477_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.REG_FILE._08187_  (.A1(\u_cpu.REG_FILE._03403_ ),
    .A2(\u_cpu.REG_FILE._03476_ ),
    .A3(\u_cpu.REG_FILE._03477_ ),
    .B1(\u_cpu.REG_FILE._03221_ ),
    .Y(\u_cpu.REG_FILE._03478_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.REG_FILE._08188_  (.A1(\u_cpu.REG_FILE._02937_ ),
    .A2(\u_cpu.REG_FILE._03473_ ),
    .B1(\u_cpu.REG_FILE._03475_ ),
    .B2(\u_cpu.REG_FILE._03478_ ),
    .C1(\u_cpu.REG_FILE._03023_ ),
    .X(\u_cpu.REG_FILE._03479_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08189_  (.A(\u_cpu.REG_FILE.rf[28][11] ),
    .B(\u_cpu.REG_FILE._03058_ ),
    .Y(\u_cpu.REG_FILE._03480_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08190_  (.A_N(\u_cpu.REG_FILE.rf[29][11] ),
    .B(\u_cpu.REG_FILE._03060_ ),
    .X(\u_cpu.REG_FILE._03481_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08191_  (.A(\u_cpu.REG_FILE.rf[31][11] ),
    .B_N(\u_cpu.REG_FILE._03065_ ),
    .X(\u_cpu.REG_FILE._03482_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08192_  (.A1(\u_cpu.REG_FILE.rf[30][11] ),
    .A2(\u_cpu.REG_FILE._03063_ ),
    .B1(\u_cpu.REG_FILE._03064_ ),
    .C1(\u_cpu.REG_FILE._03482_ ),
    .Y(\u_cpu.REG_FILE._03483_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._08193_  (.A1(\u_cpu.REG_FILE._03057_ ),
    .A2(\u_cpu.REG_FILE._03480_ ),
    .A3(\u_cpu.REG_FILE._03481_ ),
    .B1(\u_cpu.REG_FILE._03221_ ),
    .C1(\u_cpu.REG_FILE._03483_ ),
    .Y(\u_cpu.REG_FILE._03484_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08194_  (.A_N(\u_cpu.REG_FILE.rf[25][11] ),
    .B(\u_cpu.REG_FILE._02980_ ),
    .X(\u_cpu.REG_FILE._03485_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08195_  (.A1(\u_cpu.REG_FILE.rf[24][11] ),
    .A2(\u_cpu.REG_FILE._02982_ ),
    .B1_N(\u_cpu.REG_FILE._02983_ ),
    .Y(\u_cpu.REG_FILE._03486_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08196_  (.A(\u_cpu.REG_FILE.rf[27][11] ),
    .B_N(\u_cpu.REG_FILE._03077_ ),
    .X(\u_cpu.REG_FILE._03487_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08197_  (.A1(\u_cpu.REG_FILE.rf[26][11] ),
    .A2(\u_cpu.REG_FILE._03125_ ),
    .B1(\u_cpu.REG_FILE._02988_ ),
    .C1(\u_cpu.REG_FILE._03487_ ),
    .Y(\u_cpu.REG_FILE._03488_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08198_  (.A1(\u_cpu.REG_FILE._03485_ ),
    .A2(\u_cpu.REG_FILE._03486_ ),
    .B1(\u_cpu.REG_FILE._02985_ ),
    .C1(\u_cpu.REG_FILE._03488_ ),
    .Y(\u_cpu.REG_FILE._03489_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._08199_  (.A1(\u_cpu.REG_FILE._03484_ ),
    .A2(\u_cpu.REG_FILE._03489_ ),
    .A3(\u_cpu.REG_FILE._03129_ ),
    .B1(\u_cpu.REG_FILE._03081_ ),
    .X(\u_cpu.REG_FILE._03490_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08200_  (.A(\u_cpu.REG_FILE.rf[14][11] ),
    .B(\u_cpu.REG_FILE._02998_ ),
    .Y(\u_cpu.REG_FILE._03491_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08201_  (.A1(\u_cpu.REG_FILE.rf[15][11] ),
    .A2(\u_cpu.REG_FILE._02960_ ),
    .B1(\u_cpu.REG_FILE._02961_ ),
    .Y(\u_cpu.REG_FILE._03492_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08202_  (.A1(\u_cpu.REG_FILE.rf[12][11] ),
    .A2(\u_cpu.REG_FILE._03003_ ),
    .B1_N(\u_cpu.REG_FILE._02817_ ),
    .X(\u_cpu.REG_FILE._03493_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08203_  (.A1(\u_cpu.REG_FILE.rf[13][11] ),
    .A2(\u_cpu.REG_FILE._03002_ ),
    .B1(\u_cpu.REG_FILE._03493_ ),
    .Y(\u_cpu.REG_FILE._03494_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08204_  (.A1(\u_cpu.REG_FILE._03491_ ),
    .A2(\u_cpu.REG_FILE._03492_ ),
    .B1(\u_cpu.REG_FILE._03494_ ),
    .C1(\u_cpu.REG_FILE._02963_ ),
    .Y(\u_cpu.REG_FILE._03495_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08205_  (.A(\u_cpu.REG_FILE.rf[11][11] ),
    .B_N(\u_cpu.REG_FILE._03012_ ),
    .X(\u_cpu.REG_FILE._03496_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08206_  (.A1(\u_cpu.REG_FILE.rf[10][11] ),
    .A2(\u_cpu.REG_FILE._03010_ ),
    .B1(\u_cpu.REG_FILE._03011_ ),
    .C1(\u_cpu.REG_FILE._03496_ ),
    .Y(\u_cpu.REG_FILE._03497_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08207_  (.A1(\u_cpu.REG_FILE.rf[8][11] ),
    .A2(\u_cpu.REG_FILE._03090_ ),
    .B1_N(\u_cpu.REG_FILE._03017_ ),
    .X(\u_cpu.REG_FILE._03498_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08208_  (.A1(\u_cpu.REG_FILE.rf[9][11] ),
    .A2(\u_cpu.REG_FILE._03015_ ),
    .B1(\u_cpu.REG_FILE._03498_ ),
    .Y(\u_cpu.REG_FILE._03499_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08209_  (.A(\u_cpu.REG_FILE._03135_ ),
    .B(\u_cpu.REG_FILE._03497_ ),
    .C(\u_cpu.REG_FILE._03499_ ),
    .Y(\u_cpu.REG_FILE._03500_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08210_  (.A(\u_cpu.REG_FILE._03495_ ),
    .B(\u_cpu.REG_FILE._03500_ ),
    .C(\u_cpu.REG_FILE._03021_ ),
    .Y(\u_cpu.REG_FILE._03501_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08211_  (.A(\u_cpu.REG_FILE.rf[0][11] ),
    .B(\u_cpu.REG_FILE._03309_ ),
    .Y(\u_cpu.REG_FILE._03502_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08212_  (.A_N(\u_cpu.REG_FILE.rf[1][11] ),
    .B(\u_cpu.REG_FILE._03311_ ),
    .X(\u_cpu.REG_FILE._03503_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08213_  (.A(\u_cpu.REG_FILE.rf[3][11] ),
    .B_N(\u_cpu.REG_FILE._02852_ ),
    .X(\u_cpu.REG_FILE._03504_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08214_  (.A1(\u_cpu.REG_FILE.rf[2][11] ),
    .A2(\u_cpu.REG_FILE._03309_ ),
    .B1(\u_cpu.REG_FILE._03407_ ),
    .C1(\u_cpu.REG_FILE._03504_ ),
    .Y(\u_cpu.REG_FILE._03505_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._08215_  (.A1(\u_cpu.REG_FILE._03308_ ),
    .A2(\u_cpu.REG_FILE._03502_ ),
    .A3(\u_cpu.REG_FILE._03503_ ),
    .B1(\u_cpu.REG_FILE._03008_ ),
    .C1(\u_cpu.REG_FILE._03505_ ),
    .Y(\u_cpu.REG_FILE._03506_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08216_  (.A(\u_cpu.REG_FILE.rf[4][11] ),
    .B(\u_cpu.REG_FILE._03404_ ),
    .Y(\u_cpu.REG_FILE._03507_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08217_  (.A_N(\u_cpu.REG_FILE.rf[5][11] ),
    .B(\u_cpu.REG_FILE._02748_ ),
    .X(\u_cpu.REG_FILE._03508_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.REG_FILE._08218_  (.A1(\u_cpu.REG_FILE.rf[6][11] ),
    .A2(\u_cpu.REG_FILE._02779_ ),
    .B1(\u_cpu.REG_FILE._02781_ ),
    .X(\u_cpu.REG_FILE._03509_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08219_  (.A1(\u_cpu.REG_FILE.rf[7][11] ),
    .A2(\u_cpu.REG_FILE._03351_ ),
    .B1(\u_cpu.REG_FILE._03509_ ),
    .Y(\u_cpu.REG_FILE._03510_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._08220_  (.A1(\u_cpu.REG_FILE._03403_ ),
    .A2(\u_cpu.REG_FILE._03507_ ),
    .A3(\u_cpu.REG_FILE._03508_ ),
    .B1(\u_cpu.REG_FILE._02834_ ),
    .C1(\u_cpu.REG_FILE._03510_ ),
    .Y(\u_cpu.REG_FILE._03511_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08221_  (.A(\u_cpu.REG_FILE._02851_ ),
    .B(\u_cpu.REG_FILE._03506_ ),
    .C(\u_cpu.REG_FILE._03511_ ),
    .Y(\u_cpu.REG_FILE._03512_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08222_  (.A(\u_cpu.REG_FILE._02997_ ),
    .B(\u_cpu.REG_FILE._03501_ ),
    .C(\u_cpu.REG_FILE._03512_ ),
    .Y(\u_cpu.REG_FILE._03513_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08223_  (.A1(\u_cpu.REG_FILE._03479_ ),
    .A2(\u_cpu.REG_FILE._03490_ ),
    .B1(\u_cpu.REG_FILE._03513_ ),
    .C1(\u_cpu.REG_FILE._03467_ ),
    .X(\u_cpu.ALU.SrcB[11] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08224_  (.A(\u_cpu.REG_FILE.rf[15][12] ),
    .B_N(\u_cpu.REG_FILE._02754_ ),
    .X(\u_cpu.REG_FILE._03514_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08225_  (.A1(\u_cpu.REG_FILE.rf[14][12] ),
    .A2(\u_cpu.REG_FILE._03418_ ),
    .B1(\u_cpu.REG_FILE._02752_ ),
    .C1(\u_cpu.REG_FILE._03514_ ),
    .Y(\u_cpu.REG_FILE._03515_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08226_  (.A1(\u_cpu.REG_FILE.rf[12][12] ),
    .A2(\u_cpu.REG_FILE._02760_ ),
    .B1_N(\u_cpu.REG_FILE._02761_ ),
    .X(\u_cpu.REG_FILE._03516_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08227_  (.A1(\u_cpu.REG_FILE.rf[13][12] ),
    .A2(\u_cpu.REG_FILE._02759_ ),
    .B1(\u_cpu.REG_FILE._03516_ ),
    .Y(\u_cpu.REG_FILE._03517_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08228_  (.A(\u_cpu.REG_FILE._03515_ ),
    .B(\u_cpu.REG_FILE._03517_ ),
    .C(\u_cpu.REG_FILE._02978_ ),
    .Y(\u_cpu.REG_FILE._03518_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08229_  (.A_N(\u_cpu.REG_FILE.rf[9][12] ),
    .B(\u_cpu.REG_FILE._02768_ ),
    .X(\u_cpu.REG_FILE._03519_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08230_  (.A1(\u_cpu.REG_FILE.rf[8][12] ),
    .A2(\u_cpu.REG_FILE._02772_ ),
    .B1_N(\u_cpu.REG_FILE._02774_ ),
    .Y(\u_cpu.REG_FILE._03520_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08231_  (.A(\u_cpu.REG_FILE.rf[11][12] ),
    .B_N(\u_cpu.REG_FILE._02986_ ),
    .X(\u_cpu.REG_FILE._03521_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08232_  (.A1(\u_cpu.REG_FILE.rf[10][12] ),
    .A2(\u_cpu.REG_FILE._02780_ ),
    .B1(\u_cpu.REG_FILE._02782_ ),
    .C1(\u_cpu.REG_FILE._03521_ ),
    .Y(\u_cpu.REG_FILE._03522_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08233_  (.A1(\u_cpu.REG_FILE._03519_ ),
    .A2(\u_cpu.REG_FILE._03520_ ),
    .B1(\u_cpu.REG_FILE._03062_ ),
    .C1(\u_cpu.REG_FILE._03522_ ),
    .Y(\u_cpu.REG_FILE._03523_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08234_  (.A(\u_cpu.REG_FILE._03518_ ),
    .B(\u_cpu.REG_FILE._03523_ ),
    .C(\u_cpu.REG_FILE._02788_ ),
    .Y(\u_cpu.REG_FILE._03524_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08235_  (.A1(\u_cpu.REG_FILE.rf[4][12] ),
    .A2(\u_cpu.REG_FILE._02793_ ),
    .B1_N(\u_cpu.REG_FILE._02954_ ),
    .Y(\u_cpu.REG_FILE._03525_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._08236_  (.A1(\u_cpu.REG_FILE._01798_ ),
    .A2(\u_cpu.REG_FILE._02946_ ),
    .B1(\u_cpu.REG_FILE._03525_ ),
    .Y(\u_cpu.REG_FILE._03526_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08237_  (.A1(\u_cpu.REG_FILE.rf[6][12] ),
    .A2(\u_cpu.REG_FILE._03331_ ),
    .B1(\u_cpu.REG_FILE._02799_ ),
    .Y(\u_cpu.REG_FILE._03527_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08238_  (.A_N(\u_cpu.REG_FILE.rf[7][12] ),
    .B(\u_cpu.REG_FILE._02801_ ),
    .X(\u_cpu.REG_FILE._03528_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08239_  (.A1(\u_cpu.REG_FILE._03527_ ),
    .A2(\u_cpu.REG_FILE._03528_ ),
    .B1(\u_cpu.REG_FILE._03434_ ),
    .Y(\u_cpu.REG_FILE._03529_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08240_  (.A(\u_cpu.REG_FILE._02747_ ),
    .X(\u_cpu.REG_FILE._03530_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08241_  (.A_N(\u_cpu.REG_FILE.rf[1][12] ),
    .B(\u_cpu.REG_FILE._03530_ ),
    .X(\u_cpu.REG_FILE._03531_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08242_  (.A1(\u_cpu.REG_FILE.rf[0][12] ),
    .A2(\u_cpu.REG_FILE._02811_ ),
    .B1_N(\u_cpu.REG_FILE._02812_ ),
    .Y(\u_cpu.REG_FILE._03532_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08243_  (.A(\u_cpu.REG_FILE.rf[3][12] ),
    .B_N(\u_cpu.REG_FILE._03337_ ),
    .X(\u_cpu.REG_FILE._03533_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08244_  (.A1(\u_cpu.REG_FILE.rf[2][12] ),
    .A2(\u_cpu.REG_FILE._02903_ ),
    .B1(\u_cpu.REG_FILE._02818_ ),
    .C1(\u_cpu.REG_FILE._03533_ ),
    .Y(\u_cpu.REG_FILE._03534_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08245_  (.A1(\u_cpu.REG_FILE._03531_ ),
    .A2(\u_cpu.REG_FILE._03532_ ),
    .B1(\u_cpu.REG_FILE._02814_ ),
    .C1(\u_cpu.REG_FILE._03534_ ),
    .Y(\u_cpu.REG_FILE._03535_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08246_  (.A1(\u_cpu.REG_FILE._03526_ ),
    .A2(\u_cpu.REG_FILE._03529_ ),
    .B1(\u_cpu.REG_FILE._02965_ ),
    .C1(\u_cpu.REG_FILE._03535_ ),
    .Y(\u_cpu.REG_FILE._03536_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._08247_  (.A(\u_cpu.REG_FILE._03524_ ),
    .B(\u_cpu.REG_FILE._03536_ ),
    .Y(\u_cpu.REG_FILE._03537_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08248_  (.A(\u_cpu.REG_FILE.rf[27][12] ),
    .B_N(\u_cpu.REG_FILE._02827_ ),
    .X(\u_cpu.REG_FILE._03538_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08249_  (.A1(\u_cpu.REG_FILE.rf[26][12] ),
    .A2(\u_cpu.REG_FILE._02824_ ),
    .B1(\u_cpu.REG_FILE._03000_ ),
    .C1(\u_cpu.REG_FILE._03538_ ),
    .X(\u_cpu.REG_FILE._03539_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08250_  (.A1(\u_cpu.REG_FILE.rf[24][12] ),
    .A2(\u_cpu.REG_FILE._03445_ ),
    .B1_N(\u_cpu.REG_FILE._02865_ ),
    .X(\u_cpu.REG_FILE._03540_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08251_  (.A(\u_cpu.REG_FILE.rf[25][12] ),
    .B_N(\u_cpu.REG_FILE._02832_ ),
    .X(\u_cpu.REG_FILE._03541_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._08252_  (.A1(\u_cpu.REG_FILE._03540_ ),
    .A2(\u_cpu.REG_FILE._03541_ ),
    .B1(\u_cpu.REG_FILE._02764_ ),
    .X(\u_cpu.REG_FILE._03542_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08253_  (.A(\u_cpu.REG_FILE.rf[30][12] ),
    .B(\u_cpu.REG_FILE._03063_ ),
    .Y(\u_cpu.REG_FILE._03543_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08254_  (.A1(\u_cpu.REG_FILE.rf[31][12] ),
    .A2(\u_cpu.REG_FILE._03297_ ),
    .B1(\u_cpu.REG_FILE._02854_ ),
    .Y(\u_cpu.REG_FILE._03544_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08255_  (.A(\u_cpu.REG_FILE.rf[28][12] ),
    .B(\u_cpu.REG_FILE._02916_ ),
    .Y(\u_cpu.REG_FILE._03545_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08256_  (.A1(\u_cpu.REG_FILE.rf[29][12] ),
    .A2(\u_cpu.REG_FILE._03351_ ),
    .B1_N(\u_cpu.REG_FILE._02947_ ),
    .Y(\u_cpu.REG_FILE._03546_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._08257_  (.A1(\u_cpu.REG_FILE._03543_ ),
    .A2(\u_cpu.REG_FILE._03544_ ),
    .B1(\u_cpu.REG_FILE._03545_ ),
    .B2(\u_cpu.REG_FILE._03546_ ),
    .C1(\u_cpu.REG_FILE._02919_ ),
    .Y(\u_cpu.REG_FILE._03547_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08258_  (.A1(\u_cpu.REG_FILE._03539_ ),
    .A2(\u_cpu.REG_FILE._03542_ ),
    .B1(\u_cpu.REG_FILE._02836_ ),
    .C1(\u_cpu.REG_FILE._03547_ ),
    .Y(\u_cpu.REG_FILE._03548_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08259_  (.A1(\u_cpu.REG_FILE.rf[18][12] ),
    .A2(\u_cpu.REG_FILE._02923_ ),
    .B1(\u_cpu.REG_FILE._03249_ ),
    .Y(\u_cpu.REG_FILE._03549_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08260_  (.A(\u_cpu.REG_FILE.rf[19][12] ),
    .B(\u_cpu.REG_FILE._02856_ ),
    .Y(\u_cpu.REG_FILE._03550_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08261_  (.A1(\u_cpu.REG_FILE.rf[16][12] ),
    .A2(\u_cpu.REG_FILE._03038_ ),
    .B1_N(\u_cpu.REG_FILE._02861_ ),
    .X(\u_cpu.REG_FILE._03551_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08262_  (.A1(\u_cpu.REG_FILE.rf[17][12] ),
    .A2(\u_cpu.REG_FILE._03304_ ),
    .B1(\u_cpu.REG_FILE._03551_ ),
    .Y(\u_cpu.REG_FILE._03552_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08263_  (.A1(\u_cpu.REG_FILE._03549_ ),
    .A2(\u_cpu.REG_FILE._03550_ ),
    .B1(\u_cpu.REG_FILE._03292_ ),
    .C1(\u_cpu.REG_FILE._03552_ ),
    .Y(\u_cpu.REG_FILE._03553_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._08264_  (.A(\u_cpu.REG_FILE.rf[22][12] ),
    .B(\u_cpu.REG_FILE._03143_ ),
    .X(\u_cpu.REG_FILE._03554_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08265_  (.A1(\u_cpu.REG_FILE.rf[23][12] ),
    .A2(\u_cpu.REG_FILE._03142_ ),
    .B1(\u_cpu.REG_FILE._03255_ ),
    .C1(\u_cpu.REG_FILE._03554_ ),
    .Y(\u_cpu.REG_FILE._03555_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08266_  (.A1(\u_cpu.REG_FILE.rf[20][12] ),
    .A2(\u_cpu.REG_FILE._03016_ ),
    .B1_N(\u_cpu.REG_FILE._02931_ ),
    .X(\u_cpu.REG_FILE._03556_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08267_  (.A1(\u_cpu.REG_FILE.rf[21][12] ),
    .A2(\u_cpu.REG_FILE._02870_ ),
    .B1(\u_cpu.REG_FILE._03556_ ),
    .Y(\u_cpu.REG_FILE._03557_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08268_  (.A(\u_cpu.REG_FILE._03555_ ),
    .B(\u_cpu.REG_FILE._03557_ ),
    .C(\u_cpu.REG_FILE._02875_ ),
    .Y(\u_cpu.REG_FILE._03558_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08269_  (.A(\u_cpu.REG_FILE._02922_ ),
    .B(\u_cpu.REG_FILE._03553_ ),
    .C(\u_cpu.REG_FILE._03558_ ),
    .Y(\u_cpu.REG_FILE._03559_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08270_  (.A(\u_cpu.REG_FILE._03548_ ),
    .B(\u_cpu.REG_FILE._03559_ ),
    .C(\u_cpu.REG_FILE._02878_ ),
    .Y(\u_cpu.REG_FILE._03560_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08271_  (.A1(\u_cpu.REG_FILE._02746_ ),
    .A2(\u_cpu.REG_FILE._03537_ ),
    .B1(\u_cpu.REG_FILE._03560_ ),
    .C1(\u_cpu.REG_FILE._03467_ ),
    .X(\u_cpu.ALU.SrcB[12] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08272_  (.A(\u_cpu.REG_FILE.rf[15][13] ),
    .B_N(\u_cpu.REG_FILE._02754_ ),
    .X(\u_cpu.REG_FILE._03561_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08273_  (.A1(\u_cpu.REG_FILE.rf[14][13] ),
    .A2(\u_cpu.REG_FILE._03418_ ),
    .B1(\u_cpu.REG_FILE._02752_ ),
    .C1(\u_cpu.REG_FILE._03561_ ),
    .Y(\u_cpu.REG_FILE._03562_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08274_  (.A1(\u_cpu.REG_FILE.rf[12][13] ),
    .A2(\u_cpu.REG_FILE._02760_ ),
    .B1_N(\u_cpu.REG_FILE._02761_ ),
    .X(\u_cpu.REG_FILE._03563_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08275_  (.A1(\u_cpu.REG_FILE.rf[13][13] ),
    .A2(\u_cpu.REG_FILE._02759_ ),
    .B1(\u_cpu.REG_FILE._03563_ ),
    .Y(\u_cpu.REG_FILE._03564_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08276_  (.A(\u_cpu.REG_FILE._03562_ ),
    .B(\u_cpu.REG_FILE._03564_ ),
    .C(\u_cpu.REG_FILE._02978_ ),
    .Y(\u_cpu.REG_FILE._03565_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08277_  (.A_N(\u_cpu.REG_FILE.rf[9][13] ),
    .B(\u_cpu.REG_FILE._02945_ ),
    .X(\u_cpu.REG_FILE._03566_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08278_  (.A1(\u_cpu.REG_FILE.rf[8][13] ),
    .A2(\u_cpu.REG_FILE._02816_ ),
    .B1_N(\u_cpu.REG_FILE._02774_ ),
    .Y(\u_cpu.REG_FILE._03567_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08279_  (.A(\u_cpu.REG_FILE.rf[11][13] ),
    .B_N(\u_cpu.REG_FILE._02986_ ),
    .X(\u_cpu.REG_FILE._03568_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08280_  (.A1(\u_cpu.REG_FILE.rf[10][13] ),
    .A2(\u_cpu.REG_FILE._02780_ ),
    .B1(\u_cpu.REG_FILE._02782_ ),
    .C1(\u_cpu.REG_FILE._03568_ ),
    .Y(\u_cpu.REG_FILE._03569_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08281_  (.A1(\u_cpu.REG_FILE._03566_ ),
    .A2(\u_cpu.REG_FILE._03567_ ),
    .B1(\u_cpu.REG_FILE._03062_ ),
    .C1(\u_cpu.REG_FILE._03569_ ),
    .Y(\u_cpu.REG_FILE._03570_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08282_  (.A(\u_cpu.REG_FILE._03565_ ),
    .B(\u_cpu.REG_FILE._03570_ ),
    .C(\u_cpu.REG_FILE._02788_ ),
    .Y(\u_cpu.REG_FILE._03571_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08283_  (.A1(\u_cpu.REG_FILE.rf[4][13] ),
    .A2(\u_cpu.REG_FILE._02793_ ),
    .B1_N(\u_cpu.REG_FILE._02954_ ),
    .Y(\u_cpu.REG_FILE._03572_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._08284_  (.A1(\u_cpu.REG_FILE._01849_ ),
    .A2(\u_cpu.REG_FILE._02946_ ),
    .B1(\u_cpu.REG_FILE._03572_ ),
    .Y(\u_cpu.REG_FILE._03573_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08285_  (.A1(\u_cpu.REG_FILE.rf[6][13] ),
    .A2(\u_cpu.REG_FILE._03331_ ),
    .B1(\u_cpu.REG_FILE._03407_ ),
    .Y(\u_cpu.REG_FILE._03574_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08286_  (.A_N(\u_cpu.REG_FILE.rf[7][13] ),
    .B(\u_cpu.REG_FILE._02801_ ),
    .X(\u_cpu.REG_FILE._03575_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08287_  (.A1(\u_cpu.REG_FILE._03574_ ),
    .A2(\u_cpu.REG_FILE._03575_ ),
    .B1(\u_cpu.REG_FILE._03434_ ),
    .Y(\u_cpu.REG_FILE._03576_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08288_  (.A_N(\u_cpu.REG_FILE.rf[1][13] ),
    .B(\u_cpu.REG_FILE._03530_ ),
    .X(\u_cpu.REG_FILE._03577_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08289_  (.A1(\u_cpu.REG_FILE.rf[0][13] ),
    .A2(\u_cpu.REG_FILE._02811_ ),
    .B1_N(\u_cpu.REG_FILE._02812_ ),
    .Y(\u_cpu.REG_FILE._03578_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08290_  (.A(\u_cpu.REG_FILE.rf[3][13] ),
    .B_N(\u_cpu.REG_FILE._03337_ ),
    .X(\u_cpu.REG_FILE._03579_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08291_  (.A1(\u_cpu.REG_FILE.rf[2][13] ),
    .A2(\u_cpu.REG_FILE._02903_ ),
    .B1(\u_cpu.REG_FILE._03026_ ),
    .C1(\u_cpu.REG_FILE._03579_ ),
    .Y(\u_cpu.REG_FILE._03580_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08292_  (.A1(\u_cpu.REG_FILE._03577_ ),
    .A2(\u_cpu.REG_FILE._03578_ ),
    .B1(\u_cpu.REG_FILE._02814_ ),
    .C1(\u_cpu.REG_FILE._03580_ ),
    .Y(\u_cpu.REG_FILE._03581_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08293_  (.A1(\u_cpu.REG_FILE._03573_ ),
    .A2(\u_cpu.REG_FILE._03576_ ),
    .B1(\u_cpu.REG_FILE._02965_ ),
    .C1(\u_cpu.REG_FILE._03581_ ),
    .Y(\u_cpu.REG_FILE._03582_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._08294_  (.A(\u_cpu.REG_FILE._03571_ ),
    .B(\u_cpu.REG_FILE._03582_ ),
    .Y(\u_cpu.REG_FILE._03583_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08295_  (.A(\u_cpu.REG_FILE.rf[27][13] ),
    .B_N(\u_cpu.REG_FILE._02827_ ),
    .X(\u_cpu.REG_FILE._03584_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08296_  (.A1(\u_cpu.REG_FILE.rf[26][13] ),
    .A2(\u_cpu.REG_FILE._02824_ ),
    .B1(\u_cpu.REG_FILE._03000_ ),
    .C1(\u_cpu.REG_FILE._03584_ ),
    .X(\u_cpu.REG_FILE._03585_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08297_  (.A1(\u_cpu.REG_FILE.rf[24][13] ),
    .A2(\u_cpu.REG_FILE._03445_ ),
    .B1_N(\u_cpu.REG_FILE._02865_ ),
    .X(\u_cpu.REG_FILE._03586_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08298_  (.A(\u_cpu.REG_FILE.rf[25][13] ),
    .B_N(\u_cpu.REG_FILE._02832_ ),
    .X(\u_cpu.REG_FILE._03587_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._08299_  (.A1(\u_cpu.REG_FILE._03586_ ),
    .A2(\u_cpu.REG_FILE._03587_ ),
    .B1(\u_cpu.REG_FILE._02764_ ),
    .X(\u_cpu.REG_FILE._03588_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08300_  (.A1(\u_cpu.REG_FILE.rf[28][13] ),
    .A2(\u_cpu.REG_FILE._02837_ ),
    .B1_N(\u_cpu.REG_FILE._03201_ ),
    .Y(\u_cpu.REG_FILE._03589_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08301_  (.A(\u_cpu.REG_FILE.rf[29][13] ),
    .B(\u_cpu.REG_FILE._02841_ ),
    .Y(\u_cpu.REG_FILE._03590_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08302_  (.A(\u_cpu.REG_FILE.rf[30][13] ),
    .B(\u_cpu.REG_FILE._02916_ ),
    .Y(\u_cpu.REG_FILE._03591_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08303_  (.A1(\u_cpu.REG_FILE.rf[31][13] ),
    .A2(\u_cpu.REG_FILE._02845_ ),
    .B1(\u_cpu.REG_FILE._02846_ ),
    .Y(\u_cpu.REG_FILE._03592_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._08304_  (.A1(\u_cpu.REG_FILE._03589_ ),
    .A2(\u_cpu.REG_FILE._03590_ ),
    .B1(\u_cpu.REG_FILE._03591_ ),
    .B2(\u_cpu.REG_FILE._03592_ ),
    .C1(\u_cpu.REG_FILE._02919_ ),
    .Y(\u_cpu.REG_FILE._03593_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08305_  (.A1(\u_cpu.REG_FILE._03585_ ),
    .A2(\u_cpu.REG_FILE._03588_ ),
    .B1(\u_cpu.REG_FILE._02836_ ),
    .C1(\u_cpu.REG_FILE._03593_ ),
    .Y(\u_cpu.REG_FILE._03594_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08306_  (.A1(\u_cpu.REG_FILE.rf[18][13] ),
    .A2(\u_cpu.REG_FILE._02923_ ),
    .B1(\u_cpu.REG_FILE._03249_ ),
    .Y(\u_cpu.REG_FILE._03595_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08307_  (.A(\u_cpu.REG_FILE.rf[19][13] ),
    .B(\u_cpu.REG_FILE._02856_ ),
    .Y(\u_cpu.REG_FILE._03596_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08308_  (.A1(\u_cpu.REG_FILE.rf[16][13] ),
    .A2(\u_cpu.REG_FILE._03038_ ),
    .B1_N(\u_cpu.REG_FILE._02861_ ),
    .X(\u_cpu.REG_FILE._03597_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08309_  (.A1(\u_cpu.REG_FILE.rf[17][13] ),
    .A2(\u_cpu.REG_FILE._03304_ ),
    .B1(\u_cpu.REG_FILE._03597_ ),
    .Y(\u_cpu.REG_FILE._03598_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08310_  (.A1(\u_cpu.REG_FILE._03595_ ),
    .A2(\u_cpu.REG_FILE._03596_ ),
    .B1(\u_cpu.REG_FILE._03292_ ),
    .C1(\u_cpu.REG_FILE._03598_ ),
    .Y(\u_cpu.REG_FILE._03599_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._08311_  (.A(\u_cpu.REG_FILE.rf[22][13] ),
    .B(\u_cpu.REG_FILE._03143_ ),
    .X(\u_cpu.REG_FILE._03600_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08312_  (.A1(\u_cpu.REG_FILE.rf[23][13] ),
    .A2(\u_cpu.REG_FILE._03142_ ),
    .B1(\u_cpu.REG_FILE._03255_ ),
    .C1(\u_cpu.REG_FILE._03600_ ),
    .Y(\u_cpu.REG_FILE._03601_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08313_  (.A1(\u_cpu.REG_FILE.rf[20][13] ),
    .A2(\u_cpu.REG_FILE._03016_ ),
    .B1_N(\u_cpu.REG_FILE._02931_ ),
    .X(\u_cpu.REG_FILE._03602_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08314_  (.A1(\u_cpu.REG_FILE.rf[21][13] ),
    .A2(\u_cpu.REG_FILE._02870_ ),
    .B1(\u_cpu.REG_FILE._03602_ ),
    .Y(\u_cpu.REG_FILE._03603_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08315_  (.A(\u_cpu.REG_FILE._03601_ ),
    .B(\u_cpu.REG_FILE._03603_ ),
    .C(\u_cpu.REG_FILE._02875_ ),
    .Y(\u_cpu.REG_FILE._03604_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08316_  (.A(\u_cpu.REG_FILE._02922_ ),
    .B(\u_cpu.REG_FILE._03599_ ),
    .C(\u_cpu.REG_FILE._03604_ ),
    .Y(\u_cpu.REG_FILE._03605_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08317_  (.A(\u_cpu.REG_FILE._03594_ ),
    .B(\u_cpu.REG_FILE._03605_ ),
    .C(\u_cpu.REG_FILE._02878_ ),
    .Y(\u_cpu.REG_FILE._03606_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08318_  (.A1(\u_cpu.REG_FILE._02746_ ),
    .A2(\u_cpu.REG_FILE._03583_ ),
    .B1(\u_cpu.REG_FILE._03606_ ),
    .C1(\u_cpu.REG_FILE._03467_ ),
    .X(\u_cpu.ALU.SrcB[13] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08319_  (.A(\u_cpu.REG_FILE.rf[15][14] ),
    .B_N(\u_cpu.REG_FILE._02754_ ),
    .X(\u_cpu.REG_FILE._03607_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08320_  (.A1(\u_cpu.REG_FILE.rf[14][14] ),
    .A2(\u_cpu.REG_FILE._03418_ ),
    .B1(\u_cpu.REG_FILE._02752_ ),
    .C1(\u_cpu.REG_FILE._03607_ ),
    .Y(\u_cpu.REG_FILE._03608_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08321_  (.A1(\u_cpu.REG_FILE.rf[12][14] ),
    .A2(\u_cpu.REG_FILE._02974_ ),
    .B1_N(\u_cpu.REG_FILE._02761_ ),
    .X(\u_cpu.REG_FILE._03609_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08322_  (.A1(\u_cpu.REG_FILE.rf[13][14] ),
    .A2(\u_cpu.REG_FILE._02759_ ),
    .B1(\u_cpu.REG_FILE._03609_ ),
    .Y(\u_cpu.REG_FILE._03610_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08323_  (.A(\u_cpu.REG_FILE._03608_ ),
    .B(\u_cpu.REG_FILE._03610_ ),
    .C(\u_cpu.REG_FILE._02978_ ),
    .Y(\u_cpu.REG_FILE._03611_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08324_  (.A_N(\u_cpu.REG_FILE.rf[9][14] ),
    .B(\u_cpu.REG_FILE._02945_ ),
    .X(\u_cpu.REG_FILE._03612_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08325_  (.A1(\u_cpu.REG_FILE.rf[8][14] ),
    .A2(\u_cpu.REG_FILE._02816_ ),
    .B1_N(\u_cpu.REG_FILE._02947_ ),
    .Y(\u_cpu.REG_FILE._03613_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08326_  (.A(\u_cpu.REG_FILE.rf[11][14] ),
    .B_N(\u_cpu.REG_FILE._02986_ ),
    .X(\u_cpu.REG_FILE._03614_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08327_  (.A1(\u_cpu.REG_FILE.rf[10][14] ),
    .A2(\u_cpu.REG_FILE._02780_ ),
    .B1(\u_cpu.REG_FILE._02846_ ),
    .C1(\u_cpu.REG_FILE._03614_ ),
    .Y(\u_cpu.REG_FILE._03615_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08328_  (.A1(\u_cpu.REG_FILE._03612_ ),
    .A2(\u_cpu.REG_FILE._03613_ ),
    .B1(\u_cpu.REG_FILE._03062_ ),
    .C1(\u_cpu.REG_FILE._03615_ ),
    .Y(\u_cpu.REG_FILE._03616_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08329_  (.A(\u_cpu.REG_FILE._03611_ ),
    .B(\u_cpu.REG_FILE._03616_ ),
    .C(\u_cpu.REG_FILE._03218_ ),
    .Y(\u_cpu.REG_FILE._03617_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08330_  (.A1(\u_cpu.REG_FILE.rf[4][14] ),
    .A2(\u_cpu.REG_FILE._02793_ ),
    .B1_N(\u_cpu.REG_FILE._02954_ ),
    .Y(\u_cpu.REG_FILE._03618_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._08331_  (.A1(\u_cpu.REG_FILE._01902_ ),
    .A2(\u_cpu.REG_FILE._02946_ ),
    .B1(\u_cpu.REG_FILE._03618_ ),
    .Y(\u_cpu.REG_FILE._03619_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08332_  (.A1(\u_cpu.REG_FILE.rf[6][14] ),
    .A2(\u_cpu.REG_FILE._03331_ ),
    .B1(\u_cpu.REG_FILE._03407_ ),
    .Y(\u_cpu.REG_FILE._03620_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08333_  (.A_N(\u_cpu.REG_FILE.rf[7][14] ),
    .B(\u_cpu.REG_FILE._02808_ ),
    .X(\u_cpu.REG_FILE._03621_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08334_  (.A1(\u_cpu.REG_FILE._03620_ ),
    .A2(\u_cpu.REG_FILE._03621_ ),
    .B1(\u_cpu.REG_FILE._03434_ ),
    .Y(\u_cpu.REG_FILE._03622_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08335_  (.A_N(\u_cpu.REG_FILE.rf[1][14] ),
    .B(\u_cpu.REG_FILE._03530_ ),
    .X(\u_cpu.REG_FILE._03623_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08336_  (.A1(\u_cpu.REG_FILE.rf[0][14] ),
    .A2(\u_cpu.REG_FILE._02811_ ),
    .B1_N(\u_cpu.REG_FILE._02794_ ),
    .Y(\u_cpu.REG_FILE._03624_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08337_  (.A(\u_cpu.REG_FILE.rf[3][14] ),
    .B_N(\u_cpu.REG_FILE._03337_ ),
    .X(\u_cpu.REG_FILE._03625_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08338_  (.A1(\u_cpu.REG_FILE.rf[2][14] ),
    .A2(\u_cpu.REG_FILE._02903_ ),
    .B1(\u_cpu.REG_FILE._03026_ ),
    .C1(\u_cpu.REG_FILE._03625_ ),
    .Y(\u_cpu.REG_FILE._03626_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08339_  (.A1(\u_cpu.REG_FILE._03623_ ),
    .A2(\u_cpu.REG_FILE._03624_ ),
    .B1(\u_cpu.REG_FILE._02858_ ),
    .C1(\u_cpu.REG_FILE._03626_ ),
    .Y(\u_cpu.REG_FILE._03627_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08340_  (.A1(\u_cpu.REG_FILE._03619_ ),
    .A2(\u_cpu.REG_FILE._03622_ ),
    .B1(\u_cpu.REG_FILE._02965_ ),
    .C1(\u_cpu.REG_FILE._03627_ ),
    .Y(\u_cpu.REG_FILE._03628_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._08341_  (.A(\u_cpu.REG_FILE._03617_ ),
    .B(\u_cpu.REG_FILE._03628_ ),
    .Y(\u_cpu.REG_FILE._03629_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08342_  (.A(\u_cpu.REG_FILE.rf[27][14] ),
    .B_N(\u_cpu.REG_FILE._02771_ ),
    .X(\u_cpu.REG_FILE._03630_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08343_  (.A1(\u_cpu.REG_FILE.rf[26][14] ),
    .A2(\u_cpu.REG_FILE._03287_ ),
    .B1(\u_cpu.REG_FILE._02854_ ),
    .C1(\u_cpu.REG_FILE._03630_ ),
    .X(\u_cpu.REG_FILE._03631_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08344_  (.A1(\u_cpu.REG_FILE.rf[24][14] ),
    .A2(\u_cpu.REG_FILE._03204_ ),
    .B1_N(\u_cpu.REG_FILE._03201_ ),
    .Y(\u_cpu.REG_FILE._03632_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08345_  (.A_N(\u_cpu.REG_FILE.rf[25][14] ),
    .B(\u_cpu.REG_FILE._02880_ ),
    .X(\u_cpu.REG_FILE._03633_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08346_  (.A1(\u_cpu.REG_FILE._03632_ ),
    .A2(\u_cpu.REG_FILE._03633_ ),
    .B1(\u_cpu.REG_FILE._03292_ ),
    .Y(\u_cpu.REG_FILE._03634_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08347_  (.A1(\u_cpu.REG_FILE.rf[28][14] ),
    .A2(\u_cpu.REG_FILE._02790_ ),
    .B1_N(\u_cpu.REG_FILE._02751_ ),
    .Y(\u_cpu.REG_FILE._03635_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08348_  (.A_N(\u_cpu.REG_FILE.rf[29][14] ),
    .B(\u_cpu.REG_FILE._02754_ ),
    .X(\u_cpu.REG_FILE._03636_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08349_  (.A(\u_cpu.REG_FILE.rf[30][14] ),
    .B(\u_cpu.REG_FILE._03071_ ),
    .Y(\u_cpu.REG_FILE._03637_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08350_  (.A1(\u_cpu.REG_FILE.rf[31][14] ),
    .A2(\u_cpu.REG_FILE._03297_ ),
    .B1(\u_cpu.REG_FILE._03064_ ),
    .Y(\u_cpu.REG_FILE._03638_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.REG_FILE._08351_  (.A1(\u_cpu.REG_FILE._03635_ ),
    .A2(\u_cpu.REG_FILE._03636_ ),
    .B1(\u_cpu.REG_FILE._03637_ ),
    .B2(\u_cpu.REG_FILE._03638_ ),
    .Y(\u_cpu.REG_FILE._03639_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._08352_  (.A1(\u_cpu.REG_FILE._03631_ ),
    .A2(\u_cpu.REG_FILE._03634_ ),
    .B1(\u_cpu.REG_FILE._03024_ ),
    .B2(\u_cpu.REG_FILE._03639_ ),
    .C1(\u_cpu.REG_FILE._03218_ ),
    .Y(\u_cpu.REG_FILE._03640_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08353_  (.A1(\u_cpu.REG_FILE.rf[18][14] ),
    .A2(\u_cpu.REG_FILE._02923_ ),
    .B1(\u_cpu.REG_FILE._03249_ ),
    .Y(\u_cpu.REG_FILE._03641_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08354_  (.A(\u_cpu.REG_FILE.rf[19][14] ),
    .B(\u_cpu.REG_FILE._02856_ ),
    .Y(\u_cpu.REG_FILE._03642_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08355_  (.A1(\u_cpu.REG_FILE.rf[16][14] ),
    .A2(\u_cpu.REG_FILE._03038_ ),
    .B1_N(\u_cpu.REG_FILE._02861_ ),
    .X(\u_cpu.REG_FILE._03643_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08356_  (.A1(\u_cpu.REG_FILE.rf[17][14] ),
    .A2(\u_cpu.REG_FILE._03304_ ),
    .B1(\u_cpu.REG_FILE._03643_ ),
    .Y(\u_cpu.REG_FILE._03644_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08357_  (.A1(\u_cpu.REG_FILE._03641_ ),
    .A2(\u_cpu.REG_FILE._03642_ ),
    .B1(\u_cpu.REG_FILE._03292_ ),
    .C1(\u_cpu.REG_FILE._03644_ ),
    .Y(\u_cpu.REG_FILE._03645_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08358_  (.A(\u_cpu.REG_FILE.rf[20][14] ),
    .B(\u_cpu.REG_FILE._03309_ ),
    .Y(\u_cpu.REG_FILE._03646_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08359_  (.A_N(\u_cpu.REG_FILE.rf[21][14] ),
    .B(\u_cpu.REG_FILE._03311_ ),
    .X(\u_cpu.REG_FILE._03647_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08360_  (.A(\u_cpu.REG_FILE.rf[23][14] ),
    .B_N(\u_cpu.REG_FILE._02852_ ),
    .X(\u_cpu.REG_FILE._03648_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08361_  (.A1(\u_cpu.REG_FILE.rf[22][14] ),
    .A2(\u_cpu.REG_FILE._02797_ ),
    .B1(\u_cpu.REG_FILE._03198_ ),
    .C1(\u_cpu.REG_FILE._03648_ ),
    .Y(\u_cpu.REG_FILE._03649_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._08362_  (.A1(\u_cpu.REG_FILE._03308_ ),
    .A2(\u_cpu.REG_FILE._03646_ ),
    .A3(\u_cpu.REG_FILE._03647_ ),
    .B1(\u_cpu.REG_FILE._02834_ ),
    .C1(\u_cpu.REG_FILE._03649_ ),
    .Y(\u_cpu.REG_FILE._03650_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08363_  (.A(\u_cpu.REG_FILE._02922_ ),
    .B(\u_cpu.REG_FILE._03645_ ),
    .C(\u_cpu.REG_FILE._03650_ ),
    .Y(\u_cpu.REG_FILE._03651_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08364_  (.A(\u_cpu.REG_FILE._03640_ ),
    .B(\u_cpu.REG_FILE._03651_ ),
    .C(\u_cpu.REG_FILE._02745_ ),
    .Y(\u_cpu.REG_FILE._03652_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08365_  (.A1(\u_cpu.REG_FILE._02746_ ),
    .A2(\u_cpu.REG_FILE._03629_ ),
    .B1(\u_cpu.REG_FILE._03652_ ),
    .C1(\u_cpu.REG_FILE._03467_ ),
    .X(\u_cpu.ALU.SrcB[14] ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08366_  (.A(\u_cpu.REG_FILE._02810_ ),
    .X(\u_cpu.REG_FILE._03653_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08367_  (.A1(\u_cpu.REG_FILE.rf[18][15] ),
    .A2(\u_cpu.REG_FILE._03653_ ),
    .B1(\u_cpu.REG_FILE._02941_ ),
    .Y(\u_cpu.REG_FILE._03654_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._08368_  (.A1(\u_cpu.REG_FILE._01975_ ),
    .A2(\u_cpu.REG_FILE._02939_ ),
    .B1(\u_cpu.REG_FILE._03654_ ),
    .Y(\u_cpu.REG_FILE._03655_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08369_  (.A(\u_cpu.REG_FILE.rf[16][15] ),
    .B(\u_cpu.REG_FILE._03371_ ),
    .Y(\u_cpu.REG_FILE._03656_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._08370_  (.A1(\u_cpu.REG_FILE._01978_ ),
    .A2(\u_cpu.REG_FILE._03166_ ),
    .B1(\u_cpu.REG_FILE._02948_ ),
    .C1(\u_cpu.REG_FILE._03656_ ),
    .Y(\u_cpu.REG_FILE._03657_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08371_  (.A1(\u_cpu.REG_FILE.rf[20][15] ),
    .A2(\u_cpu.REG_FILE._02953_ ),
    .B1_N(\u_cpu.REG_FILE._03050_ ),
    .Y(\u_cpu.REG_FILE._03658_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08372_  (.A(\u_cpu.REG_FILE.rf[21][15] ),
    .B(\u_cpu.REG_FILE._02956_ ),
    .Y(\u_cpu.REG_FILE._03659_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08373_  (.A(\u_cpu.REG_FILE.rf[22][15] ),
    .B(\u_cpu.REG_FILE._02958_ ),
    .Y(\u_cpu.REG_FILE._03660_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08374_  (.A1(\u_cpu.REG_FILE.rf[23][15] ),
    .A2(\u_cpu.REG_FILE._03114_ ),
    .B1(\u_cpu.REG_FILE._03377_ ),
    .Y(\u_cpu.REG_FILE._03661_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._08375_  (.A1(\u_cpu.REG_FILE._03658_ ),
    .A2(\u_cpu.REG_FILE._03659_ ),
    .B1(\u_cpu.REG_FILE._03660_ ),
    .B2(\u_cpu.REG_FILE._03661_ ),
    .C1(\u_cpu.REG_FILE._02848_ ),
    .Y(\u_cpu.REG_FILE._03662_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.REG_FILE._08376_  (.A1(\u_cpu.REG_FILE._02937_ ),
    .A2(\u_cpu.REG_FILE._03655_ ),
    .A3(\u_cpu.REG_FILE._03657_ ),
    .B1(\u_cpu.REG_FILE._03662_ ),
    .C1(\u_cpu.REG_FILE._02966_ ),
    .X(\u_cpu.REG_FILE._03663_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08377_  (.A(\u_cpu.REG_FILE.rf[31][15] ),
    .B_N(\u_cpu.REG_FILE._02970_ ),
    .X(\u_cpu.REG_FILE._03664_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08378_  (.A1(\u_cpu.REG_FILE.rf[30][15] ),
    .A2(\u_cpu.REG_FILE._02749_ ),
    .B1(\u_cpu.REG_FILE._02969_ ),
    .C1(\u_cpu.REG_FILE._03664_ ),
    .Y(\u_cpu.REG_FILE._03665_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08379_  (.A1(\u_cpu.REG_FILE.rf[28][15] ),
    .A2(\u_cpu.REG_FILE._02974_ ),
    .B1_N(\u_cpu.REG_FILE._02975_ ),
    .X(\u_cpu.REG_FILE._03666_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08380_  (.A1(\u_cpu.REG_FILE.rf[29][15] ),
    .A2(\u_cpu.REG_FILE._02973_ ),
    .B1(\u_cpu.REG_FILE._03666_ ),
    .Y(\u_cpu.REG_FILE._03667_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08381_  (.A(\u_cpu.REG_FILE._03665_ ),
    .B(\u_cpu.REG_FILE._03667_ ),
    .C(\u_cpu.REG_FILE._03006_ ),
    .Y(\u_cpu.REG_FILE._03668_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08382_  (.A_N(\u_cpu.REG_FILE.rf[25][15] ),
    .B(\u_cpu.REG_FILE._02980_ ),
    .X(\u_cpu.REG_FILE._03669_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08383_  (.A1(\u_cpu.REG_FILE.rf[24][15] ),
    .A2(\u_cpu.REG_FILE._02982_ ),
    .B1_N(\u_cpu.REG_FILE._02983_ ),
    .Y(\u_cpu.REG_FILE._03670_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08384_  (.A(\u_cpu.REG_FILE.rf[27][15] ),
    .B_N(\u_cpu.REG_FILE._03077_ ),
    .X(\u_cpu.REG_FILE._03671_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08385_  (.A1(\u_cpu.REG_FILE.rf[26][15] ),
    .A2(\u_cpu.REG_FILE._03125_ ),
    .B1(\u_cpu.REG_FILE._02988_ ),
    .C1(\u_cpu.REG_FILE._03671_ ),
    .Y(\u_cpu.REG_FILE._03672_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08386_  (.A1(\u_cpu.REG_FILE._03669_ ),
    .A2(\u_cpu.REG_FILE._03670_ ),
    .B1(\u_cpu.REG_FILE._02985_ ),
    .C1(\u_cpu.REG_FILE._03672_ ),
    .Y(\u_cpu.REG_FILE._03673_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._08387_  (.A1(\u_cpu.REG_FILE._03668_ ),
    .A2(\u_cpu.REG_FILE._03673_ ),
    .A3(\u_cpu.REG_FILE._03129_ ),
    .B1(\u_cpu.REG_FILE._03081_ ),
    .X(\u_cpu.REG_FILE._03674_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08388_  (.A(\u_cpu.REG_FILE.rf[8][15] ),
    .B(\u_cpu.REG_FILE._02998_ ),
    .Y(\u_cpu.REG_FILE._03675_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08389_  (.A1(\u_cpu.REG_FILE.rf[9][15] ),
    .A2(\u_cpu.REG_FILE._03132_ ),
    .B1_N(\u_cpu.REG_FILE._03133_ ),
    .Y(\u_cpu.REG_FILE._03676_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._08390_  (.A(\u_cpu.REG_FILE.rf[10][15] ),
    .B(\u_cpu.REG_FILE._02867_ ),
    .X(\u_cpu.REG_FILE._03677_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08391_  (.A1(\u_cpu.REG_FILE.rf[11][15] ),
    .A2(\u_cpu.REG_FILE._03136_ ),
    .B1(\u_cpu.REG_FILE._03137_ ),
    .C1(\u_cpu.REG_FILE._03677_ ),
    .Y(\u_cpu.REG_FILE._03678_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08392_  (.A1(\u_cpu.REG_FILE._03675_ ),
    .A2(\u_cpu.REG_FILE._03676_ ),
    .B1(\u_cpu.REG_FILE._03135_ ),
    .C1(\u_cpu.REG_FILE._03678_ ),
    .Y(\u_cpu.REG_FILE._03679_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._08393_  (.A(\u_cpu.REG_FILE.rf[14][15] ),
    .B(\u_cpu.REG_FILE._03143_ ),
    .X(\u_cpu.REG_FILE._03680_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08394_  (.A1(\u_cpu.REG_FILE.rf[15][15] ),
    .A2(\u_cpu.REG_FILE._03142_ ),
    .B1(\u_cpu.REG_FILE._03255_ ),
    .C1(\u_cpu.REG_FILE._03680_ ),
    .Y(\u_cpu.REG_FILE._03681_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08395_  (.A1(\u_cpu.REG_FILE.rf[12][15] ),
    .A2(\u_cpu.REG_FILE._03016_ ),
    .B1_N(\u_cpu.REG_FILE._02931_ ),
    .X(\u_cpu.REG_FILE._03682_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08396_  (.A1(\u_cpu.REG_FILE.rf[13][15] ),
    .A2(\u_cpu.REG_FILE._02870_ ),
    .B1(\u_cpu.REG_FILE._03682_ ),
    .Y(\u_cpu.REG_FILE._03683_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08397_  (.A(\u_cpu.REG_FILE._03681_ ),
    .B(\u_cpu.REG_FILE._03683_ ),
    .C(\u_cpu.REG_FILE._03074_ ),
    .Y(\u_cpu.REG_FILE._03684_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08398_  (.A(\u_cpu.REG_FILE._03679_ ),
    .B(\u_cpu.REG_FILE._03141_ ),
    .C(\u_cpu.REG_FILE._03684_ ),
    .Y(\u_cpu.REG_FILE._03685_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08399_  (.A(\u_cpu.REG_FILE.rf[3][15] ),
    .B_N(\u_cpu.REG_FILE._02815_ ),
    .X(\u_cpu.REG_FILE._03686_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08400_  (.A1(\u_cpu.REG_FILE.rf[2][15] ),
    .A2(\u_cpu.REG_FILE._03025_ ),
    .B1(\u_cpu.REG_FILE._03026_ ),
    .C1(\u_cpu.REG_FILE._03686_ ),
    .Y(\u_cpu.REG_FILE._03687_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08401_  (.A1(\u_cpu.REG_FILE.rf[0][15] ),
    .A2(\u_cpu.REG_FILE._03030_ ),
    .B1_N(\u_cpu.REG_FILE._02872_ ),
    .X(\u_cpu.REG_FILE._03688_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08402_  (.A1(\u_cpu.REG_FILE.rf[1][15] ),
    .A2(\u_cpu.REG_FILE._03029_ ),
    .B1(\u_cpu.REG_FILE._03688_ ),
    .Y(\u_cpu.REG_FILE._03689_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08403_  (.A(\u_cpu.REG_FILE._03009_ ),
    .B(\u_cpu.REG_FILE._03687_ ),
    .C(\u_cpu.REG_FILE._03689_ ),
    .Y(\u_cpu.REG_FILE._03690_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08404_  (.A(\u_cpu.REG_FILE.rf[7][15] ),
    .B_N(\u_cpu.REG_FILE._02783_ ),
    .X(\u_cpu.REG_FILE._03691_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08405_  (.A1(\u_cpu.REG_FILE.rf[6][15] ),
    .A2(\u_cpu.REG_FILE._02843_ ),
    .B1(\u_cpu.REG_FILE._02866_ ),
    .C1(\u_cpu.REG_FILE._03691_ ),
    .Y(\u_cpu.REG_FILE._03692_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08406_  (.A1(\u_cpu.REG_FILE.rf[4][15] ),
    .A2(\u_cpu.REG_FILE._03030_ ),
    .B1_N(\u_cpu.REG_FILE._03039_ ),
    .X(\u_cpu.REG_FILE._03693_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08407_  (.A1(\u_cpu.REG_FILE.rf[5][15] ),
    .A2(\u_cpu.REG_FILE._03037_ ),
    .B1(\u_cpu.REG_FILE._03693_ ),
    .Y(\u_cpu.REG_FILE._03694_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08408_  (.A(\u_cpu.REG_FILE._03692_ ),
    .B(\u_cpu.REG_FILE._03694_ ),
    .C(\u_cpu.REG_FILE._03042_ ),
    .Y(\u_cpu.REG_FILE._03695_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08409_  (.A(\u_cpu.REG_FILE._02851_ ),
    .B(\u_cpu.REG_FILE._03690_ ),
    .C(\u_cpu.REG_FILE._03695_ ),
    .Y(\u_cpu.REG_FILE._03696_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08410_  (.A(\u_cpu.REG_FILE._02997_ ),
    .B(\u_cpu.REG_FILE._03685_ ),
    .C(\u_cpu.REG_FILE._03696_ ),
    .Y(\u_cpu.REG_FILE._03697_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08411_  (.A1(\u_cpu.REG_FILE._03663_ ),
    .A2(\u_cpu.REG_FILE._03674_ ),
    .B1(\u_cpu.REG_FILE._03697_ ),
    .C1(\u_cpu.REG_FILE._03467_ ),
    .X(\u_cpu.ALU.SrcB[15] ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08412_  (.A1(\u_cpu.REG_FILE.rf[16][16] ),
    .A2(\u_cpu.REG_FILE._02790_ ),
    .B1_N(\u_cpu.REG_FILE._02751_ ),
    .Y(\u_cpu.REG_FILE._03698_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08413_  (.A_N(\u_cpu.REG_FILE.rf[17][16] ),
    .B(\u_cpu.REG_FILE._03445_ ),
    .X(\u_cpu.REG_FILE._03699_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08414_  (.A1(\u_cpu.REG_FILE.rf[18][16] ),
    .A2(\u_cpu.REG_FILE._03404_ ),
    .B1(\u_cpu.REG_FILE._03470_ ),
    .Y(\u_cpu.REG_FILE._03700_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08415_  (.A_N(\u_cpu.REG_FILE.rf[19][16] ),
    .B(\u_cpu.REG_FILE._02980_ ),
    .X(\u_cpu.REG_FILE._03701_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.REG_FILE._08416_  (.A1(\u_cpu.REG_FILE._03698_ ),
    .A2(\u_cpu.REG_FILE._03699_ ),
    .B1(\u_cpu.REG_FILE._03700_ ),
    .B2(\u_cpu.REG_FILE._03701_ ),
    .Y(\u_cpu.REG_FILE._03702_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08417_  (.A(\u_cpu.REG_FILE.rf[23][16] ),
    .B_N(\u_cpu.REG_FILE._03003_ ),
    .X(\u_cpu.REG_FILE._03703_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08418_  (.A1(\u_cpu.REG_FILE.rf[22][16] ),
    .A2(\u_cpu.REG_FILE._02987_ ),
    .B1(\u_cpu.REG_FILE._02826_ ),
    .C1(\u_cpu.REG_FILE._03703_ ),
    .X(\u_cpu.REG_FILE._03704_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08419_  (.A(\u_cpu.REG_FILE.rf[20][16] ),
    .B(\u_cpu.REG_FILE._02940_ ),
    .Y(\u_cpu.REG_FILE._03705_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08420_  (.A_N(\u_cpu.REG_FILE.rf[21][16] ),
    .B(\u_cpu.REG_FILE._02880_ ),
    .X(\u_cpu.REG_FILE._03706_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.REG_FILE._08421_  (.A1(\u_cpu.REG_FILE._03403_ ),
    .A2(\u_cpu.REG_FILE._03705_ ),
    .A3(\u_cpu.REG_FILE._03706_ ),
    .B1(\u_cpu.REG_FILE._02804_ ),
    .Y(\u_cpu.REG_FILE._03707_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.REG_FILE._08422_  (.A1(\u_cpu.REG_FILE._02937_ ),
    .A2(\u_cpu.REG_FILE._03702_ ),
    .B1(\u_cpu.REG_FILE._03704_ ),
    .B2(\u_cpu.REG_FILE._03707_ ),
    .C1(\u_cpu.REG_FILE._03023_ ),
    .X(\u_cpu.REG_FILE._03708_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08423_  (.A(\u_cpu.REG_FILE._03201_ ),
    .X(\u_cpu.REG_FILE._03709_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08424_  (.A(\u_cpu.REG_FILE.rf[24][16] ),
    .B(\u_cpu.REG_FILE._03058_ ),
    .Y(\u_cpu.REG_FILE._03710_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08425_  (.A_N(\u_cpu.REG_FILE.rf[25][16] ),
    .B(\u_cpu.REG_FILE._03060_ ),
    .X(\u_cpu.REG_FILE._03711_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08426_  (.A(\u_cpu.REG_FILE.rf[27][16] ),
    .B_N(\u_cpu.REG_FILE._03065_ ),
    .X(\u_cpu.REG_FILE._03712_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08427_  (.A1(\u_cpu.REG_FILE.rf[26][16] ),
    .A2(\u_cpu.REG_FILE._03063_ ),
    .B1(\u_cpu.REG_FILE._03064_ ),
    .C1(\u_cpu.REG_FILE._03712_ ),
    .Y(\u_cpu.REG_FILE._03713_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._08428_  (.A1(\u_cpu.REG_FILE._03709_ ),
    .A2(\u_cpu.REG_FILE._03710_ ),
    .A3(\u_cpu.REG_FILE._03711_ ),
    .B1(\u_cpu.REG_FILE._03062_ ),
    .C1(\u_cpu.REG_FILE._03713_ ),
    .Y(\u_cpu.REG_FILE._03714_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08429_  (.A_N(\u_cpu.REG_FILE.rf[29][16] ),
    .B(\u_cpu.REG_FILE._03069_ ),
    .X(\u_cpu.REG_FILE._03715_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08430_  (.A1(\u_cpu.REG_FILE.rf[28][16] ),
    .A2(\u_cpu.REG_FILE._03071_ ),
    .B1_N(\u_cpu.REG_FILE._03072_ ),
    .Y(\u_cpu.REG_FILE._03716_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08431_  (.A(\u_cpu.REG_FILE.rf[31][16] ),
    .B_N(\u_cpu.REG_FILE._03034_ ),
    .X(\u_cpu.REG_FILE._03717_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08432_  (.A1(\u_cpu.REG_FILE.rf[30][16] ),
    .A2(\u_cpu.REG_FILE._03075_ ),
    .B1(\u_cpu.REG_FILE._03076_ ),
    .C1(\u_cpu.REG_FILE._03717_ ),
    .Y(\u_cpu.REG_FILE._03718_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08433_  (.A1(\u_cpu.REG_FILE._03715_ ),
    .A2(\u_cpu.REG_FILE._03716_ ),
    .B1(\u_cpu.REG_FILE._03074_ ),
    .C1(\u_cpu.REG_FILE._03718_ ),
    .Y(\u_cpu.REG_FILE._03719_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._08434_  (.A1(\u_cpu.REG_FILE._03714_ ),
    .A2(\u_cpu.REG_FILE._02992_ ),
    .A3(\u_cpu.REG_FILE._03719_ ),
    .B1(\u_cpu.REG_FILE._03081_ ),
    .X(\u_cpu.REG_FILE._03720_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08435_  (.A(\u_cpu.REG_FILE.rf[8][16] ),
    .B(\u_cpu.REG_FILE._02998_ ),
    .Y(\u_cpu.REG_FILE._03721_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08436_  (.A1(\u_cpu.REG_FILE.rf[9][16] ),
    .A2(\u_cpu.REG_FILE._03132_ ),
    .B1_N(\u_cpu.REG_FILE._03133_ ),
    .Y(\u_cpu.REG_FILE._03722_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._08437_  (.A(\u_cpu.REG_FILE.rf[10][16] ),
    .B(\u_cpu.REG_FILE._02867_ ),
    .X(\u_cpu.REG_FILE._03723_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08438_  (.A1(\u_cpu.REG_FILE.rf[11][16] ),
    .A2(\u_cpu.REG_FILE._03136_ ),
    .B1(\u_cpu.REG_FILE._03137_ ),
    .C1(\u_cpu.REG_FILE._03723_ ),
    .Y(\u_cpu.REG_FILE._03724_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08439_  (.A1(\u_cpu.REG_FILE._03721_ ),
    .A2(\u_cpu.REG_FILE._03722_ ),
    .B1(\u_cpu.REG_FILE._03135_ ),
    .C1(\u_cpu.REG_FILE._03724_ ),
    .Y(\u_cpu.REG_FILE._03725_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._08440_  (.A(\u_cpu.REG_FILE.rf[14][16] ),
    .B(\u_cpu.REG_FILE._03143_ ),
    .X(\u_cpu.REG_FILE._03726_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08441_  (.A1(\u_cpu.REG_FILE.rf[15][16] ),
    .A2(\u_cpu.REG_FILE._03142_ ),
    .B1(\u_cpu.REG_FILE._03255_ ),
    .C1(\u_cpu.REG_FILE._03726_ ),
    .Y(\u_cpu.REG_FILE._03727_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08442_  (.A1(\u_cpu.REG_FILE.rf[12][16] ),
    .A2(\u_cpu.REG_FILE._03016_ ),
    .B1_N(\u_cpu.REG_FILE._02931_ ),
    .X(\u_cpu.REG_FILE._03728_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08443_  (.A1(\u_cpu.REG_FILE.rf[13][16] ),
    .A2(\u_cpu.REG_FILE._02870_ ),
    .B1(\u_cpu.REG_FILE._03728_ ),
    .Y(\u_cpu.REG_FILE._03729_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08444_  (.A(\u_cpu.REG_FILE._03727_ ),
    .B(\u_cpu.REG_FILE._03729_ ),
    .C(\u_cpu.REG_FILE._03074_ ),
    .Y(\u_cpu.REG_FILE._03730_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08445_  (.A(\u_cpu.REG_FILE._03725_ ),
    .B(\u_cpu.REG_FILE._03141_ ),
    .C(\u_cpu.REG_FILE._03730_ ),
    .Y(\u_cpu.REG_FILE._03731_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08446_  (.A(\u_cpu.REG_FILE.rf[0][16] ),
    .B(\u_cpu.REG_FILE._03309_ ),
    .Y(\u_cpu.REG_FILE._03732_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08447_  (.A_N(\u_cpu.REG_FILE.rf[1][16] ),
    .B(\u_cpu.REG_FILE._03311_ ),
    .X(\u_cpu.REG_FILE._03733_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08448_  (.A(\u_cpu.REG_FILE.rf[3][16] ),
    .B_N(\u_cpu.REG_FILE._02852_ ),
    .X(\u_cpu.REG_FILE._03734_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08449_  (.A1(\u_cpu.REG_FILE.rf[2][16] ),
    .A2(\u_cpu.REG_FILE._02837_ ),
    .B1(\u_cpu.REG_FILE._03407_ ),
    .C1(\u_cpu.REG_FILE._03734_ ),
    .Y(\u_cpu.REG_FILE._03735_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._08450_  (.A1(\u_cpu.REG_FILE._03308_ ),
    .A2(\u_cpu.REG_FILE._03732_ ),
    .A3(\u_cpu.REG_FILE._03733_ ),
    .B1(\u_cpu.REG_FILE._03008_ ),
    .C1(\u_cpu.REG_FILE._03735_ ),
    .Y(\u_cpu.REG_FILE._03736_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08451_  (.A(\u_cpu.REG_FILE.rf[7][16] ),
    .B_N(\u_cpu.REG_FILE._02783_ ),
    .X(\u_cpu.REG_FILE._03737_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08452_  (.A1(\u_cpu.REG_FILE.rf[6][16] ),
    .A2(\u_cpu.REG_FILE._02843_ ),
    .B1(\u_cpu.REG_FILE._02866_ ),
    .C1(\u_cpu.REG_FILE._03737_ ),
    .Y(\u_cpu.REG_FILE._03738_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08453_  (.A1(\u_cpu.REG_FILE.rf[4][16] ),
    .A2(\u_cpu.REG_FILE._03030_ ),
    .B1_N(\u_cpu.REG_FILE._03039_ ),
    .X(\u_cpu.REG_FILE._03739_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08454_  (.A1(\u_cpu.REG_FILE.rf[5][16] ),
    .A2(\u_cpu.REG_FILE._03037_ ),
    .B1(\u_cpu.REG_FILE._03739_ ),
    .Y(\u_cpu.REG_FILE._03740_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08455_  (.A(\u_cpu.REG_FILE._03738_ ),
    .B(\u_cpu.REG_FILE._03740_ ),
    .C(\u_cpu.REG_FILE._03042_ ),
    .Y(\u_cpu.REG_FILE._03741_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08456_  (.A(\u_cpu.REG_FILE._02851_ ),
    .B(\u_cpu.REG_FILE._03736_ ),
    .C(\u_cpu.REG_FILE._03741_ ),
    .Y(\u_cpu.REG_FILE._03742_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08457_  (.A(\u_cpu.REG_FILE._02997_ ),
    .B(\u_cpu.REG_FILE._03731_ ),
    .C(\u_cpu.REG_FILE._03742_ ),
    .Y(\u_cpu.REG_FILE._03743_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08458_  (.A1(\u_cpu.REG_FILE._03708_ ),
    .A2(\u_cpu.REG_FILE._03720_ ),
    .B1(\u_cpu.REG_FILE._03743_ ),
    .C1(\u_cpu.REG_FILE._03467_ ),
    .X(\u_cpu.ALU.SrcB[16] ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08459_  (.A1(\u_cpu.REG_FILE.rf[18][17] ),
    .A2(\u_cpu.REG_FILE._03653_ ),
    .B1(\u_cpu.REG_FILE._02941_ ),
    .Y(\u_cpu.REG_FILE._03744_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._08460_  (.A1(\u_cpu.REG_FILE._02074_ ),
    .A2(\u_cpu.REG_FILE._02939_ ),
    .B1(\u_cpu.REG_FILE._03744_ ),
    .Y(\u_cpu.REG_FILE._03745_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08461_  (.A(\u_cpu.REG_FILE.rf[16][17] ),
    .B(\u_cpu.REG_FILE._03371_ ),
    .Y(\u_cpu.REG_FILE._03746_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._08462_  (.A1(\u_cpu.REG_FILE._02077_ ),
    .A2(\u_cpu.REG_FILE._03166_ ),
    .B1(\u_cpu.REG_FILE._02948_ ),
    .C1(\u_cpu.REG_FILE._03746_ ),
    .Y(\u_cpu.REG_FILE._03747_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08463_  (.A1(\u_cpu.REG_FILE.rf[20][17] ),
    .A2(\u_cpu.REG_FILE._02953_ ),
    .B1_N(\u_cpu.REG_FILE._03050_ ),
    .Y(\u_cpu.REG_FILE._03748_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08464_  (.A(\u_cpu.REG_FILE.rf[21][17] ),
    .B(\u_cpu.REG_FILE._02859_ ),
    .Y(\u_cpu.REG_FILE._03749_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08465_  (.A(\u_cpu.REG_FILE.rf[22][17] ),
    .B(\u_cpu.REG_FILE._02958_ ),
    .Y(\u_cpu.REG_FILE._03750_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08466_  (.A1(\u_cpu.REG_FILE.rf[23][17] ),
    .A2(\u_cpu.REG_FILE._03114_ ),
    .B1(\u_cpu.REG_FILE._03377_ ),
    .Y(\u_cpu.REG_FILE._03751_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._08467_  (.A1(\u_cpu.REG_FILE._03748_ ),
    .A2(\u_cpu.REG_FILE._03749_ ),
    .B1(\u_cpu.REG_FILE._03750_ ),
    .B2(\u_cpu.REG_FILE._03751_ ),
    .C1(\u_cpu.REG_FILE._02848_ ),
    .Y(\u_cpu.REG_FILE._03752_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.REG_FILE._08468_  (.A1(\u_cpu.REG_FILE._02937_ ),
    .A2(\u_cpu.REG_FILE._03745_ ),
    .A3(\u_cpu.REG_FILE._03747_ ),
    .B1(\u_cpu.REG_FILE._03752_ ),
    .C1(\u_cpu.REG_FILE._02966_ ),
    .X(\u_cpu.REG_FILE._03753_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08469_  (.A(\u_cpu.REG_FILE.rf[31][17] ),
    .B_N(\u_cpu.REG_FILE._02970_ ),
    .X(\u_cpu.REG_FILE._03754_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08470_  (.A1(\u_cpu.REG_FILE.rf[30][17] ),
    .A2(\u_cpu.REG_FILE._02749_ ),
    .B1(\u_cpu.REG_FILE._02969_ ),
    .C1(\u_cpu.REG_FILE._03754_ ),
    .Y(\u_cpu.REG_FILE._03755_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08471_  (.A1(\u_cpu.REG_FILE.rf[28][17] ),
    .A2(\u_cpu.REG_FILE._02974_ ),
    .B1_N(\u_cpu.REG_FILE._02975_ ),
    .X(\u_cpu.REG_FILE._03756_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08472_  (.A1(\u_cpu.REG_FILE.rf[29][17] ),
    .A2(\u_cpu.REG_FILE._02973_ ),
    .B1(\u_cpu.REG_FILE._03756_ ),
    .Y(\u_cpu.REG_FILE._03757_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08473_  (.A(\u_cpu.REG_FILE._03755_ ),
    .B(\u_cpu.REG_FILE._03757_ ),
    .C(\u_cpu.REG_FILE._03006_ ),
    .Y(\u_cpu.REG_FILE._03758_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08474_  (.A_N(\u_cpu.REG_FILE.rf[25][17] ),
    .B(\u_cpu.REG_FILE._02980_ ),
    .X(\u_cpu.REG_FILE._03759_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08475_  (.A1(\u_cpu.REG_FILE.rf[24][17] ),
    .A2(\u_cpu.REG_FILE._03212_ ),
    .B1_N(\u_cpu.REG_FILE._02983_ ),
    .Y(\u_cpu.REG_FILE._03760_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08476_  (.A(\u_cpu.REG_FILE.rf[27][17] ),
    .B_N(\u_cpu.REG_FILE._03077_ ),
    .X(\u_cpu.REG_FILE._03761_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08477_  (.A1(\u_cpu.REG_FILE.rf[26][17] ),
    .A2(\u_cpu.REG_FILE._03125_ ),
    .B1(\u_cpu.REG_FILE._02988_ ),
    .C1(\u_cpu.REG_FILE._03761_ ),
    .Y(\u_cpu.REG_FILE._03762_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08478_  (.A1(\u_cpu.REG_FILE._03759_ ),
    .A2(\u_cpu.REG_FILE._03760_ ),
    .B1(\u_cpu.REG_FILE._02985_ ),
    .C1(\u_cpu.REG_FILE._03762_ ),
    .Y(\u_cpu.REG_FILE._03763_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._08479_  (.A1(\u_cpu.REG_FILE._03758_ ),
    .A2(\u_cpu.REG_FILE._03763_ ),
    .A3(\u_cpu.REG_FILE._03129_ ),
    .B1(\u_cpu.REG_FILE._03081_ ),
    .X(\u_cpu.REG_FILE._03764_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08480_  (.A(\u_cpu.REG_FILE.rf[14][17] ),
    .B(\u_cpu.REG_FILE._02998_ ),
    .Y(\u_cpu.REG_FILE._03765_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08481_  (.A1(\u_cpu.REG_FILE.rf[15][17] ),
    .A2(\u_cpu.REG_FILE._02960_ ),
    .B1(\u_cpu.REG_FILE._02961_ ),
    .Y(\u_cpu.REG_FILE._03766_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08482_  (.A1(\u_cpu.REG_FILE.rf[12][17] ),
    .A2(\u_cpu.REG_FILE._02860_ ),
    .B1_N(\u_cpu.REG_FILE._02817_ ),
    .X(\u_cpu.REG_FILE._03767_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08483_  (.A1(\u_cpu.REG_FILE.rf[13][17] ),
    .A2(\u_cpu.REG_FILE._02956_ ),
    .B1(\u_cpu.REG_FILE._03767_ ),
    .Y(\u_cpu.REG_FILE._03768_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08484_  (.A1(\u_cpu.REG_FILE._03765_ ),
    .A2(\u_cpu.REG_FILE._03766_ ),
    .B1(\u_cpu.REG_FILE._03768_ ),
    .C1(\u_cpu.REG_FILE._02963_ ),
    .Y(\u_cpu.REG_FILE._03769_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08485_  (.A(\u_cpu.REG_FILE.rf[11][17] ),
    .B_N(\u_cpu.REG_FILE._03012_ ),
    .X(\u_cpu.REG_FILE._03770_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08486_  (.A1(\u_cpu.REG_FILE.rf[10][17] ),
    .A2(\u_cpu.REG_FILE._03010_ ),
    .B1(\u_cpu.REG_FILE._03011_ ),
    .C1(\u_cpu.REG_FILE._03770_ ),
    .Y(\u_cpu.REG_FILE._03771_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08487_  (.A1(\u_cpu.REG_FILE.rf[8][17] ),
    .A2(\u_cpu.REG_FILE._03090_ ),
    .B1_N(\u_cpu.REG_FILE._03017_ ),
    .X(\u_cpu.REG_FILE._03772_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08488_  (.A1(\u_cpu.REG_FILE.rf[9][17] ),
    .A2(\u_cpu.REG_FILE._03015_ ),
    .B1(\u_cpu.REG_FILE._03772_ ),
    .Y(\u_cpu.REG_FILE._03773_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08489_  (.A(\u_cpu.REG_FILE._03135_ ),
    .B(\u_cpu.REG_FILE._03771_ ),
    .C(\u_cpu.REG_FILE._03773_ ),
    .Y(\u_cpu.REG_FILE._03774_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08490_  (.A(\u_cpu.REG_FILE._03769_ ),
    .B(\u_cpu.REG_FILE._03774_ ),
    .C(\u_cpu.REG_FILE._03021_ ),
    .Y(\u_cpu.REG_FILE._03775_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08491_  (.A(\u_cpu.REG_FILE.rf[3][17] ),
    .B_N(\u_cpu.REG_FILE._02815_ ),
    .X(\u_cpu.REG_FILE._03776_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08492_  (.A1(\u_cpu.REG_FILE.rf[2][17] ),
    .A2(\u_cpu.REG_FILE._03025_ ),
    .B1(\u_cpu.REG_FILE._03026_ ),
    .C1(\u_cpu.REG_FILE._03776_ ),
    .Y(\u_cpu.REG_FILE._03777_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08493_  (.A1(\u_cpu.REG_FILE.rf[0][17] ),
    .A2(\u_cpu.REG_FILE._03030_ ),
    .B1_N(\u_cpu.REG_FILE._02872_ ),
    .X(\u_cpu.REG_FILE._03778_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08494_  (.A1(\u_cpu.REG_FILE.rf[1][17] ),
    .A2(\u_cpu.REG_FILE._03029_ ),
    .B1(\u_cpu.REG_FILE._03778_ ),
    .Y(\u_cpu.REG_FILE._03779_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08495_  (.A(\u_cpu.REG_FILE._03009_ ),
    .B(\u_cpu.REG_FILE._03777_ ),
    .C(\u_cpu.REG_FILE._03779_ ),
    .Y(\u_cpu.REG_FILE._03780_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08496_  (.A(\u_cpu.REG_FILE.rf[7][17] ),
    .B_N(\u_cpu.REG_FILE._02783_ ),
    .X(\u_cpu.REG_FILE._03781_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08497_  (.A1(\u_cpu.REG_FILE.rf[6][17] ),
    .A2(\u_cpu.REG_FILE._02843_ ),
    .B1(\u_cpu.REG_FILE._02866_ ),
    .C1(\u_cpu.REG_FILE._03781_ ),
    .Y(\u_cpu.REG_FILE._03782_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08498_  (.A1(\u_cpu.REG_FILE.rf[4][17] ),
    .A2(\u_cpu.REG_FILE._03030_ ),
    .B1_N(\u_cpu.REG_FILE._03039_ ),
    .X(\u_cpu.REG_FILE._03783_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08499_  (.A1(\u_cpu.REG_FILE.rf[5][17] ),
    .A2(\u_cpu.REG_FILE._03029_ ),
    .B1(\u_cpu.REG_FILE._03783_ ),
    .Y(\u_cpu.REG_FILE._03784_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08500_  (.A(\u_cpu.REG_FILE._03782_ ),
    .B(\u_cpu.REG_FILE._03784_ ),
    .C(\u_cpu.REG_FILE._03042_ ),
    .Y(\u_cpu.REG_FILE._03785_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08501_  (.A(\u_cpu.REG_FILE._02851_ ),
    .B(\u_cpu.REG_FILE._03780_ ),
    .C(\u_cpu.REG_FILE._03785_ ),
    .Y(\u_cpu.REG_FILE._03786_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08502_  (.A(\u_cpu.REG_FILE._02997_ ),
    .B(\u_cpu.REG_FILE._03775_ ),
    .C(\u_cpu.REG_FILE._03786_ ),
    .Y(\u_cpu.REG_FILE._03787_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08503_  (.A1(\u_cpu.REG_FILE._03753_ ),
    .A2(\u_cpu.REG_FILE._03764_ ),
    .B1(\u_cpu.REG_FILE._03787_ ),
    .C1(\u_cpu.REG_FILE._03467_ ),
    .X(\u_cpu.ALU.SrcB[17] ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08504_  (.A1(\u_cpu.REG_FILE.rf[18][18] ),
    .A2(\u_cpu.REG_FILE._03653_ ),
    .B1(\u_cpu.REG_FILE._03298_ ),
    .Y(\u_cpu.REG_FILE._03788_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._08505_  (.A1(\u_cpu.REG_FILE._02112_ ),
    .A2(\u_cpu.REG_FILE._02939_ ),
    .B1(\u_cpu.REG_FILE._03788_ ),
    .Y(\u_cpu.REG_FILE._03789_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08506_  (.A(\u_cpu.REG_FILE.rf[16][18] ),
    .B(\u_cpu.REG_FILE._03371_ ),
    .Y(\u_cpu.REG_FILE._03790_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._08507_  (.A1(\u_cpu.REG_FILE._02115_ ),
    .A2(\u_cpu.REG_FILE._03166_ ),
    .B1(\u_cpu.REG_FILE._02948_ ),
    .C1(\u_cpu.REG_FILE._03790_ ),
    .Y(\u_cpu.REG_FILE._03791_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08508_  (.A1(\u_cpu.REG_FILE.rf[20][18] ),
    .A2(\u_cpu.REG_FILE._02853_ ),
    .B1_N(\u_cpu.REG_FILE._03050_ ),
    .Y(\u_cpu.REG_FILE._03792_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08509_  (.A(\u_cpu.REG_FILE.rf[21][18] ),
    .B(\u_cpu.REG_FILE._02859_ ),
    .Y(\u_cpu.REG_FILE._03793_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08510_  (.A(\u_cpu.REG_FILE.rf[22][18] ),
    .B(\u_cpu.REG_FILE._02958_ ),
    .Y(\u_cpu.REG_FILE._03794_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08511_  (.A1(\u_cpu.REG_FILE.rf[23][18] ),
    .A2(\u_cpu.REG_FILE._03114_ ),
    .B1(\u_cpu.REG_FILE._03377_ ),
    .Y(\u_cpu.REG_FILE._03795_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._08512_  (.A1(\u_cpu.REG_FILE._03792_ ),
    .A2(\u_cpu.REG_FILE._03793_ ),
    .B1(\u_cpu.REG_FILE._03794_ ),
    .B2(\u_cpu.REG_FILE._03795_ ),
    .C1(\u_cpu.REG_FILE._02848_ ),
    .Y(\u_cpu.REG_FILE._03796_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.REG_FILE._08513_  (.A1(\u_cpu.REG_FILE._02765_ ),
    .A2(\u_cpu.REG_FILE._03789_ ),
    .A3(\u_cpu.REG_FILE._03791_ ),
    .B1(\u_cpu.REG_FILE._03796_ ),
    .C1(\u_cpu.REG_FILE._02966_ ),
    .X(\u_cpu.REG_FILE._03797_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08514_  (.A(\u_cpu.REG_FILE.rf[24][18] ),
    .B(\u_cpu.REG_FILE._03058_ ),
    .Y(\u_cpu.REG_FILE._03798_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08515_  (.A_N(\u_cpu.REG_FILE.rf[25][18] ),
    .B(\u_cpu.REG_FILE._03060_ ),
    .X(\u_cpu.REG_FILE._03799_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08516_  (.A(\u_cpu.REG_FILE._02776_ ),
    .X(\u_cpu.REG_FILE._03800_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08517_  (.A(\u_cpu.REG_FILE.rf[27][18] ),
    .B_N(\u_cpu.REG_FILE._03065_ ),
    .X(\u_cpu.REG_FILE._03801_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08518_  (.A1(\u_cpu.REG_FILE.rf[26][18] ),
    .A2(\u_cpu.REG_FILE._03063_ ),
    .B1(\u_cpu.REG_FILE._03064_ ),
    .C1(\u_cpu.REG_FILE._03801_ ),
    .Y(\u_cpu.REG_FILE._03802_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._08519_  (.A1(\u_cpu.REG_FILE._03709_ ),
    .A2(\u_cpu.REG_FILE._03798_ ),
    .A3(\u_cpu.REG_FILE._03799_ ),
    .B1(\u_cpu.REG_FILE._03800_ ),
    .C1(\u_cpu.REG_FILE._03802_ ),
    .Y(\u_cpu.REG_FILE._03803_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08520_  (.A_N(\u_cpu.REG_FILE.rf[29][18] ),
    .B(\u_cpu.REG_FILE._03069_ ),
    .X(\u_cpu.REG_FILE._03804_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08521_  (.A1(\u_cpu.REG_FILE.rf[28][18] ),
    .A2(\u_cpu.REG_FILE._03071_ ),
    .B1_N(\u_cpu.REG_FILE._03072_ ),
    .Y(\u_cpu.REG_FILE._03805_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08522_  (.A(\u_cpu.REG_FILE.rf[31][18] ),
    .B_N(\u_cpu.REG_FILE._03034_ ),
    .X(\u_cpu.REG_FILE._03806_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08523_  (.A1(\u_cpu.REG_FILE.rf[30][18] ),
    .A2(\u_cpu.REG_FILE._03075_ ),
    .B1(\u_cpu.REG_FILE._03076_ ),
    .C1(\u_cpu.REG_FILE._03806_ ),
    .Y(\u_cpu.REG_FILE._03807_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08524_  (.A1(\u_cpu.REG_FILE._03804_ ),
    .A2(\u_cpu.REG_FILE._03805_ ),
    .B1(\u_cpu.REG_FILE._03074_ ),
    .C1(\u_cpu.REG_FILE._03807_ ),
    .Y(\u_cpu.REG_FILE._03808_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._08525_  (.A1(\u_cpu.REG_FILE._03803_ ),
    .A2(\u_cpu.REG_FILE._02992_ ),
    .A3(\u_cpu.REG_FILE._03808_ ),
    .B1(\u_cpu.REG_FILE._03081_ ),
    .X(\u_cpu.REG_FILE._03809_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08526_  (.A(\u_cpu.REG_FILE.rf[0][18] ),
    .B(\u_cpu.REG_FILE._02816_ ),
    .Y(\u_cpu.REG_FILE._03810_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08527_  (.A_N(\u_cpu.REG_FILE.rf[1][18] ),
    .B(\u_cpu.REG_FILE._03530_ ),
    .X(\u_cpu.REG_FILE._03811_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08528_  (.A(\u_cpu.REG_FILE.rf[3][18] ),
    .B_N(\u_cpu.REG_FILE._02949_ ),
    .X(\u_cpu.REG_FILE._03812_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08529_  (.A1(\u_cpu.REG_FILE.rf[2][18] ),
    .A2(\u_cpu.REG_FILE._02987_ ),
    .B1(\u_cpu.REG_FILE._03377_ ),
    .C1(\u_cpu.REG_FILE._03812_ ),
    .Y(\u_cpu.REG_FILE._03813_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.REG_FILE._08530_  (.A1(\u_cpu.REG_FILE._03709_ ),
    .A2(\u_cpu.REG_FILE._03810_ ),
    .A3(\u_cpu.REG_FILE._03811_ ),
    .B1(\u_cpu.REG_FILE._03800_ ),
    .C1(\u_cpu.REG_FILE._03813_ ),
    .X(\u_cpu.REG_FILE._03814_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08531_  (.A(\u_cpu.REG_FILE._02792_ ),
    .X(\u_cpu.REG_FILE._03815_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08532_  (.A(\u_cpu.REG_FILE.rf[4][18] ),
    .B(\u_cpu.REG_FILE._03815_ ),
    .Y(\u_cpu.REG_FILE._03816_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._08533_  (.A1(\u_cpu.REG_FILE._02098_ ),
    .A2(\u_cpu.REG_FILE._03418_ ),
    .B1(\u_cpu.REG_FILE._03308_ ),
    .C1(\u_cpu.REG_FILE._03816_ ),
    .Y(\u_cpu.REG_FILE._03817_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08534_  (.A1(\u_cpu.REG_FILE.rf[6][18] ),
    .A2(\u_cpu.REG_FILE._03204_ ),
    .B1(\u_cpu.REG_FILE._03198_ ),
    .Y(\u_cpu.REG_FILE._03818_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08535_  (.A_N(\u_cpu.REG_FILE.rf[7][18] ),
    .B(\u_cpu.REG_FILE._02880_ ),
    .X(\u_cpu.REG_FILE._03819_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08536_  (.A1(\u_cpu.REG_FILE._03818_ ),
    .A2(\u_cpu.REG_FILE._03819_ ),
    .B1(\u_cpu.REG_FILE._03434_ ),
    .Y(\u_cpu.REG_FILE._03820_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08537_  (.A1(\u_cpu.REG_FILE._03817_ ),
    .A2(\u_cpu.REG_FILE._03820_ ),
    .B1_N(\u_cpu.REG_FILE._03141_ ),
    .Y(\u_cpu.REG_FILE._03821_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08538_  (.A_N(\u_cpu.REG_FILE.rf[13][18] ),
    .B(\u_cpu.REG_FILE._02760_ ),
    .X(\u_cpu.REG_FILE._03822_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08539_  (.A1(\u_cpu.REG_FILE.rf[12][18] ),
    .A2(\u_cpu.REG_FILE._03815_ ),
    .B1_N(\u_cpu.REG_FILE._02954_ ),
    .Y(\u_cpu.REG_FILE._03823_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08540_  (.A(\u_cpu.REG_FILE.rf[15][18] ),
    .B_N(\u_cpu.REG_FILE._02810_ ),
    .X(\u_cpu.REG_FILE._03824_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08541_  (.A1(\u_cpu.REG_FILE.rf[14][18] ),
    .A2(\u_cpu.REG_FILE._03287_ ),
    .B1(\u_cpu.REG_FILE._03470_ ),
    .C1(\u_cpu.REG_FILE._03824_ ),
    .Y(\u_cpu.REG_FILE._03825_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08542_  (.A1(\u_cpu.REG_FILE._03822_ ),
    .A2(\u_cpu.REG_FILE._03823_ ),
    .B1(\u_cpu.REG_FILE._03825_ ),
    .Y(\u_cpu.REG_FILE._03826_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08543_  (.A(\u_cpu.REG_FILE.rf[10][18] ),
    .B(\u_cpu.REG_FILE._03025_ ),
    .Y(\u_cpu.REG_FILE._03827_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08544_  (.A1(\u_cpu.REG_FILE.rf[11][18] ),
    .A2(\u_cpu.REG_FILE._03297_ ),
    .B1(\u_cpu.REG_FILE._03470_ ),
    .Y(\u_cpu.REG_FILE._03828_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08545_  (.A1(\u_cpu.REG_FILE.rf[8][18] ),
    .A2(\u_cpu.REG_FILE._03337_ ),
    .B1_N(\u_cpu.REG_FILE._02798_ ),
    .X(\u_cpu.REG_FILE._03829_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08546_  (.A1(\u_cpu.REG_FILE.rf[9][18] ),
    .A2(\u_cpu.REG_FILE._02845_ ),
    .B1(\u_cpu.REG_FILE._03829_ ),
    .Y(\u_cpu.REG_FILE._03830_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08547_  (.A1(\u_cpu.REG_FILE._03827_ ),
    .A2(\u_cpu.REG_FILE._03828_ ),
    .B1(\u_cpu.REG_FILE._03830_ ),
    .C1(\u_cpu.REG_FILE._03800_ ),
    .Y(\u_cpu.REG_FILE._03831_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08548_  (.A1(\u_cpu.REG_FILE._03024_ ),
    .A2(\u_cpu.REG_FILE._03826_ ),
    .B1(\u_cpu.REG_FILE._03831_ ),
    .C1(\u_cpu.REG_FILE._03218_ ),
    .Y(\u_cpu.REG_FILE._03832_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08549_  (.A1(\u_cpu.REG_FILE._03814_ ),
    .A2(\u_cpu.REG_FILE._03821_ ),
    .B1(\u_cpu.REG_FILE._02994_ ),
    .C1(\u_cpu.REG_FILE._03832_ ),
    .Y(\u_cpu.REG_FILE._03833_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08550_  (.A1(\u_cpu.REG_FILE._03797_ ),
    .A2(\u_cpu.REG_FILE._03809_ ),
    .B1(\u_cpu.REG_FILE._03833_ ),
    .C1(\u_cpu.REG_FILE._03467_ ),
    .X(\u_cpu.ALU.SrcB[18] ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._08551_  (.A(\u_cpu.REG_FILE.rf[22][19] ),
    .B(\u_cpu.REG_FILE._02853_ ),
    .X(\u_cpu.REG_FILE._03834_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08552_  (.A1(\u_cpu.REG_FILE.rf[23][19] ),
    .A2(\u_cpu.REG_FILE._02759_ ),
    .B1(\u_cpu.REG_FILE._02948_ ),
    .C1(\u_cpu.REG_FILE._03834_ ),
    .Y(\u_cpu.REG_FILE._03835_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08553_  (.A1(\u_cpu.REG_FILE.rf[20][19] ),
    .A2(\u_cpu.REG_FILE._03815_ ),
    .B1_N(\u_cpu.REG_FILE._03133_ ),
    .X(\u_cpu.REG_FILE._03836_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08554_  (.A(\u_cpu.REG_FILE.rf[21][19] ),
    .B_N(\u_cpu.REG_FILE._03331_ ),
    .X(\u_cpu.REG_FILE._03837_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._08555_  (.A1(\u_cpu.REG_FILE._03836_ ),
    .A2(\u_cpu.REG_FILE._03837_ ),
    .B1(\u_cpu.REG_FILE._03024_ ),
    .Y(\u_cpu.REG_FILE._03838_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08556_  (.A1(\u_cpu.REG_FILE.rf[16][19] ),
    .A2(\u_cpu.REG_FILE._03815_ ),
    .B1_N(\u_cpu.REG_FILE._02838_ ),
    .Y(\u_cpu.REG_FILE._03839_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08557_  (.A_N(\u_cpu.REG_FILE.rf[17][19] ),
    .B(\u_cpu.REG_FILE._03530_ ),
    .X(\u_cpu.REG_FILE._03840_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08558_  (.A1(\u_cpu.REG_FILE.rf[18][19] ),
    .A2(\u_cpu.REG_FILE._03653_ ),
    .B1(\u_cpu.REG_FILE._03298_ ),
    .Y(\u_cpu.REG_FILE._03841_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08559_  (.A_N(\u_cpu.REG_FILE.rf[19][19] ),
    .B(\u_cpu.REG_FILE._02945_ ),
    .X(\u_cpu.REG_FILE._03842_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.REG_FILE._08560_  (.A1(\u_cpu.REG_FILE._03839_ ),
    .A2(\u_cpu.REG_FILE._03840_ ),
    .B1(\u_cpu.REG_FILE._03841_ ),
    .B2(\u_cpu.REG_FILE._03842_ ),
    .C1(\u_cpu.REG_FILE._02985_ ),
    .X(\u_cpu.REG_FILE._03843_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._08561_  (.A1(\u_cpu.REG_FILE._03835_ ),
    .A2(\u_cpu.REG_FILE._03838_ ),
    .B1(\u_cpu.REG_FILE._02788_ ),
    .C1(\u_cpu.REG_FILE._03843_ ),
    .Y(\u_cpu.REG_FILE._03844_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08562_  (.A(\u_cpu.REG_FILE.rf[24][19] ),
    .B(\u_cpu.REG_FILE._03058_ ),
    .Y(\u_cpu.REG_FILE._03845_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08563_  (.A_N(\u_cpu.REG_FILE.rf[25][19] ),
    .B(\u_cpu.REG_FILE._03060_ ),
    .X(\u_cpu.REG_FILE._03846_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08564_  (.A(\u_cpu.REG_FILE.rf[27][19] ),
    .B_N(\u_cpu.REG_FILE._03065_ ),
    .X(\u_cpu.REG_FILE._03847_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08565_  (.A1(\u_cpu.REG_FILE.rf[26][19] ),
    .A2(\u_cpu.REG_FILE._03063_ ),
    .B1(\u_cpu.REG_FILE._03064_ ),
    .C1(\u_cpu.REG_FILE._03847_ ),
    .Y(\u_cpu.REG_FILE._03848_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._08566_  (.A1(\u_cpu.REG_FILE._03709_ ),
    .A2(\u_cpu.REG_FILE._03845_ ),
    .A3(\u_cpu.REG_FILE._03846_ ),
    .B1(\u_cpu.REG_FILE._03800_ ),
    .C1(\u_cpu.REG_FILE._03848_ ),
    .Y(\u_cpu.REG_FILE._03849_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08567_  (.A_N(\u_cpu.REG_FILE.rf[29][19] ),
    .B(\u_cpu.REG_FILE._03069_ ),
    .X(\u_cpu.REG_FILE._03850_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08568_  (.A1(\u_cpu.REG_FILE.rf[28][19] ),
    .A2(\u_cpu.REG_FILE._03071_ ),
    .B1_N(\u_cpu.REG_FILE._03072_ ),
    .Y(\u_cpu.REG_FILE._03851_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08569_  (.A(\u_cpu.REG_FILE.rf[31][19] ),
    .B_N(\u_cpu.REG_FILE._03034_ ),
    .X(\u_cpu.REG_FILE._03852_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08570_  (.A1(\u_cpu.REG_FILE.rf[30][19] ),
    .A2(\u_cpu.REG_FILE._03075_ ),
    .B1(\u_cpu.REG_FILE._03076_ ),
    .C1(\u_cpu.REG_FILE._03852_ ),
    .Y(\u_cpu.REG_FILE._03853_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08571_  (.A1(\u_cpu.REG_FILE._03850_ ),
    .A2(\u_cpu.REG_FILE._03851_ ),
    .B1(\u_cpu.REG_FILE._03221_ ),
    .C1(\u_cpu.REG_FILE._03853_ ),
    .Y(\u_cpu.REG_FILE._03854_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._08572_  (.A1(\u_cpu.REG_FILE._03849_ ),
    .A2(\u_cpu.REG_FILE._02992_ ),
    .A3(\u_cpu.REG_FILE._03854_ ),
    .B1(\u_cpu.REG_FILE._03081_ ),
    .X(\u_cpu.REG_FILE._03855_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._08573_  (.A(\u_cpu.REG_FILE.rf[5][19] ),
    .Y(\u_cpu.REG_FILE._03856_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08574_  (.A1(\u_cpu.REG_FILE.rf[4][19] ),
    .A2(\u_cpu.REG_FILE._03404_ ),
    .B1_N(\u_cpu.REG_FILE._03201_ ),
    .Y(\u_cpu.REG_FILE._03857_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._08575_  (.A1(\u_cpu.REG_FILE._03856_ ),
    .A2(\u_cpu.REG_FILE._02946_ ),
    .B1(\u_cpu.REG_FILE._03857_ ),
    .Y(\u_cpu.REG_FILE._03858_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08576_  (.A1(\u_cpu.REG_FILE.rf[6][19] ),
    .A2(\u_cpu.REG_FILE._03204_ ),
    .B1(\u_cpu.REG_FILE._03198_ ),
    .Y(\u_cpu.REG_FILE._03859_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08577_  (.A_N(\u_cpu.REG_FILE.rf[7][19] ),
    .B(\u_cpu.REG_FILE._02880_ ),
    .X(\u_cpu.REG_FILE._03860_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08578_  (.A1(\u_cpu.REG_FILE._03859_ ),
    .A2(\u_cpu.REG_FILE._03860_ ),
    .B1(\u_cpu.REG_FILE._02834_ ),
    .Y(\u_cpu.REG_FILE._03861_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08579_  (.A_N(\u_cpu.REG_FILE.rf[1][19] ),
    .B(\u_cpu.REG_FILE._02830_ ),
    .X(\u_cpu.REG_FILE._03862_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08580_  (.A1(\u_cpu.REG_FILE.rf[0][19] ),
    .A2(\u_cpu.REG_FILE._02853_ ),
    .B1_N(\u_cpu.REG_FILE._02838_ ),
    .Y(\u_cpu.REG_FILE._03863_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08581_  (.A(\u_cpu.REG_FILE.rf[3][19] ),
    .B_N(\u_cpu.REG_FILE._02810_ ),
    .X(\u_cpu.REG_FILE._03864_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08582_  (.A1(\u_cpu.REG_FILE.rf[2][19] ),
    .A2(\u_cpu.REG_FILE._03287_ ),
    .B1(\u_cpu.REG_FILE._03470_ ),
    .C1(\u_cpu.REG_FILE._03864_ ),
    .Y(\u_cpu.REG_FILE._03865_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08583_  (.A1(\u_cpu.REG_FILE._03862_ ),
    .A2(\u_cpu.REG_FILE._03863_ ),
    .B1(\u_cpu.REG_FILE._03292_ ),
    .C1(\u_cpu.REG_FILE._03865_ ),
    .Y(\u_cpu.REG_FILE._03866_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08584_  (.A1(\u_cpu.REG_FILE._03858_ ),
    .A2(\u_cpu.REG_FILE._03861_ ),
    .B1(\u_cpu.REG_FILE._03866_ ),
    .Y(\u_cpu.REG_FILE._03867_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08585_  (.A(\u_cpu.REG_FILE.rf[12][19] ),
    .B(\u_cpu.REG_FILE._02843_ ),
    .Y(\u_cpu.REG_FILE._03868_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08586_  (.A1(\u_cpu.REG_FILE.rf[13][19] ),
    .A2(\u_cpu.REG_FILE._02845_ ),
    .B1_N(\u_cpu.REG_FILE._02947_ ),
    .Y(\u_cpu.REG_FILE._03869_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._08587_  (.A(\u_cpu.REG_FILE.rf[14][19] ),
    .B(\u_cpu.REG_FILE._02792_ ),
    .X(\u_cpu.REG_FILE._03870_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08588_  (.A1(\u_cpu.REG_FILE.rf[15][19] ),
    .A2(\u_cpu.REG_FILE._03351_ ),
    .B1(\u_cpu.REG_FILE._02818_ ),
    .C1(\u_cpu.REG_FILE._03870_ ),
    .Y(\u_cpu.REG_FILE._03871_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08589_  (.A1(\u_cpu.REG_FILE._03868_ ),
    .A2(\u_cpu.REG_FILE._03869_ ),
    .B1(\u_cpu.REG_FILE._02804_ ),
    .C1(\u_cpu.REG_FILE._03871_ ),
    .Y(\u_cpu.REG_FILE._03872_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08590_  (.A(\u_cpu.REG_FILE.rf[11][19] ),
    .B_N(\u_cpu.REG_FILE._02792_ ),
    .X(\u_cpu.REG_FILE._03873_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08591_  (.A1(\u_cpu.REG_FILE.rf[10][19] ),
    .A2(\u_cpu.REG_FILE._02953_ ),
    .B1(\u_cpu.REG_FILE._02799_ ),
    .C1(\u_cpu.REG_FILE._03873_ ),
    .Y(\u_cpu.REG_FILE._03874_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08592_  (.A1(\u_cpu.REG_FILE.rf[8][19] ),
    .A2(\u_cpu.REG_FILE._02779_ ),
    .B1_N(\u_cpu.REG_FILE._02798_ ),
    .X(\u_cpu.REG_FILE._03875_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08593_  (.A1(\u_cpu.REG_FILE.rf[9][19] ),
    .A2(\u_cpu.REG_FILE._03351_ ),
    .B1(\u_cpu.REG_FILE._03875_ ),
    .Y(\u_cpu.REG_FILE._03876_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08594_  (.A(\u_cpu.REG_FILE._02985_ ),
    .B(\u_cpu.REG_FILE._03874_ ),
    .C(\u_cpu.REG_FILE._03876_ ),
    .Y(\u_cpu.REG_FILE._03877_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08595_  (.A(\u_cpu.REG_FILE._03872_ ),
    .B(\u_cpu.REG_FILE._03877_ ),
    .C(\u_cpu.REG_FILE._03141_ ),
    .Y(\u_cpu.REG_FILE._03878_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08596_  (.A1(\u_cpu.REG_FILE._02788_ ),
    .A2(\u_cpu.REG_FILE._03867_ ),
    .B1(\u_cpu.REG_FILE._03878_ ),
    .C1(\u_cpu.REG_FILE._02994_ ),
    .Y(\u_cpu.REG_FILE._03879_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08597_  (.A1(\u_cpu.REG_FILE._03844_ ),
    .A2(\u_cpu.REG_FILE._03855_ ),
    .B1(\u_cpu.REG_FILE._03879_ ),
    .C1(\u_cpu.REG_FILE._03467_ ),
    .X(\u_cpu.ALU.SrcB[19] ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._08598_  (.A(\u_cpu.REG_FILE.rf[22][20] ),
    .B(\u_cpu.REG_FILE._02853_ ),
    .X(\u_cpu.REG_FILE._03880_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08599_  (.A1(\u_cpu.REG_FILE.rf[23][20] ),
    .A2(\u_cpu.REG_FILE._02759_ ),
    .B1(\u_cpu.REG_FILE._02948_ ),
    .C1(\u_cpu.REG_FILE._03880_ ),
    .Y(\u_cpu.REG_FILE._03881_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08600_  (.A1(\u_cpu.REG_FILE.rf[20][20] ),
    .A2(\u_cpu.REG_FILE._03815_ ),
    .B1_N(\u_cpu.REG_FILE._03133_ ),
    .X(\u_cpu.REG_FILE._03882_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08601_  (.A(\u_cpu.REG_FILE.rf[21][20] ),
    .B_N(\u_cpu.REG_FILE._03331_ ),
    .X(\u_cpu.REG_FILE._03883_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._08602_  (.A1(\u_cpu.REG_FILE._03882_ ),
    .A2(\u_cpu.REG_FILE._03883_ ),
    .B1(\u_cpu.REG_FILE._03024_ ),
    .Y(\u_cpu.REG_FILE._03884_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08603_  (.A1(\u_cpu.REG_FILE.rf[16][20] ),
    .A2(\u_cpu.REG_FILE._03815_ ),
    .B1_N(\u_cpu.REG_FILE._02838_ ),
    .Y(\u_cpu.REG_FILE._03885_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08604_  (.A_N(\u_cpu.REG_FILE.rf[17][20] ),
    .B(\u_cpu.REG_FILE._03530_ ),
    .X(\u_cpu.REG_FILE._03886_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08605_  (.A1(\u_cpu.REG_FILE.rf[18][20] ),
    .A2(\u_cpu.REG_FILE._02811_ ),
    .B1(\u_cpu.REG_FILE._03298_ ),
    .Y(\u_cpu.REG_FILE._03887_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08606_  (.A_N(\u_cpu.REG_FILE.rf[19][20] ),
    .B(\u_cpu.REG_FILE._02945_ ),
    .X(\u_cpu.REG_FILE._03888_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.REG_FILE._08607_  (.A1(\u_cpu.REG_FILE._03885_ ),
    .A2(\u_cpu.REG_FILE._03886_ ),
    .B1(\u_cpu.REG_FILE._03887_ ),
    .B2(\u_cpu.REG_FILE._03888_ ),
    .C1(\u_cpu.REG_FILE._02985_ ),
    .X(\u_cpu.REG_FILE._03889_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._08608_  (.A1(\u_cpu.REG_FILE._03881_ ),
    .A2(\u_cpu.REG_FILE._03884_ ),
    .B1(\u_cpu.REG_FILE._02788_ ),
    .C1(\u_cpu.REG_FILE._03889_ ),
    .Y(\u_cpu.REG_FILE._03890_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08609_  (.A(\u_cpu.REG_FILE.rf[24][20] ),
    .B(\u_cpu.REG_FILE._03058_ ),
    .Y(\u_cpu.REG_FILE._03891_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08610_  (.A_N(\u_cpu.REG_FILE.rf[25][20] ),
    .B(\u_cpu.REG_FILE._03060_ ),
    .X(\u_cpu.REG_FILE._03892_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08611_  (.A(\u_cpu.REG_FILE.rf[27][20] ),
    .B_N(\u_cpu.REG_FILE._03065_ ),
    .X(\u_cpu.REG_FILE._03893_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08612_  (.A1(\u_cpu.REG_FILE.rf[26][20] ),
    .A2(\u_cpu.REG_FILE._02772_ ),
    .B1(\u_cpu.REG_FILE._03064_ ),
    .C1(\u_cpu.REG_FILE._03893_ ),
    .Y(\u_cpu.REG_FILE._03894_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._08613_  (.A1(\u_cpu.REG_FILE._03709_ ),
    .A2(\u_cpu.REG_FILE._03891_ ),
    .A3(\u_cpu.REG_FILE._03892_ ),
    .B1(\u_cpu.REG_FILE._03800_ ),
    .C1(\u_cpu.REG_FILE._03894_ ),
    .Y(\u_cpu.REG_FILE._03895_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08614_  (.A_N(\u_cpu.REG_FILE.rf[29][20] ),
    .B(\u_cpu.REG_FILE._02768_ ),
    .X(\u_cpu.REG_FILE._03896_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08615_  (.A1(\u_cpu.REG_FILE.rf[28][20] ),
    .A2(\u_cpu.REG_FILE._03071_ ),
    .B1_N(\u_cpu.REG_FILE._03072_ ),
    .Y(\u_cpu.REG_FILE._03897_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08616_  (.A(\u_cpu.REG_FILE.rf[31][20] ),
    .B_N(\u_cpu.REG_FILE._03034_ ),
    .X(\u_cpu.REG_FILE._03898_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08617_  (.A1(\u_cpu.REG_FILE.rf[30][20] ),
    .A2(\u_cpu.REG_FILE._03075_ ),
    .B1(\u_cpu.REG_FILE._03076_ ),
    .C1(\u_cpu.REG_FILE._03898_ ),
    .Y(\u_cpu.REG_FILE._03899_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08618_  (.A1(\u_cpu.REG_FILE._03896_ ),
    .A2(\u_cpu.REG_FILE._03897_ ),
    .B1(\u_cpu.REG_FILE._03221_ ),
    .C1(\u_cpu.REG_FILE._03899_ ),
    .Y(\u_cpu.REG_FILE._03900_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._08619_  (.A1(\u_cpu.REG_FILE._03895_ ),
    .A2(\u_cpu.REG_FILE._02992_ ),
    .A3(\u_cpu.REG_FILE._03900_ ),
    .B1(\u_cpu.REG_FILE._02996_ ),
    .X(\u_cpu.REG_FILE._03901_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08620_  (.A(\u_cpu.REG_FILE.rf[8][20] ),
    .B(\u_cpu.REG_FILE._02998_ ),
    .Y(\u_cpu.REG_FILE._03902_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08621_  (.A1(\u_cpu.REG_FILE.rf[9][20] ),
    .A2(\u_cpu.REG_FILE._03132_ ),
    .B1_N(\u_cpu.REG_FILE._03133_ ),
    .Y(\u_cpu.REG_FILE._03903_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._08622_  (.A(\u_cpu.REG_FILE.rf[10][20] ),
    .B(\u_cpu.REG_FILE._02867_ ),
    .X(\u_cpu.REG_FILE._03904_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08623_  (.A1(\u_cpu.REG_FILE.rf[11][20] ),
    .A2(\u_cpu.REG_FILE._03136_ ),
    .B1(\u_cpu.REG_FILE._03137_ ),
    .C1(\u_cpu.REG_FILE._03904_ ),
    .Y(\u_cpu.REG_FILE._03905_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08624_  (.A1(\u_cpu.REG_FILE._03902_ ),
    .A2(\u_cpu.REG_FILE._03903_ ),
    .B1(\u_cpu.REG_FILE._03135_ ),
    .C1(\u_cpu.REG_FILE._03905_ ),
    .Y(\u_cpu.REG_FILE._03906_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._08625_  (.A(\u_cpu.REG_FILE.rf[14][20] ),
    .B(\u_cpu.REG_FILE._03143_ ),
    .X(\u_cpu.REG_FILE._03907_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08626_  (.A1(\u_cpu.REG_FILE.rf[15][20] ),
    .A2(\u_cpu.REG_FILE._03142_ ),
    .B1(\u_cpu.REG_FILE._03255_ ),
    .C1(\u_cpu.REG_FILE._03907_ ),
    .Y(\u_cpu.REG_FILE._03908_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08627_  (.A1(\u_cpu.REG_FILE.rf[12][20] ),
    .A2(\u_cpu.REG_FILE._03016_ ),
    .B1_N(\u_cpu.REG_FILE._02931_ ),
    .X(\u_cpu.REG_FILE._03909_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08628_  (.A1(\u_cpu.REG_FILE.rf[13][20] ),
    .A2(\u_cpu.REG_FILE._03015_ ),
    .B1(\u_cpu.REG_FILE._03909_ ),
    .Y(\u_cpu.REG_FILE._03910_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08629_  (.A(\u_cpu.REG_FILE._03908_ ),
    .B(\u_cpu.REG_FILE._03910_ ),
    .C(\u_cpu.REG_FILE._03074_ ),
    .Y(\u_cpu.REG_FILE._03911_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08630_  (.A(\u_cpu.REG_FILE._03906_ ),
    .B(\u_cpu.REG_FILE._03141_ ),
    .C(\u_cpu.REG_FILE._03911_ ),
    .Y(\u_cpu.REG_FILE._03912_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08631_  (.A(\u_cpu.REG_FILE.rf[3][20] ),
    .B_N(\u_cpu.REG_FILE._02815_ ),
    .X(\u_cpu.REG_FILE._03913_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08632_  (.A1(\u_cpu.REG_FILE.rf[2][20] ),
    .A2(\u_cpu.REG_FILE._03010_ ),
    .B1(\u_cpu.REG_FILE._03011_ ),
    .C1(\u_cpu.REG_FILE._03913_ ),
    .Y(\u_cpu.REG_FILE._03914_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08633_  (.A1(\u_cpu.REG_FILE.rf[0][20] ),
    .A2(\u_cpu.REG_FILE._03030_ ),
    .B1_N(\u_cpu.REG_FILE._02872_ ),
    .X(\u_cpu.REG_FILE._03915_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08634_  (.A1(\u_cpu.REG_FILE.rf[1][20] ),
    .A2(\u_cpu.REG_FILE._03029_ ),
    .B1(\u_cpu.REG_FILE._03915_ ),
    .Y(\u_cpu.REG_FILE._03916_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08635_  (.A(\u_cpu.REG_FILE._03009_ ),
    .B(\u_cpu.REG_FILE._03914_ ),
    .C(\u_cpu.REG_FILE._03916_ ),
    .Y(\u_cpu.REG_FILE._03917_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08636_  (.A(\u_cpu.REG_FILE.rf[7][20] ),
    .B_N(\u_cpu.REG_FILE._02783_ ),
    .X(\u_cpu.REG_FILE._03918_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08637_  (.A1(\u_cpu.REG_FILE.rf[6][20] ),
    .A2(\u_cpu.REG_FILE._02843_ ),
    .B1(\u_cpu.REG_FILE._02866_ ),
    .C1(\u_cpu.REG_FILE._03918_ ),
    .Y(\u_cpu.REG_FILE._03919_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08638_  (.A1(\u_cpu.REG_FILE.rf[4][20] ),
    .A2(\u_cpu.REG_FILE._03030_ ),
    .B1_N(\u_cpu.REG_FILE._02872_ ),
    .X(\u_cpu.REG_FILE._03920_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08639_  (.A1(\u_cpu.REG_FILE.rf[5][20] ),
    .A2(\u_cpu.REG_FILE._03029_ ),
    .B1(\u_cpu.REG_FILE._03920_ ),
    .Y(\u_cpu.REG_FILE._03921_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08640_  (.A(\u_cpu.REG_FILE._03919_ ),
    .B(\u_cpu.REG_FILE._03921_ ),
    .C(\u_cpu.REG_FILE._03042_ ),
    .Y(\u_cpu.REG_FILE._03922_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08641_  (.A(\u_cpu.REG_FILE._02851_ ),
    .B(\u_cpu.REG_FILE._03917_ ),
    .C(\u_cpu.REG_FILE._03922_ ),
    .Y(\u_cpu.REG_FILE._03923_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08642_  (.A(\u_cpu.REG_FILE._02997_ ),
    .B(\u_cpu.REG_FILE._03912_ ),
    .C(\u_cpu.REG_FILE._03923_ ),
    .Y(\u_cpu.REG_FILE._03924_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._08643_  (.A(\u_cpu.REG_FILE._02883_ ),
    .X(\u_cpu.REG_FILE._03925_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08644_  (.A1(\u_cpu.REG_FILE._03890_ ),
    .A2(\u_cpu.REG_FILE._03901_ ),
    .B1(\u_cpu.REG_FILE._03924_ ),
    .C1(\u_cpu.REG_FILE._03925_ ),
    .X(\u_cpu.ALU.SrcB[20] ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08645_  (.A1(\u_cpu.REG_FILE.rf[18][21] ),
    .A2(\u_cpu.REG_FILE._03653_ ),
    .B1(\u_cpu.REG_FILE._03298_ ),
    .Y(\u_cpu.REG_FILE._03926_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._08646_  (.A1(\u_cpu.REG_FILE._02250_ ),
    .A2(\u_cpu.REG_FILE._02939_ ),
    .B1(\u_cpu.REG_FILE._03926_ ),
    .Y(\u_cpu.REG_FILE._03927_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08647_  (.A(\u_cpu.REG_FILE.rf[16][21] ),
    .B(\u_cpu.REG_FILE._03371_ ),
    .Y(\u_cpu.REG_FILE._03928_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._08648_  (.A1(\u_cpu.REG_FILE._02253_ ),
    .A2(\u_cpu.REG_FILE._03166_ ),
    .B1(\u_cpu.REG_FILE._03057_ ),
    .C1(\u_cpu.REG_FILE._03928_ ),
    .Y(\u_cpu.REG_FILE._03929_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08649_  (.A(\u_cpu.REG_FILE.rf[20][21] ),
    .B(\u_cpu.REG_FILE._02816_ ),
    .Y(\u_cpu.REG_FILE._03930_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08650_  (.A_N(\u_cpu.REG_FILE.rf[21][21] ),
    .B(\u_cpu.REG_FILE._02801_ ),
    .X(\u_cpu.REG_FILE._03931_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08651_  (.A(\u_cpu.REG_FILE.rf[23][21] ),
    .B_N(\u_cpu.REG_FILE._02771_ ),
    .X(\u_cpu.REG_FILE._03932_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08652_  (.A1(\u_cpu.REG_FILE.rf[22][21] ),
    .A2(\u_cpu.REG_FILE._02816_ ),
    .B1(\u_cpu.REG_FILE._02818_ ),
    .C1(\u_cpu.REG_FILE._03932_ ),
    .Y(\u_cpu.REG_FILE._03933_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._08653_  (.A1(\u_cpu.REG_FILE._03709_ ),
    .A2(\u_cpu.REG_FILE._03930_ ),
    .A3(\u_cpu.REG_FILE._03931_ ),
    .B1(\u_cpu.REG_FILE._02804_ ),
    .C1(\u_cpu.REG_FILE._03933_ ),
    .Y(\u_cpu.REG_FILE._03934_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.REG_FILE._08654_  (.A1(\u_cpu.REG_FILE._02765_ ),
    .A2(\u_cpu.REG_FILE._03927_ ),
    .A3(\u_cpu.REG_FILE._03929_ ),
    .B1(\u_cpu.REG_FILE._03934_ ),
    .C1(\u_cpu.REG_FILE._02966_ ),
    .X(\u_cpu.REG_FILE._03935_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08655_  (.A(\u_cpu.REG_FILE.rf[24][21] ),
    .B(\u_cpu.REG_FILE._03058_ ),
    .Y(\u_cpu.REG_FILE._03936_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08656_  (.A_N(\u_cpu.REG_FILE.rf[25][21] ),
    .B(\u_cpu.REG_FILE._03060_ ),
    .X(\u_cpu.REG_FILE._03937_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08657_  (.A(\u_cpu.REG_FILE.rf[27][21] ),
    .B_N(\u_cpu.REG_FILE._03065_ ),
    .X(\u_cpu.REG_FILE._03938_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08658_  (.A1(\u_cpu.REG_FILE.rf[26][21] ),
    .A2(\u_cpu.REG_FILE._02772_ ),
    .B1(\u_cpu.REG_FILE._03064_ ),
    .C1(\u_cpu.REG_FILE._03938_ ),
    .Y(\u_cpu.REG_FILE._03939_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._08659_  (.A1(\u_cpu.REG_FILE._03709_ ),
    .A2(\u_cpu.REG_FILE._03936_ ),
    .A3(\u_cpu.REG_FILE._03937_ ),
    .B1(\u_cpu.REG_FILE._03800_ ),
    .C1(\u_cpu.REG_FILE._03939_ ),
    .Y(\u_cpu.REG_FILE._03940_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08660_  (.A_N(\u_cpu.REG_FILE.rf[29][21] ),
    .B(\u_cpu.REG_FILE._02768_ ),
    .X(\u_cpu.REG_FILE._03941_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08661_  (.A1(\u_cpu.REG_FILE.rf[28][21] ),
    .A2(\u_cpu.REG_FILE._03071_ ),
    .B1_N(\u_cpu.REG_FILE._03072_ ),
    .Y(\u_cpu.REG_FILE._03942_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08662_  (.A(\u_cpu.REG_FILE.rf[31][21] ),
    .B_N(\u_cpu.REG_FILE._03034_ ),
    .X(\u_cpu.REG_FILE._03943_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08663_  (.A1(\u_cpu.REG_FILE.rf[30][21] ),
    .A2(\u_cpu.REG_FILE._03075_ ),
    .B1(\u_cpu.REG_FILE._03076_ ),
    .C1(\u_cpu.REG_FILE._03943_ ),
    .Y(\u_cpu.REG_FILE._03944_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08664_  (.A1(\u_cpu.REG_FILE._03941_ ),
    .A2(\u_cpu.REG_FILE._03942_ ),
    .B1(\u_cpu.REG_FILE._03221_ ),
    .C1(\u_cpu.REG_FILE._03944_ ),
    .Y(\u_cpu.REG_FILE._03945_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._08665_  (.A1(\u_cpu.REG_FILE._03940_ ),
    .A2(\u_cpu.REG_FILE._02992_ ),
    .A3(\u_cpu.REG_FILE._03945_ ),
    .B1(\u_cpu.REG_FILE._02996_ ),
    .X(\u_cpu.REG_FILE._03946_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08666_  (.A(\u_cpu.REG_FILE.rf[12][21] ),
    .B(\u_cpu.REG_FILE._02950_ ),
    .Y(\u_cpu.REG_FILE._03947_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08667_  (.A1(\u_cpu.REG_FILE.rf[13][21] ),
    .A2(\u_cpu.REG_FILE._03132_ ),
    .B1_N(\u_cpu.REG_FILE._03133_ ),
    .Y(\u_cpu.REG_FILE._03948_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._08668_  (.A(\u_cpu.REG_FILE.rf[14][21] ),
    .B(\u_cpu.REG_FILE._02867_ ),
    .X(\u_cpu.REG_FILE._03949_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08669_  (.A1(\u_cpu.REG_FILE.rf[15][21] ),
    .A2(\u_cpu.REG_FILE._03136_ ),
    .B1(\u_cpu.REG_FILE._03076_ ),
    .C1(\u_cpu.REG_FILE._03949_ ),
    .Y(\u_cpu.REG_FILE._03950_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08670_  (.A1(\u_cpu.REG_FILE._03947_ ),
    .A2(\u_cpu.REG_FILE._03948_ ),
    .B1(\u_cpu.REG_FILE._03042_ ),
    .C1(\u_cpu.REG_FILE._03950_ ),
    .Y(\u_cpu.REG_FILE._03951_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08671_  (.A(\u_cpu.REG_FILE.rf[11][21] ),
    .B_N(\u_cpu.REG_FILE._03012_ ),
    .X(\u_cpu.REG_FILE._03952_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08672_  (.A1(\u_cpu.REG_FILE.rf[10][21] ),
    .A2(\u_cpu.REG_FILE._03010_ ),
    .B1(\u_cpu.REG_FILE._03011_ ),
    .C1(\u_cpu.REG_FILE._03952_ ),
    .Y(\u_cpu.REG_FILE._03953_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08673_  (.A1(\u_cpu.REG_FILE.rf[8][21] ),
    .A2(\u_cpu.REG_FILE._03090_ ),
    .B1_N(\u_cpu.REG_FILE._03017_ ),
    .X(\u_cpu.REG_FILE._03954_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08674_  (.A1(\u_cpu.REG_FILE.rf[9][21] ),
    .A2(\u_cpu.REG_FILE._03136_ ),
    .B1(\u_cpu.REG_FILE._03954_ ),
    .Y(\u_cpu.REG_FILE._03955_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08675_  (.A(\u_cpu.REG_FILE._03135_ ),
    .B(\u_cpu.REG_FILE._03953_ ),
    .C(\u_cpu.REG_FILE._03955_ ),
    .Y(\u_cpu.REG_FILE._03956_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08676_  (.A(\u_cpu.REG_FILE._03951_ ),
    .B(\u_cpu.REG_FILE._03956_ ),
    .C(\u_cpu.REG_FILE._03021_ ),
    .Y(\u_cpu.REG_FILE._03957_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08677_  (.A(\u_cpu.REG_FILE.rf[3][21] ),
    .B_N(\u_cpu.REG_FILE._02815_ ),
    .X(\u_cpu.REG_FILE._03958_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08678_  (.A1(\u_cpu.REG_FILE.rf[2][21] ),
    .A2(\u_cpu.REG_FILE._03010_ ),
    .B1(\u_cpu.REG_FILE._03011_ ),
    .C1(\u_cpu.REG_FILE._03958_ ),
    .Y(\u_cpu.REG_FILE._03959_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08679_  (.A1(\u_cpu.REG_FILE.rf[0][21] ),
    .A2(\u_cpu.REG_FILE._02827_ ),
    .B1_N(\u_cpu.REG_FILE._02872_ ),
    .X(\u_cpu.REG_FILE._03960_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08680_  (.A1(\u_cpu.REG_FILE.rf[1][21] ),
    .A2(\u_cpu.REG_FILE._03029_ ),
    .B1(\u_cpu.REG_FILE._03960_ ),
    .Y(\u_cpu.REG_FILE._03961_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08681_  (.A(\u_cpu.REG_FILE._03009_ ),
    .B(\u_cpu.REG_FILE._03959_ ),
    .C(\u_cpu.REG_FILE._03961_ ),
    .Y(\u_cpu.REG_FILE._03962_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08682_  (.A(\u_cpu.REG_FILE.rf[4][21] ),
    .B(\u_cpu.REG_FILE._03404_ ),
    .Y(\u_cpu.REG_FILE._03963_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08683_  (.A_N(\u_cpu.REG_FILE.rf[5][21] ),
    .B(\u_cpu.REG_FILE._02748_ ),
    .X(\u_cpu.REG_FILE._03964_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.REG_FILE._08684_  (.A1(\u_cpu.REG_FILE.rf[6][21] ),
    .A2(\u_cpu.REG_FILE._02779_ ),
    .B1(\u_cpu.REG_FILE._02781_ ),
    .X(\u_cpu.REG_FILE._03965_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08685_  (.A1(\u_cpu.REG_FILE.rf[7][21] ),
    .A2(\u_cpu.REG_FILE._03351_ ),
    .B1(\u_cpu.REG_FILE._03965_ ),
    .Y(\u_cpu.REG_FILE._03966_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._08686_  (.A1(\u_cpu.REG_FILE._03403_ ),
    .A2(\u_cpu.REG_FILE._03963_ ),
    .A3(\u_cpu.REG_FILE._03964_ ),
    .B1(\u_cpu.REG_FILE._02834_ ),
    .C1(\u_cpu.REG_FILE._03966_ ),
    .Y(\u_cpu.REG_FILE._03967_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08687_  (.A(\u_cpu.REG_FILE._02851_ ),
    .B(\u_cpu.REG_FILE._03962_ ),
    .C(\u_cpu.REG_FILE._03967_ ),
    .Y(\u_cpu.REG_FILE._03968_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08688_  (.A(\u_cpu.REG_FILE._02994_ ),
    .B(\u_cpu.REG_FILE._03957_ ),
    .C(\u_cpu.REG_FILE._03968_ ),
    .Y(\u_cpu.REG_FILE._03969_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08689_  (.A1(\u_cpu.REG_FILE._03935_ ),
    .A2(\u_cpu.REG_FILE._03946_ ),
    .B1(\u_cpu.REG_FILE._03969_ ),
    .C1(\u_cpu.REG_FILE._03925_ ),
    .X(\u_cpu.ALU.SrcB[21] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08690_  (.A(\u_cpu.REG_FILE.rf[11][22] ),
    .B_N(\u_cpu.REG_FILE._03311_ ),
    .X(\u_cpu.REG_FILE._03970_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08691_  (.A1(\u_cpu.REG_FILE.rf[10][22] ),
    .A2(\u_cpu.REG_FILE._02950_ ),
    .B1(\u_cpu.REG_FILE._02826_ ),
    .C1(\u_cpu.REG_FILE._03970_ ),
    .X(\u_cpu.REG_FILE._03971_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08692_  (.A1(\u_cpu.REG_FILE.rf[8][22] ),
    .A2(\u_cpu.REG_FILE._02760_ ),
    .B1_N(\u_cpu.REG_FILE._02825_ ),
    .X(\u_cpu.REG_FILE._03972_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08693_  (.A(\u_cpu.REG_FILE.rf[9][22] ),
    .B_N(\u_cpu.REG_FILE._02832_ ),
    .X(\u_cpu.REG_FILE._03973_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._08694_  (.A1(\u_cpu.REG_FILE._03972_ ),
    .A2(\u_cpu.REG_FILE._03973_ ),
    .B1(\u_cpu.REG_FILE._02834_ ),
    .X(\u_cpu.REG_FILE._03974_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08695_  (.A(\u_cpu.REG_FILE.rf[14][22] ),
    .B(\u_cpu.REG_FILE._02968_ ),
    .Y(\u_cpu.REG_FILE._03975_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08696_  (.A1(\u_cpu.REG_FILE.rf[15][22] ),
    .A2(\u_cpu.REG_FILE._03002_ ),
    .B1(\u_cpu.REG_FILE._02826_ ),
    .Y(\u_cpu.REG_FILE._03976_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08697_  (.A1(\u_cpu.REG_FILE.rf[12][22] ),
    .A2(\u_cpu.REG_FILE._03445_ ),
    .B1_N(\u_cpu.REG_FILE._02825_ ),
    .X(\u_cpu.REG_FILE._03977_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08698_  (.A1(\u_cpu.REG_FILE.rf[13][22] ),
    .A2(\u_cpu.REG_FILE._03002_ ),
    .B1(\u_cpu.REG_FILE._03977_ ),
    .Y(\u_cpu.REG_FILE._03978_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08699_  (.A1(\u_cpu.REG_FILE._03975_ ),
    .A2(\u_cpu.REG_FILE._03976_ ),
    .B1(\u_cpu.REG_FILE._03978_ ),
    .C1(\u_cpu.REG_FILE._02765_ ),
    .Y(\u_cpu.REG_FILE._03979_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08700_  (.A1(\u_cpu.REG_FILE._03971_ ),
    .A2(\u_cpu.REG_FILE._03974_ ),
    .B1(\u_cpu.REG_FILE._03218_ ),
    .C1(\u_cpu.REG_FILE._03979_ ),
    .X(\u_cpu.REG_FILE._03980_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08701_  (.A_N(\u_cpu.REG_FILE.rf[1][22] ),
    .B(\u_cpu.REG_FILE._02980_ ),
    .X(\u_cpu.REG_FILE._03981_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08702_  (.A1(\u_cpu.REG_FILE.rf[0][22] ),
    .A2(\u_cpu.REG_FILE._03212_ ),
    .B1_N(\u_cpu.REG_FILE._02983_ ),
    .Y(\u_cpu.REG_FILE._03982_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08703_  (.A(\u_cpu.REG_FILE.rf[3][22] ),
    .B_N(\u_cpu.REG_FILE._03077_ ),
    .X(\u_cpu.REG_FILE._03983_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08704_  (.A1(\u_cpu.REG_FILE.rf[2][22] ),
    .A2(\u_cpu.REG_FILE._03125_ ),
    .B1(\u_cpu.REG_FILE._02988_ ),
    .C1(\u_cpu.REG_FILE._03983_ ),
    .Y(\u_cpu.REG_FILE._03984_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08705_  (.A1(\u_cpu.REG_FILE._03981_ ),
    .A2(\u_cpu.REG_FILE._03982_ ),
    .B1(\u_cpu.REG_FILE._02777_ ),
    .C1(\u_cpu.REG_FILE._03984_ ),
    .Y(\u_cpu.REG_FILE._03985_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08706_  (.A_N(\u_cpu.REG_FILE.rf[5][22] ),
    .B(\u_cpu.REG_FILE._02768_ ),
    .X(\u_cpu.REG_FILE._03986_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08707_  (.A1(\u_cpu.REG_FILE.rf[4][22] ),
    .A2(\u_cpu.REG_FILE._03071_ ),
    .B1_N(\u_cpu.REG_FILE._02774_ ),
    .Y(\u_cpu.REG_FILE._03987_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08708_  (.A(\u_cpu.REG_FILE.rf[7][22] ),
    .B_N(\u_cpu.REG_FILE._03034_ ),
    .X(\u_cpu.REG_FILE._03988_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08709_  (.A1(\u_cpu.REG_FILE.rf[6][22] ),
    .A2(\u_cpu.REG_FILE._03075_ ),
    .B1(\u_cpu.REG_FILE._03076_ ),
    .C1(\u_cpu.REG_FILE._03988_ ),
    .Y(\u_cpu.REG_FILE._03989_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08710_  (.A1(\u_cpu.REG_FILE._03986_ ),
    .A2(\u_cpu.REG_FILE._03987_ ),
    .B1(\u_cpu.REG_FILE._03221_ ),
    .C1(\u_cpu.REG_FILE._03989_ ),
    .Y(\u_cpu.REG_FILE._03990_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._08711_  (.A1(\u_cpu.REG_FILE._02807_ ),
    .A2(\u_cpu.REG_FILE._03985_ ),
    .A3(\u_cpu.REG_FILE._03990_ ),
    .B1(\u_cpu.REG_FILE._02745_ ),
    .X(\u_cpu.REG_FILE._03991_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08712_  (.A(\u_cpu.REG_FILE.rf[27][22] ),
    .B_N(\u_cpu.REG_FILE._02871_ ),
    .X(\u_cpu.REG_FILE._03992_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08713_  (.A1(\u_cpu.REG_FILE.rf[26][22] ),
    .A2(\u_cpu.REG_FILE._02982_ ),
    .B1(\u_cpu.REG_FILE._03000_ ),
    .C1(\u_cpu.REG_FILE._03992_ ),
    .X(\u_cpu.REG_FILE._03993_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08714_  (.A(\u_cpu.REG_FILE.rf[24][22] ),
    .B(\u_cpu.REG_FILE._03287_ ),
    .Y(\u_cpu.REG_FILE._03994_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08715_  (.A_N(\u_cpu.REG_FILE.rf[25][22] ),
    .B(\u_cpu.REG_FILE._02830_ ),
    .X(\u_cpu.REG_FILE._03995_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.REG_FILE._08716_  (.A1(\u_cpu.REG_FILE._03403_ ),
    .A2(\u_cpu.REG_FILE._03994_ ),
    .A3(\u_cpu.REG_FILE._03995_ ),
    .B1(\u_cpu.REG_FILE._03800_ ),
    .Y(\u_cpu.REG_FILE._03996_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08717_  (.A(\u_cpu.REG_FILE.rf[30][22] ),
    .B(\u_cpu.REG_FILE._03063_ ),
    .Y(\u_cpu.REG_FILE._03997_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08718_  (.A1(\u_cpu.REG_FILE.rf[31][22] ),
    .A2(\u_cpu.REG_FILE._03297_ ),
    .B1(\u_cpu.REG_FILE._02854_ ),
    .Y(\u_cpu.REG_FILE._03998_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08719_  (.A(\u_cpu.REG_FILE.rf[28][22] ),
    .B(\u_cpu.REG_FILE._02916_ ),
    .Y(\u_cpu.REG_FILE._03999_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08720_  (.A1(\u_cpu.REG_FILE.rf[29][22] ),
    .A2(\u_cpu.REG_FILE._03351_ ),
    .B1_N(\u_cpu.REG_FILE._02947_ ),
    .Y(\u_cpu.REG_FILE._04000_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._08721_  (.A1(\u_cpu.REG_FILE._03997_ ),
    .A2(\u_cpu.REG_FILE._03998_ ),
    .B1(\u_cpu.REG_FILE._03999_ ),
    .B2(\u_cpu.REG_FILE._04000_ ),
    .C1(\u_cpu.REG_FILE._02919_ ),
    .Y(\u_cpu.REG_FILE._04001_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08722_  (.A1(\u_cpu.REG_FILE._03993_ ),
    .A2(\u_cpu.REG_FILE._03996_ ),
    .B1(\u_cpu.REG_FILE._02836_ ),
    .C1(\u_cpu.REG_FILE._04001_ ),
    .Y(\u_cpu.REG_FILE._04002_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08723_  (.A1(\u_cpu.REG_FILE.rf[18][22] ),
    .A2(\u_cpu.REG_FILE._02923_ ),
    .B1(\u_cpu.REG_FILE._03249_ ),
    .Y(\u_cpu.REG_FILE._04003_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08724_  (.A(\u_cpu.REG_FILE.rf[19][22] ),
    .B(\u_cpu.REG_FILE._02856_ ),
    .Y(\u_cpu.REG_FILE._04004_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08725_  (.A1(\u_cpu.REG_FILE.rf[16][22] ),
    .A2(\u_cpu.REG_FILE._03038_ ),
    .B1_N(\u_cpu.REG_FILE._03039_ ),
    .X(\u_cpu.REG_FILE._04005_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08726_  (.A1(\u_cpu.REG_FILE.rf[17][22] ),
    .A2(\u_cpu.REG_FILE._03304_ ),
    .B1(\u_cpu.REG_FILE._04005_ ),
    .Y(\u_cpu.REG_FILE._04006_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08727_  (.A1(\u_cpu.REG_FILE._04003_ ),
    .A2(\u_cpu.REG_FILE._04004_ ),
    .B1(\u_cpu.REG_FILE._03292_ ),
    .C1(\u_cpu.REG_FILE._04006_ ),
    .Y(\u_cpu.REG_FILE._04007_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._08728_  (.A(\u_cpu.REG_FILE.rf[22][22] ),
    .B(\u_cpu.REG_FILE._03143_ ),
    .X(\u_cpu.REG_FILE._04008_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08729_  (.A1(\u_cpu.REG_FILE.rf[23][22] ),
    .A2(\u_cpu.REG_FILE._03142_ ),
    .B1(\u_cpu.REG_FILE._03255_ ),
    .C1(\u_cpu.REG_FILE._04008_ ),
    .Y(\u_cpu.REG_FILE._04009_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08730_  (.A1(\u_cpu.REG_FILE.rf[20][22] ),
    .A2(\u_cpu.REG_FILE._03016_ ),
    .B1_N(\u_cpu.REG_FILE._03017_ ),
    .X(\u_cpu.REG_FILE._04010_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08731_  (.A1(\u_cpu.REG_FILE.rf[21][22] ),
    .A2(\u_cpu.REG_FILE._03015_ ),
    .B1(\u_cpu.REG_FILE._04010_ ),
    .Y(\u_cpu.REG_FILE._04011_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08732_  (.A(\u_cpu.REG_FILE._04009_ ),
    .B(\u_cpu.REG_FILE._04011_ ),
    .C(\u_cpu.REG_FILE._03074_ ),
    .Y(\u_cpu.REG_FILE._04012_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08733_  (.A(\u_cpu.REG_FILE._02922_ ),
    .B(\u_cpu.REG_FILE._04007_ ),
    .C(\u_cpu.REG_FILE._04012_ ),
    .Y(\u_cpu.REG_FILE._04013_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08734_  (.A(\u_cpu.REG_FILE._04002_ ),
    .B(\u_cpu.REG_FILE._04013_ ),
    .C(\u_cpu.REG_FILE._02745_ ),
    .Y(\u_cpu.REG_FILE._04014_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08735_  (.A1(\u_cpu.REG_FILE._03980_ ),
    .A2(\u_cpu.REG_FILE._03991_ ),
    .B1(\u_cpu.REG_FILE._04014_ ),
    .C1(\u_cpu.REG_FILE._03925_ ),
    .X(\u_cpu.ALU.SrcB[22] ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08736_  (.A1(\u_cpu.REG_FILE.rf[16][23] ),
    .A2(\u_cpu.REG_FILE._02790_ ),
    .B1_N(\u_cpu.REG_FILE._02751_ ),
    .Y(\u_cpu.REG_FILE._04015_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08737_  (.A_N(\u_cpu.REG_FILE.rf[17][23] ),
    .B(\u_cpu.REG_FILE._03445_ ),
    .X(\u_cpu.REG_FILE._04016_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08738_  (.A1(\u_cpu.REG_FILE.rf[18][23] ),
    .A2(\u_cpu.REG_FILE._03404_ ),
    .B1(\u_cpu.REG_FILE._03470_ ),
    .Y(\u_cpu.REG_FILE._04017_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08739_  (.A_N(\u_cpu.REG_FILE.rf[19][23] ),
    .B(\u_cpu.REG_FILE._02980_ ),
    .X(\u_cpu.REG_FILE._04018_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu.REG_FILE._08740_  (.A1(\u_cpu.REG_FILE._04015_ ),
    .A2(\u_cpu.REG_FILE._04016_ ),
    .B1(\u_cpu.REG_FILE._04017_ ),
    .B2(\u_cpu.REG_FILE._04018_ ),
    .Y(\u_cpu.REG_FILE._04019_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08741_  (.A(\u_cpu.REG_FILE.rf[23][23] ),
    .B_N(\u_cpu.REG_FILE._03003_ ),
    .X(\u_cpu.REG_FILE._04020_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08742_  (.A1(\u_cpu.REG_FILE.rf[22][23] ),
    .A2(\u_cpu.REG_FILE._02987_ ),
    .B1(\u_cpu.REG_FILE._02826_ ),
    .C1(\u_cpu.REG_FILE._04020_ ),
    .X(\u_cpu.REG_FILE._04021_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08743_  (.A(\u_cpu.REG_FILE.rf[20][23] ),
    .B(\u_cpu.REG_FILE._02940_ ),
    .Y(\u_cpu.REG_FILE._04022_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08744_  (.A_N(\u_cpu.REG_FILE.rf[21][23] ),
    .B(\u_cpu.REG_FILE._02880_ ),
    .X(\u_cpu.REG_FILE._04023_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu.REG_FILE._08745_  (.A1(\u_cpu.REG_FILE._03403_ ),
    .A2(\u_cpu.REG_FILE._04022_ ),
    .A3(\u_cpu.REG_FILE._04023_ ),
    .B1(\u_cpu.REG_FILE._02804_ ),
    .Y(\u_cpu.REG_FILE._04024_ ));
 sky130_fd_sc_hd__o221a_2 \u_cpu.REG_FILE._08746_  (.A1(\u_cpu.REG_FILE._02937_ ),
    .A2(\u_cpu.REG_FILE._04019_ ),
    .B1(\u_cpu.REG_FILE._04021_ ),
    .B2(\u_cpu.REG_FILE._04024_ ),
    .C1(\u_cpu.REG_FILE._03023_ ),
    .X(\u_cpu.REG_FILE._04025_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08747_  (.A(\u_cpu.REG_FILE.rf[24][23] ),
    .B(\u_cpu.REG_FILE._03058_ ),
    .Y(\u_cpu.REG_FILE._04026_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08748_  (.A_N(\u_cpu.REG_FILE.rf[25][23] ),
    .B(\u_cpu.REG_FILE._03060_ ),
    .X(\u_cpu.REG_FILE._04027_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08749_  (.A(\u_cpu.REG_FILE.rf[27][23] ),
    .B_N(\u_cpu.REG_FILE._03065_ ),
    .X(\u_cpu.REG_FILE._04028_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08750_  (.A1(\u_cpu.REG_FILE.rf[26][23] ),
    .A2(\u_cpu.REG_FILE._02772_ ),
    .B1(\u_cpu.REG_FILE._03064_ ),
    .C1(\u_cpu.REG_FILE._04028_ ),
    .Y(\u_cpu.REG_FILE._04029_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._08751_  (.A1(\u_cpu.REG_FILE._03709_ ),
    .A2(\u_cpu.REG_FILE._04026_ ),
    .A3(\u_cpu.REG_FILE._04027_ ),
    .B1(\u_cpu.REG_FILE._03800_ ),
    .C1(\u_cpu.REG_FILE._04029_ ),
    .Y(\u_cpu.REG_FILE._04030_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08752_  (.A_N(\u_cpu.REG_FILE.rf[29][23] ),
    .B(\u_cpu.REG_FILE._02768_ ),
    .X(\u_cpu.REG_FILE._04031_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08753_  (.A1(\u_cpu.REG_FILE.rf[28][23] ),
    .A2(\u_cpu.REG_FILE._03071_ ),
    .B1_N(\u_cpu.REG_FILE._02774_ ),
    .Y(\u_cpu.REG_FILE._04032_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08754_  (.A(\u_cpu.REG_FILE.rf[31][23] ),
    .B_N(\u_cpu.REG_FILE._03034_ ),
    .X(\u_cpu.REG_FILE._04033_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08755_  (.A1(\u_cpu.REG_FILE.rf[30][23] ),
    .A2(\u_cpu.REG_FILE._02843_ ),
    .B1(\u_cpu.REG_FILE._03076_ ),
    .C1(\u_cpu.REG_FILE._04033_ ),
    .Y(\u_cpu.REG_FILE._04034_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08756_  (.A1(\u_cpu.REG_FILE._04031_ ),
    .A2(\u_cpu.REG_FILE._04032_ ),
    .B1(\u_cpu.REG_FILE._03221_ ),
    .C1(\u_cpu.REG_FILE._04034_ ),
    .Y(\u_cpu.REG_FILE._04035_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._08757_  (.A1(\u_cpu.REG_FILE._04030_ ),
    .A2(\u_cpu.REG_FILE._02992_ ),
    .A3(\u_cpu.REG_FILE._04035_ ),
    .B1(\u_cpu.REG_FILE._02996_ ),
    .X(\u_cpu.REG_FILE._04036_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08758_  (.A(\u_cpu.REG_FILE.rf[14][23] ),
    .B(\u_cpu.REG_FILE._02950_ ),
    .Y(\u_cpu.REG_FILE._04037_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08759_  (.A1(\u_cpu.REG_FILE.rf[15][23] ),
    .A2(\u_cpu.REG_FILE._02960_ ),
    .B1(\u_cpu.REG_FILE._02961_ ),
    .Y(\u_cpu.REG_FILE._04038_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08760_  (.A1(\u_cpu.REG_FILE.rf[12][23] ),
    .A2(\u_cpu.REG_FILE._02860_ ),
    .B1_N(\u_cpu.REG_FILE._02817_ ),
    .X(\u_cpu.REG_FILE._04039_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08761_  (.A1(\u_cpu.REG_FILE.rf[13][23] ),
    .A2(\u_cpu.REG_FILE._02956_ ),
    .B1(\u_cpu.REG_FILE._04039_ ),
    .Y(\u_cpu.REG_FILE._04040_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08762_  (.A1(\u_cpu.REG_FILE._04037_ ),
    .A2(\u_cpu.REG_FILE._04038_ ),
    .B1(\u_cpu.REG_FILE._04040_ ),
    .C1(\u_cpu.REG_FILE._02963_ ),
    .Y(\u_cpu.REG_FILE._04041_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08763_  (.A(\u_cpu.REG_FILE.rf[11][23] ),
    .B_N(\u_cpu.REG_FILE._03012_ ),
    .X(\u_cpu.REG_FILE._04042_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08764_  (.A1(\u_cpu.REG_FILE.rf[10][23] ),
    .A2(\u_cpu.REG_FILE._03010_ ),
    .B1(\u_cpu.REG_FILE._03011_ ),
    .C1(\u_cpu.REG_FILE._04042_ ),
    .Y(\u_cpu.REG_FILE._04043_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08765_  (.A1(\u_cpu.REG_FILE.rf[8][23] ),
    .A2(\u_cpu.REG_FILE._03090_ ),
    .B1_N(\u_cpu.REG_FILE._02798_ ),
    .X(\u_cpu.REG_FILE._04044_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08766_  (.A1(\u_cpu.REG_FILE.rf[9][23] ),
    .A2(\u_cpu.REG_FILE._03136_ ),
    .B1(\u_cpu.REG_FILE._04044_ ),
    .Y(\u_cpu.REG_FILE._04045_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08767_  (.A(\u_cpu.REG_FILE._03135_ ),
    .B(\u_cpu.REG_FILE._04043_ ),
    .C(\u_cpu.REG_FILE._04045_ ),
    .Y(\u_cpu.REG_FILE._04046_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08768_  (.A(\u_cpu.REG_FILE._04041_ ),
    .B(\u_cpu.REG_FILE._04046_ ),
    .C(\u_cpu.REG_FILE._03021_ ),
    .Y(\u_cpu.REG_FILE._04047_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08769_  (.A(\u_cpu.REG_FILE.rf[3][23] ),
    .B_N(\u_cpu.REG_FILE._02815_ ),
    .X(\u_cpu.REG_FILE._04048_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08770_  (.A1(\u_cpu.REG_FILE.rf[2][23] ),
    .A2(\u_cpu.REG_FILE._03010_ ),
    .B1(\u_cpu.REG_FILE._03011_ ),
    .C1(\u_cpu.REG_FILE._04048_ ),
    .Y(\u_cpu.REG_FILE._04049_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08771_  (.A1(\u_cpu.REG_FILE.rf[0][23] ),
    .A2(\u_cpu.REG_FILE._02827_ ),
    .B1_N(\u_cpu.REG_FILE._02872_ ),
    .X(\u_cpu.REG_FILE._04050_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08772_  (.A1(\u_cpu.REG_FILE.rf[1][23] ),
    .A2(\u_cpu.REG_FILE._03029_ ),
    .B1(\u_cpu.REG_FILE._04050_ ),
    .Y(\u_cpu.REG_FILE._04051_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08773_  (.A(\u_cpu.REG_FILE._03009_ ),
    .B(\u_cpu.REG_FILE._04049_ ),
    .C(\u_cpu.REG_FILE._04051_ ),
    .Y(\u_cpu.REG_FILE._04052_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08774_  (.A(\u_cpu.REG_FILE.rf[4][23] ),
    .B(\u_cpu.REG_FILE._03404_ ),
    .Y(\u_cpu.REG_FILE._04053_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08775_  (.A_N(\u_cpu.REG_FILE.rf[5][23] ),
    .B(\u_cpu.REG_FILE._02748_ ),
    .X(\u_cpu.REG_FILE._04054_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08776_  (.A(\u_cpu.REG_FILE.rf[7][23] ),
    .B_N(\u_cpu.REG_FILE._02792_ ),
    .X(\u_cpu.REG_FILE._04055_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08777_  (.A1(\u_cpu.REG_FILE.rf[6][23] ),
    .A2(\u_cpu.REG_FILE._03309_ ),
    .B1(\u_cpu.REG_FILE._03407_ ),
    .C1(\u_cpu.REG_FILE._04055_ ),
    .Y(\u_cpu.REG_FILE._04056_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._08778_  (.A1(\u_cpu.REG_FILE._03403_ ),
    .A2(\u_cpu.REG_FILE._04053_ ),
    .A3(\u_cpu.REG_FILE._04054_ ),
    .B1(\u_cpu.REG_FILE._02834_ ),
    .C1(\u_cpu.REG_FILE._04056_ ),
    .Y(\u_cpu.REG_FILE._04057_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08779_  (.A(\u_cpu.REG_FILE._02851_ ),
    .B(\u_cpu.REG_FILE._04052_ ),
    .C(\u_cpu.REG_FILE._04057_ ),
    .Y(\u_cpu.REG_FILE._04058_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08780_  (.A(\u_cpu.REG_FILE._02994_ ),
    .B(\u_cpu.REG_FILE._04047_ ),
    .C(\u_cpu.REG_FILE._04058_ ),
    .Y(\u_cpu.REG_FILE._04059_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08781_  (.A1(\u_cpu.REG_FILE._04025_ ),
    .A2(\u_cpu.REG_FILE._04036_ ),
    .B1(\u_cpu.REG_FILE._04059_ ),
    .C1(\u_cpu.REG_FILE._03925_ ),
    .X(\u_cpu.ALU.SrcB[23] ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08782_  (.A1(\u_cpu.REG_FILE.rf[18][24] ),
    .A2(\u_cpu.REG_FILE._03653_ ),
    .B1(\u_cpu.REG_FILE._03298_ ),
    .Y(\u_cpu.REG_FILE._04060_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._08783_  (.A1(\u_cpu.REG_FILE._02402_ ),
    .A2(\u_cpu.REG_FILE._02939_ ),
    .B1(\u_cpu.REG_FILE._04060_ ),
    .Y(\u_cpu.REG_FILE._04061_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08784_  (.A(\u_cpu.REG_FILE.rf[16][24] ),
    .B(\u_cpu.REG_FILE._03371_ ),
    .Y(\u_cpu.REG_FILE._04062_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._08785_  (.A1(\u_cpu.REG_FILE._02405_ ),
    .A2(\u_cpu.REG_FILE._03166_ ),
    .B1(\u_cpu.REG_FILE._03057_ ),
    .C1(\u_cpu.REG_FILE._04062_ ),
    .Y(\u_cpu.REG_FILE._04063_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08786_  (.A1(\u_cpu.REG_FILE.rf[20][24] ),
    .A2(\u_cpu.REG_FILE._02853_ ),
    .B1_N(\u_cpu.REG_FILE._03050_ ),
    .Y(\u_cpu.REG_FILE._04064_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08787_  (.A(\u_cpu.REG_FILE.rf[21][24] ),
    .B(\u_cpu.REG_FILE._02859_ ),
    .Y(\u_cpu.REG_FILE._04065_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08788_  (.A(\u_cpu.REG_FILE.rf[22][24] ),
    .B(\u_cpu.REG_FILE._02958_ ),
    .Y(\u_cpu.REG_FILE._04066_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08789_  (.A1(\u_cpu.REG_FILE.rf[23][24] ),
    .A2(\u_cpu.REG_FILE._03114_ ),
    .B1(\u_cpu.REG_FILE._03377_ ),
    .Y(\u_cpu.REG_FILE._04067_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._08790_  (.A1(\u_cpu.REG_FILE._04064_ ),
    .A2(\u_cpu.REG_FILE._04065_ ),
    .B1(\u_cpu.REG_FILE._04066_ ),
    .B2(\u_cpu.REG_FILE._04067_ ),
    .C1(\u_cpu.REG_FILE._02848_ ),
    .Y(\u_cpu.REG_FILE._04068_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.REG_FILE._08791_  (.A1(\u_cpu.REG_FILE._02765_ ),
    .A2(\u_cpu.REG_FILE._04061_ ),
    .A3(\u_cpu.REG_FILE._04063_ ),
    .B1(\u_cpu.REG_FILE._04068_ ),
    .C1(\u_cpu.REG_FILE._02966_ ),
    .X(\u_cpu.REG_FILE._04069_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08792_  (.A(\u_cpu.REG_FILE.rf[31][24] ),
    .B_N(\u_cpu.REG_FILE._02970_ ),
    .X(\u_cpu.REG_FILE._04070_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08793_  (.A1(\u_cpu.REG_FILE.rf[30][24] ),
    .A2(\u_cpu.REG_FILE._02749_ ),
    .B1(\u_cpu.REG_FILE._02969_ ),
    .C1(\u_cpu.REG_FILE._04070_ ),
    .Y(\u_cpu.REG_FILE._04071_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08794_  (.A1(\u_cpu.REG_FILE.rf[28][24] ),
    .A2(\u_cpu.REG_FILE._02830_ ),
    .B1_N(\u_cpu.REG_FILE._02975_ ),
    .X(\u_cpu.REG_FILE._04072_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08795_  (.A1(\u_cpu.REG_FILE.rf[29][24] ),
    .A2(\u_cpu.REG_FILE._02973_ ),
    .B1(\u_cpu.REG_FILE._04072_ ),
    .Y(\u_cpu.REG_FILE._04073_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08796_  (.A(\u_cpu.REG_FILE._04071_ ),
    .B(\u_cpu.REG_FILE._04073_ ),
    .C(\u_cpu.REG_FILE._03006_ ),
    .Y(\u_cpu.REG_FILE._04074_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08797_  (.A_N(\u_cpu.REG_FILE.rf[25][24] ),
    .B(\u_cpu.REG_FILE._03069_ ),
    .X(\u_cpu.REG_FILE._04075_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08798_  (.A1(\u_cpu.REG_FILE.rf[24][24] ),
    .A2(\u_cpu.REG_FILE._03212_ ),
    .B1_N(\u_cpu.REG_FILE._02983_ ),
    .Y(\u_cpu.REG_FILE._04076_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08799_  (.A(\u_cpu.REG_FILE.rf[27][24] ),
    .B_N(\u_cpu.REG_FILE._03077_ ),
    .X(\u_cpu.REG_FILE._04077_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08800_  (.A1(\u_cpu.REG_FILE.rf[26][24] ),
    .A2(\u_cpu.REG_FILE._03125_ ),
    .B1(\u_cpu.REG_FILE._03137_ ),
    .C1(\u_cpu.REG_FILE._04077_ ),
    .Y(\u_cpu.REG_FILE._04078_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08801_  (.A1(\u_cpu.REG_FILE._04075_ ),
    .A2(\u_cpu.REG_FILE._04076_ ),
    .B1(\u_cpu.REG_FILE._02777_ ),
    .C1(\u_cpu.REG_FILE._04078_ ),
    .Y(\u_cpu.REG_FILE._04079_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._08802_  (.A1(\u_cpu.REG_FILE._04074_ ),
    .A2(\u_cpu.REG_FILE._04079_ ),
    .A3(\u_cpu.REG_FILE._03129_ ),
    .B1(\u_cpu.REG_FILE._02996_ ),
    .X(\u_cpu.REG_FILE._04080_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08803_  (.A(\u_cpu.REG_FILE.rf[14][24] ),
    .B(\u_cpu.REG_FILE._02950_ ),
    .Y(\u_cpu.REG_FILE._04081_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08804_  (.A1(\u_cpu.REG_FILE.rf[15][24] ),
    .A2(\u_cpu.REG_FILE._02960_ ),
    .B1(\u_cpu.REG_FILE._02961_ ),
    .Y(\u_cpu.REG_FILE._04082_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08805_  (.A1(\u_cpu.REG_FILE.rf[12][24] ),
    .A2(\u_cpu.REG_FILE._02860_ ),
    .B1_N(\u_cpu.REG_FILE._02817_ ),
    .X(\u_cpu.REG_FILE._04083_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08806_  (.A1(\u_cpu.REG_FILE.rf[13][24] ),
    .A2(\u_cpu.REG_FILE._02956_ ),
    .B1(\u_cpu.REG_FILE._04083_ ),
    .Y(\u_cpu.REG_FILE._04084_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08807_  (.A1(\u_cpu.REG_FILE._04081_ ),
    .A2(\u_cpu.REG_FILE._04082_ ),
    .B1(\u_cpu.REG_FILE._04084_ ),
    .C1(\u_cpu.REG_FILE._02963_ ),
    .Y(\u_cpu.REG_FILE._04085_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08808_  (.A(\u_cpu.REG_FILE.rf[11][24] ),
    .B_N(\u_cpu.REG_FILE._03012_ ),
    .X(\u_cpu.REG_FILE._04086_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08809_  (.A1(\u_cpu.REG_FILE.rf[10][24] ),
    .A2(\u_cpu.REG_FILE._02940_ ),
    .B1(\u_cpu.REG_FILE._02854_ ),
    .C1(\u_cpu.REG_FILE._04086_ ),
    .Y(\u_cpu.REG_FILE._04087_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08810_  (.A1(\u_cpu.REG_FILE.rf[8][24] ),
    .A2(\u_cpu.REG_FILE._03090_ ),
    .B1_N(\u_cpu.REG_FILE._02798_ ),
    .X(\u_cpu.REG_FILE._04088_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08811_  (.A1(\u_cpu.REG_FILE.rf[9][24] ),
    .A2(\u_cpu.REG_FILE._03136_ ),
    .B1(\u_cpu.REG_FILE._04088_ ),
    .Y(\u_cpu.REG_FILE._04089_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08812_  (.A(\u_cpu.REG_FILE._03135_ ),
    .B(\u_cpu.REG_FILE._04087_ ),
    .C(\u_cpu.REG_FILE._04089_ ),
    .Y(\u_cpu.REG_FILE._04090_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08813_  (.A(\u_cpu.REG_FILE._04085_ ),
    .B(\u_cpu.REG_FILE._04090_ ),
    .C(\u_cpu.REG_FILE._03021_ ),
    .Y(\u_cpu.REG_FILE._04091_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._08814_  (.A(\u_cpu.REG_FILE.rf[7][24] ),
    .Y(\u_cpu.REG_FILE._04092_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08815_  (.A1(\u_cpu.REG_FILE.rf[6][24] ),
    .A2(\u_cpu.REG_FILE._02790_ ),
    .B1(\u_cpu.REG_FILE._03198_ ),
    .Y(\u_cpu.REG_FILE._04093_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._08816_  (.A1(\u_cpu.REG_FILE._04092_ ),
    .A2(\u_cpu.REG_FILE._02968_ ),
    .B1(\u_cpu.REG_FILE._04093_ ),
    .Y(\u_cpu.REG_FILE._04094_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08817_  (.A1(\u_cpu.REG_FILE.rf[4][24] ),
    .A2(\u_cpu.REG_FILE._02797_ ),
    .B1_N(\u_cpu.REG_FILE._03201_ ),
    .Y(\u_cpu.REG_FILE._04095_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._08818_  (.A1(\u_cpu.REG_FILE._02378_ ),
    .A2(\u_cpu.REG_FILE._02968_ ),
    .B1(\u_cpu.REG_FILE._04095_ ),
    .Y(\u_cpu.REG_FILE._04096_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08819_  (.A(\u_cpu.REG_FILE.rf[0][24] ),
    .B(\u_cpu.REG_FILE._03204_ ),
    .Y(\u_cpu.REG_FILE._04097_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08820_  (.A_N(\u_cpu.REG_FILE.rf[1][24] ),
    .B(\u_cpu.REG_FILE._03090_ ),
    .X(\u_cpu.REG_FILE._04098_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08821_  (.A(\u_cpu.REG_FILE.rf[3][24] ),
    .B_N(\u_cpu.REG_FILE._02767_ ),
    .X(\u_cpu.REG_FILE._04099_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08822_  (.A1(\u_cpu.REG_FILE.rf[2][24] ),
    .A2(\u_cpu.REG_FILE._03204_ ),
    .B1(\u_cpu.REG_FILE._03133_ ),
    .C1(\u_cpu.REG_FILE._04099_ ),
    .Y(\u_cpu.REG_FILE._04100_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._08823_  (.A1(\u_cpu.REG_FILE._02826_ ),
    .A2(\u_cpu.REG_FILE._04097_ ),
    .A3(\u_cpu.REG_FILE._04098_ ),
    .B1(\u_cpu.REG_FILE._03008_ ),
    .C1(\u_cpu.REG_FILE._04100_ ),
    .Y(\u_cpu.REG_FILE._04101_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._08824_  (.A1(\u_cpu.REG_FILE._03024_ ),
    .A2(\u_cpu.REG_FILE._04094_ ),
    .A3(\u_cpu.REG_FILE._04096_ ),
    .B1(\u_cpu.REG_FILE._02965_ ),
    .C1(\u_cpu.REG_FILE._04101_ ),
    .Y(\u_cpu.REG_FILE._04102_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08825_  (.A(\u_cpu.REG_FILE._02994_ ),
    .B(\u_cpu.REG_FILE._04091_ ),
    .C(\u_cpu.REG_FILE._04102_ ),
    .Y(\u_cpu.REG_FILE._04103_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08826_  (.A1(\u_cpu.REG_FILE._04069_ ),
    .A2(\u_cpu.REG_FILE._04080_ ),
    .B1(\u_cpu.REG_FILE._04103_ ),
    .C1(\u_cpu.REG_FILE._03925_ ),
    .X(\u_cpu.ALU.SrcB[24] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08827_  (.A(\u_cpu.REG_FILE.rf[15][25] ),
    .B_N(\u_cpu.REG_FILE._02754_ ),
    .X(\u_cpu.REG_FILE._04104_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08828_  (.A1(\u_cpu.REG_FILE.rf[14][25] ),
    .A2(\u_cpu.REG_FILE._03418_ ),
    .B1(\u_cpu.REG_FILE._02752_ ),
    .C1(\u_cpu.REG_FILE._04104_ ),
    .Y(\u_cpu.REG_FILE._04105_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08829_  (.A1(\u_cpu.REG_FILE.rf[12][25] ),
    .A2(\u_cpu.REG_FILE._02974_ ),
    .B1_N(\u_cpu.REG_FILE._02761_ ),
    .X(\u_cpu.REG_FILE._04106_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08830_  (.A1(\u_cpu.REG_FILE.rf[13][25] ),
    .A2(\u_cpu.REG_FILE._02759_ ),
    .B1(\u_cpu.REG_FILE._04106_ ),
    .Y(\u_cpu.REG_FILE._04107_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08831_  (.A(\u_cpu.REG_FILE._04105_ ),
    .B(\u_cpu.REG_FILE._04107_ ),
    .C(\u_cpu.REG_FILE._02978_ ),
    .Y(\u_cpu.REG_FILE._04108_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08832_  (.A_N(\u_cpu.REG_FILE.rf[9][25] ),
    .B(\u_cpu.REG_FILE._02945_ ),
    .X(\u_cpu.REG_FILE._04109_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08833_  (.A1(\u_cpu.REG_FILE.rf[8][25] ),
    .A2(\u_cpu.REG_FILE._02816_ ),
    .B1_N(\u_cpu.REG_FILE._02947_ ),
    .Y(\u_cpu.REG_FILE._04110_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08834_  (.A(\u_cpu.REG_FILE.rf[11][25] ),
    .B_N(\u_cpu.REG_FILE._02986_ ),
    .X(\u_cpu.REG_FILE._04111_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08835_  (.A1(\u_cpu.REG_FILE.rf[10][25] ),
    .A2(\u_cpu.REG_FILE._02824_ ),
    .B1(\u_cpu.REG_FILE._02846_ ),
    .C1(\u_cpu.REG_FILE._04111_ ),
    .Y(\u_cpu.REG_FILE._04112_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08836_  (.A1(\u_cpu.REG_FILE._04109_ ),
    .A2(\u_cpu.REG_FILE._04110_ ),
    .B1(\u_cpu.REG_FILE._03062_ ),
    .C1(\u_cpu.REG_FILE._04112_ ),
    .Y(\u_cpu.REG_FILE._04113_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08837_  (.A(\u_cpu.REG_FILE._04108_ ),
    .B(\u_cpu.REG_FILE._04113_ ),
    .C(\u_cpu.REG_FILE._03218_ ),
    .Y(\u_cpu.REG_FILE._04114_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08838_  (.A1(\u_cpu.REG_FILE.rf[4][25] ),
    .A2(\u_cpu.REG_FILE._02793_ ),
    .B1_N(\u_cpu.REG_FILE._02954_ ),
    .Y(\u_cpu.REG_FILE._04115_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._08839_  (.A1(\u_cpu.REG_FILE._02426_ ),
    .A2(\u_cpu.REG_FILE._02946_ ),
    .B1(\u_cpu.REG_FILE._04115_ ),
    .Y(\u_cpu.REG_FILE._04116_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08840_  (.A1(\u_cpu.REG_FILE.rf[6][25] ),
    .A2(\u_cpu.REG_FILE._03331_ ),
    .B1(\u_cpu.REG_FILE._03407_ ),
    .Y(\u_cpu.REG_FILE._04117_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08841_  (.A_N(\u_cpu.REG_FILE.rf[7][25] ),
    .B(\u_cpu.REG_FILE._02808_ ),
    .X(\u_cpu.REG_FILE._04118_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08842_  (.A1(\u_cpu.REG_FILE._04117_ ),
    .A2(\u_cpu.REG_FILE._04118_ ),
    .B1(\u_cpu.REG_FILE._03434_ ),
    .Y(\u_cpu.REG_FILE._04119_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08843_  (.A_N(\u_cpu.REG_FILE.rf[1][25] ),
    .B(\u_cpu.REG_FILE._03530_ ),
    .X(\u_cpu.REG_FILE._04120_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08844_  (.A1(\u_cpu.REG_FILE.rf[0][25] ),
    .A2(\u_cpu.REG_FILE._03287_ ),
    .B1_N(\u_cpu.REG_FILE._02794_ ),
    .Y(\u_cpu.REG_FILE._04121_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08845_  (.A(\u_cpu.REG_FILE.rf[3][25] ),
    .B_N(\u_cpu.REG_FILE._03337_ ),
    .X(\u_cpu.REG_FILE._04122_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08846_  (.A1(\u_cpu.REG_FILE.rf[2][25] ),
    .A2(\u_cpu.REG_FILE._02903_ ),
    .B1(\u_cpu.REG_FILE._03026_ ),
    .C1(\u_cpu.REG_FILE._04122_ ),
    .Y(\u_cpu.REG_FILE._04123_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08847_  (.A1(\u_cpu.REG_FILE._04120_ ),
    .A2(\u_cpu.REG_FILE._04121_ ),
    .B1(\u_cpu.REG_FILE._02858_ ),
    .C1(\u_cpu.REG_FILE._04123_ ),
    .Y(\u_cpu.REG_FILE._04124_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08848_  (.A1(\u_cpu.REG_FILE._04116_ ),
    .A2(\u_cpu.REG_FILE._04119_ ),
    .B1(\u_cpu.REG_FILE._02965_ ),
    .C1(\u_cpu.REG_FILE._04124_ ),
    .Y(\u_cpu.REG_FILE._04125_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._08849_  (.A(\u_cpu.REG_FILE._04114_ ),
    .B(\u_cpu.REG_FILE._04125_ ),
    .Y(\u_cpu.REG_FILE._04126_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08850_  (.A(\u_cpu.REG_FILE.rf[27][25] ),
    .B_N(\u_cpu.REG_FILE._02871_ ),
    .X(\u_cpu.REG_FILE._04127_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08851_  (.A1(\u_cpu.REG_FILE.rf[26][25] ),
    .A2(\u_cpu.REG_FILE._02982_ ),
    .B1(\u_cpu.REG_FILE._03000_ ),
    .C1(\u_cpu.REG_FILE._04127_ ),
    .X(\u_cpu.REG_FILE._04128_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08852_  (.A1(\u_cpu.REG_FILE.rf[24][25] ),
    .A2(\u_cpu.REG_FILE._03445_ ),
    .B1_N(\u_cpu.REG_FILE._02865_ ),
    .X(\u_cpu.REG_FILE._04129_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08853_  (.A(\u_cpu.REG_FILE.rf[25][25] ),
    .B_N(\u_cpu.REG_FILE._02832_ ),
    .X(\u_cpu.REG_FILE._04130_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._08854_  (.A1(\u_cpu.REG_FILE._04129_ ),
    .A2(\u_cpu.REG_FILE._04130_ ),
    .B1(\u_cpu.REG_FILE._02764_ ),
    .X(\u_cpu.REG_FILE._04131_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08855_  (.A(\u_cpu.REG_FILE.rf[30][25] ),
    .B(\u_cpu.REG_FILE._03063_ ),
    .Y(\u_cpu.REG_FILE._04132_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08856_  (.A1(\u_cpu.REG_FILE.rf[31][25] ),
    .A2(\u_cpu.REG_FILE._03297_ ),
    .B1(\u_cpu.REG_FILE._02854_ ),
    .Y(\u_cpu.REG_FILE._04133_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08857_  (.A(\u_cpu.REG_FILE.rf[28][25] ),
    .B(\u_cpu.REG_FILE._02916_ ),
    .Y(\u_cpu.REG_FILE._04134_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08858_  (.A1(\u_cpu.REG_FILE.rf[29][25] ),
    .A2(\u_cpu.REG_FILE._03351_ ),
    .B1_N(\u_cpu.REG_FILE._02947_ ),
    .Y(\u_cpu.REG_FILE._04135_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._08859_  (.A1(\u_cpu.REG_FILE._04132_ ),
    .A2(\u_cpu.REG_FILE._04133_ ),
    .B1(\u_cpu.REG_FILE._04134_ ),
    .B2(\u_cpu.REG_FILE._04135_ ),
    .C1(\u_cpu.REG_FILE._02919_ ),
    .Y(\u_cpu.REG_FILE._04136_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08860_  (.A1(\u_cpu.REG_FILE._04128_ ),
    .A2(\u_cpu.REG_FILE._04131_ ),
    .B1(\u_cpu.REG_FILE._02836_ ),
    .C1(\u_cpu.REG_FILE._04136_ ),
    .Y(\u_cpu.REG_FILE._04137_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08861_  (.A1(\u_cpu.REG_FILE.rf[18][25] ),
    .A2(\u_cpu.REG_FILE._02923_ ),
    .B1(\u_cpu.REG_FILE._03249_ ),
    .Y(\u_cpu.REG_FILE._04138_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08862_  (.A(\u_cpu.REG_FILE.rf[19][25] ),
    .B(\u_cpu.REG_FILE._03037_ ),
    .Y(\u_cpu.REG_FILE._04139_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08863_  (.A1(\u_cpu.REG_FILE.rf[16][25] ),
    .A2(\u_cpu.REG_FILE._03038_ ),
    .B1_N(\u_cpu.REG_FILE._03039_ ),
    .X(\u_cpu.REG_FILE._04140_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08864_  (.A1(\u_cpu.REG_FILE.rf[17][25] ),
    .A2(\u_cpu.REG_FILE._03304_ ),
    .B1(\u_cpu.REG_FILE._04140_ ),
    .Y(\u_cpu.REG_FILE._04141_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08865_  (.A1(\u_cpu.REG_FILE._04138_ ),
    .A2(\u_cpu.REG_FILE._04139_ ),
    .B1(\u_cpu.REG_FILE._03292_ ),
    .C1(\u_cpu.REG_FILE._04141_ ),
    .Y(\u_cpu.REG_FILE._04142_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._08866_  (.A(\u_cpu.REG_FILE.rf[22][25] ),
    .B(\u_cpu.REG_FILE._02810_ ),
    .X(\u_cpu.REG_FILE._04143_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08867_  (.A1(\u_cpu.REG_FILE.rf[23][25] ),
    .A2(\u_cpu.REG_FILE._03132_ ),
    .B1(\u_cpu.REG_FILE._03255_ ),
    .C1(\u_cpu.REG_FILE._04143_ ),
    .Y(\u_cpu.REG_FILE._04144_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08868_  (.A1(\u_cpu.REG_FILE.rf[20][25] ),
    .A2(\u_cpu.REG_FILE._03016_ ),
    .B1_N(\u_cpu.REG_FILE._03017_ ),
    .X(\u_cpu.REG_FILE._04145_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08869_  (.A1(\u_cpu.REG_FILE.rf[21][25] ),
    .A2(\u_cpu.REG_FILE._03015_ ),
    .B1(\u_cpu.REG_FILE._04145_ ),
    .Y(\u_cpu.REG_FILE._04146_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08870_  (.A(\u_cpu.REG_FILE._04144_ ),
    .B(\u_cpu.REG_FILE._04146_ ),
    .C(\u_cpu.REG_FILE._03074_ ),
    .Y(\u_cpu.REG_FILE._04147_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08871_  (.A(\u_cpu.REG_FILE._02922_ ),
    .B(\u_cpu.REG_FILE._04142_ ),
    .C(\u_cpu.REG_FILE._04147_ ),
    .Y(\u_cpu.REG_FILE._04148_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08872_  (.A(\u_cpu.REG_FILE._04137_ ),
    .B(\u_cpu.REG_FILE._04148_ ),
    .C(\u_cpu.REG_FILE._02745_ ),
    .Y(\u_cpu.REG_FILE._04149_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08873_  (.A1(\u_cpu.REG_FILE._02746_ ),
    .A2(\u_cpu.REG_FILE._04126_ ),
    .B1(\u_cpu.REG_FILE._04149_ ),
    .C1(\u_cpu.REG_FILE._03925_ ),
    .X(\u_cpu.ALU.SrcB[25] ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08874_  (.A1(\u_cpu.REG_FILE.rf[18][26] ),
    .A2(\u_cpu.REG_FILE._03653_ ),
    .B1(\u_cpu.REG_FILE._03298_ ),
    .Y(\u_cpu.REG_FILE._04150_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._08875_  (.A1(\u_cpu.REG_FILE._02486_ ),
    .A2(\u_cpu.REG_FILE._02791_ ),
    .B1(\u_cpu.REG_FILE._04150_ ),
    .Y(\u_cpu.REG_FILE._04151_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08876_  (.A(\u_cpu.REG_FILE.rf[16][26] ),
    .B(\u_cpu.REG_FILE._03371_ ),
    .Y(\u_cpu.REG_FILE._04152_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._08877_  (.A1(\u_cpu.REG_FILE._02489_ ),
    .A2(\u_cpu.REG_FILE._03166_ ),
    .B1(\u_cpu.REG_FILE._03057_ ),
    .C1(\u_cpu.REG_FILE._04152_ ),
    .Y(\u_cpu.REG_FILE._04153_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08878_  (.A1(\u_cpu.REG_FILE.rf[20][26] ),
    .A2(\u_cpu.REG_FILE._02853_ ),
    .B1_N(\u_cpu.REG_FILE._03050_ ),
    .Y(\u_cpu.REG_FILE._04154_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08879_  (.A(\u_cpu.REG_FILE.rf[21][26] ),
    .B(\u_cpu.REG_FILE._02859_ ),
    .Y(\u_cpu.REG_FILE._04155_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08880_  (.A(\u_cpu.REG_FILE.rf[22][26] ),
    .B(\u_cpu.REG_FILE._02958_ ),
    .Y(\u_cpu.REG_FILE._04156_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08881_  (.A1(\u_cpu.REG_FILE.rf[23][26] ),
    .A2(\u_cpu.REG_FILE._03114_ ),
    .B1(\u_cpu.REG_FILE._03377_ ),
    .Y(\u_cpu.REG_FILE._04157_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._08882_  (.A1(\u_cpu.REG_FILE._04154_ ),
    .A2(\u_cpu.REG_FILE._04155_ ),
    .B1(\u_cpu.REG_FILE._04156_ ),
    .B2(\u_cpu.REG_FILE._04157_ ),
    .C1(\u_cpu.REG_FILE._02848_ ),
    .Y(\u_cpu.REG_FILE._04158_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.REG_FILE._08883_  (.A1(\u_cpu.REG_FILE._02765_ ),
    .A2(\u_cpu.REG_FILE._04151_ ),
    .A3(\u_cpu.REG_FILE._04153_ ),
    .B1(\u_cpu.REG_FILE._04158_ ),
    .C1(\u_cpu.REG_FILE._03023_ ),
    .X(\u_cpu.REG_FILE._04159_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08884_  (.A(\u_cpu.REG_FILE.rf[28][26] ),
    .B(\u_cpu.REG_FILE._03058_ ),
    .Y(\u_cpu.REG_FILE._04160_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08885_  (.A_N(\u_cpu.REG_FILE.rf[29][26] ),
    .B(\u_cpu.REG_FILE._03060_ ),
    .X(\u_cpu.REG_FILE._04161_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08886_  (.A(\u_cpu.REG_FILE.rf[31][26] ),
    .B_N(\u_cpu.REG_FILE._03065_ ),
    .X(\u_cpu.REG_FILE._04162_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08887_  (.A1(\u_cpu.REG_FILE.rf[30][26] ),
    .A2(\u_cpu.REG_FILE._02772_ ),
    .B1(\u_cpu.REG_FILE._03064_ ),
    .C1(\u_cpu.REG_FILE._04162_ ),
    .Y(\u_cpu.REG_FILE._04163_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._08888_  (.A1(\u_cpu.REG_FILE._03709_ ),
    .A2(\u_cpu.REG_FILE._04160_ ),
    .A3(\u_cpu.REG_FILE._04161_ ),
    .B1(\u_cpu.REG_FILE._03221_ ),
    .C1(\u_cpu.REG_FILE._04163_ ),
    .Y(\u_cpu.REG_FILE._04164_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08889_  (.A_N(\u_cpu.REG_FILE.rf[25][26] ),
    .B(\u_cpu.REG_FILE._03069_ ),
    .X(\u_cpu.REG_FILE._04165_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08890_  (.A1(\u_cpu.REG_FILE.rf[24][26] ),
    .A2(\u_cpu.REG_FILE._03212_ ),
    .B1_N(\u_cpu.REG_FILE._03072_ ),
    .Y(\u_cpu.REG_FILE._04166_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08891_  (.A(\u_cpu.REG_FILE.rf[27][26] ),
    .B_N(\u_cpu.REG_FILE._03077_ ),
    .X(\u_cpu.REG_FILE._04167_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08892_  (.A1(\u_cpu.REG_FILE.rf[26][26] ),
    .A2(\u_cpu.REG_FILE._03125_ ),
    .B1(\u_cpu.REG_FILE._03137_ ),
    .C1(\u_cpu.REG_FILE._04167_ ),
    .Y(\u_cpu.REG_FILE._04168_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08893_  (.A1(\u_cpu.REG_FILE._04165_ ),
    .A2(\u_cpu.REG_FILE._04166_ ),
    .B1(\u_cpu.REG_FILE._02777_ ),
    .C1(\u_cpu.REG_FILE._04168_ ),
    .Y(\u_cpu.REG_FILE._04169_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._08894_  (.A1(\u_cpu.REG_FILE._04164_ ),
    .A2(\u_cpu.REG_FILE._04169_ ),
    .A3(\u_cpu.REG_FILE._03129_ ),
    .B1(\u_cpu.REG_FILE._02996_ ),
    .X(\u_cpu.REG_FILE._04170_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08895_  (.A_N(\u_cpu.REG_FILE.rf[1][26] ),
    .B(\u_cpu.REG_FILE._02748_ ),
    .X(\u_cpu.REG_FILE._04171_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08896_  (.A(\u_cpu.REG_FILE.rf[0][26] ),
    .B(\u_cpu.REG_FILE._03075_ ),
    .Y(\u_cpu.REG_FILE._04172_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08897_  (.A(\u_cpu.REG_FILE.rf[3][26] ),
    .B_N(\u_cpu.REG_FILE._02949_ ),
    .X(\u_cpu.REG_FILE._04173_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08898_  (.A1(\u_cpu.REG_FILE.rf[2][26] ),
    .A2(\u_cpu.REG_FILE._02987_ ),
    .B1(\u_cpu.REG_FILE._02988_ ),
    .C1(\u_cpu.REG_FILE._04173_ ),
    .Y(\u_cpu.REG_FILE._04174_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.REG_FILE._08899_  (.A1(\u_cpu.REG_FILE._03709_ ),
    .A2(\u_cpu.REG_FILE._04171_ ),
    .A3(\u_cpu.REG_FILE._04172_ ),
    .B1(\u_cpu.REG_FILE._03800_ ),
    .C1(\u_cpu.REG_FILE._04174_ ),
    .X(\u_cpu.REG_FILE._04175_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08900_  (.A(\u_cpu.REG_FILE.rf[4][26] ),
    .B(\u_cpu.REG_FILE._03815_ ),
    .Y(\u_cpu.REG_FILE._04176_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._08901_  (.A1(\u_cpu.REG_FILE._02473_ ),
    .A2(\u_cpu.REG_FILE._03418_ ),
    .B1(\u_cpu.REG_FILE._03308_ ),
    .C1(\u_cpu.REG_FILE._04176_ ),
    .Y(\u_cpu.REG_FILE._04177_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08902_  (.A1(\u_cpu.REG_FILE.rf[6][26] ),
    .A2(\u_cpu.REG_FILE._03204_ ),
    .B1(\u_cpu.REG_FILE._03198_ ),
    .Y(\u_cpu.REG_FILE._04178_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08903_  (.A_N(\u_cpu.REG_FILE.rf[7][26] ),
    .B(\u_cpu.REG_FILE._02880_ ),
    .X(\u_cpu.REG_FILE._04179_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08904_  (.A1(\u_cpu.REG_FILE._04178_ ),
    .A2(\u_cpu.REG_FILE._04179_ ),
    .B1(\u_cpu.REG_FILE._03434_ ),
    .Y(\u_cpu.REG_FILE._04180_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08905_  (.A1(\u_cpu.REG_FILE._04177_ ),
    .A2(\u_cpu.REG_FILE._04180_ ),
    .B1_N(\u_cpu.REG_FILE._03141_ ),
    .Y(\u_cpu.REG_FILE._04181_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08906_  (.A_N(\u_cpu.REG_FILE.rf[13][26] ),
    .B(\u_cpu.REG_FILE._02760_ ),
    .X(\u_cpu.REG_FILE._04182_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08907_  (.A1(\u_cpu.REG_FILE.rf[12][26] ),
    .A2(\u_cpu.REG_FILE._02953_ ),
    .B1_N(\u_cpu.REG_FILE._02954_ ),
    .Y(\u_cpu.REG_FILE._04183_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08908_  (.A(\u_cpu.REG_FILE.rf[15][26] ),
    .B_N(\u_cpu.REG_FILE._02810_ ),
    .X(\u_cpu.REG_FILE._04184_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08909_  (.A1(\u_cpu.REG_FILE.rf[14][26] ),
    .A2(\u_cpu.REG_FILE._03287_ ),
    .B1(\u_cpu.REG_FILE._03470_ ),
    .C1(\u_cpu.REG_FILE._04184_ ),
    .Y(\u_cpu.REG_FILE._04185_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08910_  (.A1(\u_cpu.REG_FILE._04182_ ),
    .A2(\u_cpu.REG_FILE._04183_ ),
    .B1(\u_cpu.REG_FILE._04185_ ),
    .Y(\u_cpu.REG_FILE._04186_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08911_  (.A(\u_cpu.REG_FILE.rf[8][26] ),
    .B(\u_cpu.REG_FILE._03025_ ),
    .Y(\u_cpu.REG_FILE._04187_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08912_  (.A1(\u_cpu.REG_FILE.rf[9][26] ),
    .A2(\u_cpu.REG_FILE._03297_ ),
    .B1_N(\u_cpu.REG_FILE._02838_ ),
    .Y(\u_cpu.REG_FILE._04188_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._08913_  (.A(\u_cpu.REG_FILE.rf[10][26] ),
    .B(\u_cpu.REG_FILE._02767_ ),
    .X(\u_cpu.REG_FILE._04189_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08914_  (.A1(\u_cpu.REG_FILE.rf[11][26] ),
    .A2(\u_cpu.REG_FILE._03297_ ),
    .B1(\u_cpu.REG_FILE._02799_ ),
    .C1(\u_cpu.REG_FILE._04189_ ),
    .Y(\u_cpu.REG_FILE._04190_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08915_  (.A1(\u_cpu.REG_FILE._04187_ ),
    .A2(\u_cpu.REG_FILE._04188_ ),
    .B1(\u_cpu.REG_FILE._03008_ ),
    .C1(\u_cpu.REG_FILE._04190_ ),
    .Y(\u_cpu.REG_FILE._04191_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08916_  (.A1(\u_cpu.REG_FILE._03024_ ),
    .A2(\u_cpu.REG_FILE._04186_ ),
    .B1(\u_cpu.REG_FILE._04191_ ),
    .C1(\u_cpu.REG_FILE._03218_ ),
    .Y(\u_cpu.REG_FILE._04192_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08917_  (.A1(\u_cpu.REG_FILE._04175_ ),
    .A2(\u_cpu.REG_FILE._04181_ ),
    .B1(\u_cpu.REG_FILE._02994_ ),
    .C1(\u_cpu.REG_FILE._04192_ ),
    .Y(\u_cpu.REG_FILE._04193_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08918_  (.A1(\u_cpu.REG_FILE._04159_ ),
    .A2(\u_cpu.REG_FILE._04170_ ),
    .B1(\u_cpu.REG_FILE._04193_ ),
    .C1(\u_cpu.REG_FILE._03925_ ),
    .X(\u_cpu.ALU.SrcB[26] ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._08919_  (.A(\u_cpu.REG_FILE.rf[19][27] ),
    .Y(\u_cpu.REG_FILE._04194_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08920_  (.A1(\u_cpu.REG_FILE.rf[18][27] ),
    .A2(\u_cpu.REG_FILE._03653_ ),
    .B1(\u_cpu.REG_FILE._03298_ ),
    .Y(\u_cpu.REG_FILE._04195_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._08921_  (.A1(\u_cpu.REG_FILE._04194_ ),
    .A2(\u_cpu.REG_FILE._02791_ ),
    .B1(\u_cpu.REG_FILE._04195_ ),
    .Y(\u_cpu.REG_FILE._04196_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu.REG_FILE._08922_  (.A(\u_cpu.REG_FILE.rf[17][27] ),
    .Y(\u_cpu.REG_FILE._04197_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08923_  (.A(\u_cpu.REG_FILE.rf[16][27] ),
    .B(\u_cpu.REG_FILE._03371_ ),
    .Y(\u_cpu.REG_FILE._04198_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._08924_  (.A1(\u_cpu.REG_FILE._04197_ ),
    .A2(\u_cpu.REG_FILE._03166_ ),
    .B1(\u_cpu.REG_FILE._03057_ ),
    .C1(\u_cpu.REG_FILE._04198_ ),
    .Y(\u_cpu.REG_FILE._04199_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08925_  (.A1(\u_cpu.REG_FILE.rf[20][27] ),
    .A2(\u_cpu.REG_FILE._02853_ ),
    .B1_N(\u_cpu.REG_FILE._03050_ ),
    .Y(\u_cpu.REG_FILE._04200_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08926_  (.A(\u_cpu.REG_FILE.rf[21][27] ),
    .B(\u_cpu.REG_FILE._02859_ ),
    .Y(\u_cpu.REG_FILE._04201_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08927_  (.A(\u_cpu.REG_FILE.rf[22][27] ),
    .B(\u_cpu.REG_FILE._02987_ ),
    .Y(\u_cpu.REG_FILE._04202_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08928_  (.A1(\u_cpu.REG_FILE.rf[23][27] ),
    .A2(\u_cpu.REG_FILE._03114_ ),
    .B1(\u_cpu.REG_FILE._03377_ ),
    .Y(\u_cpu.REG_FILE._04203_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._08929_  (.A1(\u_cpu.REG_FILE._04200_ ),
    .A2(\u_cpu.REG_FILE._04201_ ),
    .B1(\u_cpu.REG_FILE._04202_ ),
    .B2(\u_cpu.REG_FILE._04203_ ),
    .C1(\u_cpu.REG_FILE._02848_ ),
    .Y(\u_cpu.REG_FILE._04204_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.REG_FILE._08930_  (.A1(\u_cpu.REG_FILE._02765_ ),
    .A2(\u_cpu.REG_FILE._04196_ ),
    .A3(\u_cpu.REG_FILE._04199_ ),
    .B1(\u_cpu.REG_FILE._04204_ ),
    .C1(\u_cpu.REG_FILE._03023_ ),
    .X(\u_cpu.REG_FILE._04205_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08931_  (.A(\u_cpu.REG_FILE.rf[31][27] ),
    .B_N(\u_cpu.REG_FILE._02970_ ),
    .X(\u_cpu.REG_FILE._04206_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08932_  (.A1(\u_cpu.REG_FILE.rf[30][27] ),
    .A2(\u_cpu.REG_FILE._02749_ ),
    .B1(\u_cpu.REG_FILE._02969_ ),
    .C1(\u_cpu.REG_FILE._04206_ ),
    .Y(\u_cpu.REG_FILE._04207_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08933_  (.A1(\u_cpu.REG_FILE.rf[28][27] ),
    .A2(\u_cpu.REG_FILE._02830_ ),
    .B1_N(\u_cpu.REG_FILE._02975_ ),
    .X(\u_cpu.REG_FILE._04208_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08934_  (.A1(\u_cpu.REG_FILE.rf[29][27] ),
    .A2(\u_cpu.REG_FILE._02973_ ),
    .B1(\u_cpu.REG_FILE._04208_ ),
    .Y(\u_cpu.REG_FILE._04209_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08935_  (.A(\u_cpu.REG_FILE._04207_ ),
    .B(\u_cpu.REG_FILE._04209_ ),
    .C(\u_cpu.REG_FILE._03006_ ),
    .Y(\u_cpu.REG_FILE._04210_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08936_  (.A_N(\u_cpu.REG_FILE.rf[25][27] ),
    .B(\u_cpu.REG_FILE._03069_ ),
    .X(\u_cpu.REG_FILE._04211_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08937_  (.A1(\u_cpu.REG_FILE.rf[24][27] ),
    .A2(\u_cpu.REG_FILE._03212_ ),
    .B1_N(\u_cpu.REG_FILE._03072_ ),
    .Y(\u_cpu.REG_FILE._04212_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08938_  (.A(\u_cpu.REG_FILE.rf[27][27] ),
    .B_N(\u_cpu.REG_FILE._03077_ ),
    .X(\u_cpu.REG_FILE._04213_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08939_  (.A1(\u_cpu.REG_FILE.rf[26][27] ),
    .A2(\u_cpu.REG_FILE._03125_ ),
    .B1(\u_cpu.REG_FILE._03137_ ),
    .C1(\u_cpu.REG_FILE._04213_ ),
    .Y(\u_cpu.REG_FILE._04214_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08940_  (.A1(\u_cpu.REG_FILE._04211_ ),
    .A2(\u_cpu.REG_FILE._04212_ ),
    .B1(\u_cpu.REG_FILE._02777_ ),
    .C1(\u_cpu.REG_FILE._04214_ ),
    .Y(\u_cpu.REG_FILE._04215_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._08941_  (.A1(\u_cpu.REG_FILE._04210_ ),
    .A2(\u_cpu.REG_FILE._04215_ ),
    .A3(\u_cpu.REG_FILE._03129_ ),
    .B1(\u_cpu.REG_FILE._02996_ ),
    .X(\u_cpu.REG_FILE._04216_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08942_  (.A(\u_cpu.REG_FILE.rf[0][27] ),
    .B(\u_cpu.REG_FILE._02816_ ),
    .Y(\u_cpu.REG_FILE._04217_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08943_  (.A_N(\u_cpu.REG_FILE.rf[1][27] ),
    .B(\u_cpu.REG_FILE._03530_ ),
    .X(\u_cpu.REG_FILE._04218_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08944_  (.A(\u_cpu.REG_FILE.rf[3][27] ),
    .B_N(\u_cpu.REG_FILE._02949_ ),
    .X(\u_cpu.REG_FILE._04219_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08945_  (.A1(\u_cpu.REG_FILE.rf[2][27] ),
    .A2(\u_cpu.REG_FILE._02987_ ),
    .B1(\u_cpu.REG_FILE._02988_ ),
    .C1(\u_cpu.REG_FILE._04219_ ),
    .Y(\u_cpu.REG_FILE._04220_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.REG_FILE._08946_  (.A1(\u_cpu.REG_FILE._03403_ ),
    .A2(\u_cpu.REG_FILE._04217_ ),
    .A3(\u_cpu.REG_FILE._04218_ ),
    .B1(\u_cpu.REG_FILE._03800_ ),
    .C1(\u_cpu.REG_FILE._04220_ ),
    .X(\u_cpu.REG_FILE._04221_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08947_  (.A(\u_cpu.REG_FILE.rf[4][27] ),
    .B(\u_cpu.REG_FILE._03815_ ),
    .Y(\u_cpu.REG_FILE._04222_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._08948_  (.A1(\u_cpu.REG_FILE._02521_ ),
    .A2(\u_cpu.REG_FILE._03418_ ),
    .B1(\u_cpu.REG_FILE._03308_ ),
    .C1(\u_cpu.REG_FILE._04222_ ),
    .Y(\u_cpu.REG_FILE._04223_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08949_  (.A1(\u_cpu.REG_FILE.rf[6][27] ),
    .A2(\u_cpu.REG_FILE._03204_ ),
    .B1(\u_cpu.REG_FILE._03198_ ),
    .Y(\u_cpu.REG_FILE._04224_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08950_  (.A_N(\u_cpu.REG_FILE.rf[7][27] ),
    .B(\u_cpu.REG_FILE._02880_ ),
    .X(\u_cpu.REG_FILE._04225_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08951_  (.A1(\u_cpu.REG_FILE._04224_ ),
    .A2(\u_cpu.REG_FILE._04225_ ),
    .B1(\u_cpu.REG_FILE._03434_ ),
    .Y(\u_cpu.REG_FILE._04226_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08952_  (.A1(\u_cpu.REG_FILE._04223_ ),
    .A2(\u_cpu.REG_FILE._04226_ ),
    .B1_N(\u_cpu.REG_FILE._03141_ ),
    .Y(\u_cpu.REG_FILE._04227_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08953_  (.A_N(\u_cpu.REG_FILE.rf[13][27] ),
    .B(\u_cpu.REG_FILE._02760_ ),
    .X(\u_cpu.REG_FILE._04228_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08954_  (.A1(\u_cpu.REG_FILE.rf[12][27] ),
    .A2(\u_cpu.REG_FILE._02953_ ),
    .B1_N(\u_cpu.REG_FILE._02954_ ),
    .Y(\u_cpu.REG_FILE._04229_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08955_  (.A(\u_cpu.REG_FILE.rf[15][27] ),
    .B_N(\u_cpu.REG_FILE._02810_ ),
    .X(\u_cpu.REG_FILE._04230_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08956_  (.A1(\u_cpu.REG_FILE.rf[14][27] ),
    .A2(\u_cpu.REG_FILE._03287_ ),
    .B1(\u_cpu.REG_FILE._03470_ ),
    .C1(\u_cpu.REG_FILE._04230_ ),
    .Y(\u_cpu.REG_FILE._04231_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08957_  (.A1(\u_cpu.REG_FILE._04228_ ),
    .A2(\u_cpu.REG_FILE._04229_ ),
    .B1(\u_cpu.REG_FILE._04231_ ),
    .Y(\u_cpu.REG_FILE._04232_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08958_  (.A(\u_cpu.REG_FILE.rf[10][27] ),
    .B(\u_cpu.REG_FILE._03025_ ),
    .Y(\u_cpu.REG_FILE._04233_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08959_  (.A1(\u_cpu.REG_FILE.rf[11][27] ),
    .A2(\u_cpu.REG_FILE._02758_ ),
    .B1(\u_cpu.REG_FILE._03470_ ),
    .Y(\u_cpu.REG_FILE._04234_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08960_  (.A1(\u_cpu.REG_FILE.rf[8][27] ),
    .A2(\u_cpu.REG_FILE._03337_ ),
    .B1_N(\u_cpu.REG_FILE._02773_ ),
    .X(\u_cpu.REG_FILE._04235_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08961_  (.A1(\u_cpu.REG_FILE.rf[9][27] ),
    .A2(\u_cpu.REG_FILE._03297_ ),
    .B1(\u_cpu.REG_FILE._04235_ ),
    .Y(\u_cpu.REG_FILE._04236_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08962_  (.A1(\u_cpu.REG_FILE._04233_ ),
    .A2(\u_cpu.REG_FILE._04234_ ),
    .B1(\u_cpu.REG_FILE._04236_ ),
    .C1(\u_cpu.REG_FILE._02814_ ),
    .Y(\u_cpu.REG_FILE._04237_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08963_  (.A1(\u_cpu.REG_FILE._03024_ ),
    .A2(\u_cpu.REG_FILE._04232_ ),
    .B1(\u_cpu.REG_FILE._04237_ ),
    .C1(\u_cpu.REG_FILE._02836_ ),
    .Y(\u_cpu.REG_FILE._04238_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08964_  (.A1(\u_cpu.REG_FILE._04221_ ),
    .A2(\u_cpu.REG_FILE._04227_ ),
    .B1(\u_cpu.REG_FILE._02994_ ),
    .C1(\u_cpu.REG_FILE._04238_ ),
    .Y(\u_cpu.REG_FILE._04239_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._08965_  (.A1(\u_cpu.REG_FILE._04205_ ),
    .A2(\u_cpu.REG_FILE._04216_ ),
    .B1(\u_cpu.REG_FILE._04239_ ),
    .C1(\u_cpu.REG_FILE._03925_ ),
    .X(\u_cpu.ALU.SrcB[27] ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08966_  (.A1(\u_cpu.REG_FILE.rf[18][28] ),
    .A2(\u_cpu.REG_FILE._03653_ ),
    .B1(\u_cpu.REG_FILE._03298_ ),
    .Y(\u_cpu.REG_FILE._04240_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._08967_  (.A1(\u_cpu.REG_FILE._02592_ ),
    .A2(\u_cpu.REG_FILE._02791_ ),
    .B1(\u_cpu.REG_FILE._04240_ ),
    .Y(\u_cpu.REG_FILE._04241_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08968_  (.A(\u_cpu.REG_FILE.rf[16][28] ),
    .B(\u_cpu.REG_FILE._03371_ ),
    .Y(\u_cpu.REG_FILE._04242_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._08969_  (.A1(\u_cpu.REG_FILE._02595_ ),
    .A2(\u_cpu.REG_FILE._03166_ ),
    .B1(\u_cpu.REG_FILE._03057_ ),
    .C1(\u_cpu.REG_FILE._04242_ ),
    .Y(\u_cpu.REG_FILE._04243_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08970_  (.A1(\u_cpu.REG_FILE.rf[20][28] ),
    .A2(\u_cpu.REG_FILE._02853_ ),
    .B1_N(\u_cpu.REG_FILE._02838_ ),
    .Y(\u_cpu.REG_FILE._04244_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08971_  (.A(\u_cpu.REG_FILE.rf[21][28] ),
    .B(\u_cpu.REG_FILE._02859_ ),
    .Y(\u_cpu.REG_FILE._04245_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08972_  (.A(\u_cpu.REG_FILE.rf[22][28] ),
    .B(\u_cpu.REG_FILE._02987_ ),
    .Y(\u_cpu.REG_FILE._04246_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08973_  (.A1(\u_cpu.REG_FILE.rf[23][28] ),
    .A2(\u_cpu.REG_FILE._03114_ ),
    .B1(\u_cpu.REG_FILE._03377_ ),
    .Y(\u_cpu.REG_FILE._04247_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._08974_  (.A1(\u_cpu.REG_FILE._04244_ ),
    .A2(\u_cpu.REG_FILE._04245_ ),
    .B1(\u_cpu.REG_FILE._04246_ ),
    .B2(\u_cpu.REG_FILE._04247_ ),
    .C1(\u_cpu.REG_FILE._02848_ ),
    .Y(\u_cpu.REG_FILE._04248_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.REG_FILE._08975_  (.A1(\u_cpu.REG_FILE._02765_ ),
    .A2(\u_cpu.REG_FILE._04241_ ),
    .A3(\u_cpu.REG_FILE._04243_ ),
    .B1(\u_cpu.REG_FILE._04248_ ),
    .C1(\u_cpu.REG_FILE._03023_ ),
    .X(\u_cpu.REG_FILE._04249_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08976_  (.A(\u_cpu.REG_FILE.rf[31][28] ),
    .B_N(\u_cpu.REG_FILE._02970_ ),
    .X(\u_cpu.REG_FILE._04250_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08977_  (.A1(\u_cpu.REG_FILE.rf[30][28] ),
    .A2(\u_cpu.REG_FILE._02749_ ),
    .B1(\u_cpu.REG_FILE._02969_ ),
    .C1(\u_cpu.REG_FILE._04250_ ),
    .Y(\u_cpu.REG_FILE._04251_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08978_  (.A1(\u_cpu.REG_FILE.rf[28][28] ),
    .A2(\u_cpu.REG_FILE._02830_ ),
    .B1_N(\u_cpu.REG_FILE._02975_ ),
    .X(\u_cpu.REG_FILE._04252_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08979_  (.A1(\u_cpu.REG_FILE.rf[29][28] ),
    .A2(\u_cpu.REG_FILE._03002_ ),
    .B1(\u_cpu.REG_FILE._04252_ ),
    .Y(\u_cpu.REG_FILE._04253_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08980_  (.A(\u_cpu.REG_FILE._04251_ ),
    .B(\u_cpu.REG_FILE._04253_ ),
    .C(\u_cpu.REG_FILE._03006_ ),
    .Y(\u_cpu.REG_FILE._04254_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._08981_  (.A_N(\u_cpu.REG_FILE.rf[25][28] ),
    .B(\u_cpu.REG_FILE._03069_ ),
    .X(\u_cpu.REG_FILE._04255_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._08982_  (.A1(\u_cpu.REG_FILE.rf[24][28] ),
    .A2(\u_cpu.REG_FILE._03212_ ),
    .B1_N(\u_cpu.REG_FILE._03072_ ),
    .Y(\u_cpu.REG_FILE._04256_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08983_  (.A(\u_cpu.REG_FILE.rf[27][28] ),
    .B_N(\u_cpu.REG_FILE._03077_ ),
    .X(\u_cpu.REG_FILE._04257_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08984_  (.A1(\u_cpu.REG_FILE.rf[26][28] ),
    .A2(\u_cpu.REG_FILE._03075_ ),
    .B1(\u_cpu.REG_FILE._03137_ ),
    .C1(\u_cpu.REG_FILE._04257_ ),
    .Y(\u_cpu.REG_FILE._04258_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08985_  (.A1(\u_cpu.REG_FILE._04255_ ),
    .A2(\u_cpu.REG_FILE._04256_ ),
    .B1(\u_cpu.REG_FILE._02777_ ),
    .C1(\u_cpu.REG_FILE._04258_ ),
    .Y(\u_cpu.REG_FILE._04259_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._08986_  (.A1(\u_cpu.REG_FILE._04254_ ),
    .A2(\u_cpu.REG_FILE._04259_ ),
    .A3(\u_cpu.REG_FILE._03129_ ),
    .B1(\u_cpu.REG_FILE._02996_ ),
    .X(\u_cpu.REG_FILE._04260_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08987_  (.A(\u_cpu.REG_FILE.rf[14][28] ),
    .B(\u_cpu.REG_FILE._02950_ ),
    .Y(\u_cpu.REG_FILE._04261_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08988_  (.A1(\u_cpu.REG_FILE.rf[15][28] ),
    .A2(\u_cpu.REG_FILE._02960_ ),
    .B1(\u_cpu.REG_FILE._02961_ ),
    .Y(\u_cpu.REG_FILE._04262_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08989_  (.A1(\u_cpu.REG_FILE.rf[12][28] ),
    .A2(\u_cpu.REG_FILE._02860_ ),
    .B1_N(\u_cpu.REG_FILE._02861_ ),
    .X(\u_cpu.REG_FILE._04263_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08990_  (.A1(\u_cpu.REG_FILE.rf[13][28] ),
    .A2(\u_cpu.REG_FILE._02956_ ),
    .B1(\u_cpu.REG_FILE._04263_ ),
    .Y(\u_cpu.REG_FILE._04264_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08991_  (.A1(\u_cpu.REG_FILE._04261_ ),
    .A2(\u_cpu.REG_FILE._04262_ ),
    .B1(\u_cpu.REG_FILE._04264_ ),
    .C1(\u_cpu.REG_FILE._02963_ ),
    .Y(\u_cpu.REG_FILE._04265_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._08992_  (.A(\u_cpu.REG_FILE.rf[11][28] ),
    .B_N(\u_cpu.REG_FILE._03012_ ),
    .X(\u_cpu.REG_FILE._04266_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._08993_  (.A1(\u_cpu.REG_FILE.rf[10][28] ),
    .A2(\u_cpu.REG_FILE._02940_ ),
    .B1(\u_cpu.REG_FILE._02854_ ),
    .C1(\u_cpu.REG_FILE._04266_ ),
    .Y(\u_cpu.REG_FILE._04267_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._08994_  (.A1(\u_cpu.REG_FILE.rf[8][28] ),
    .A2(\u_cpu.REG_FILE._03090_ ),
    .B1_N(\u_cpu.REG_FILE._02798_ ),
    .X(\u_cpu.REG_FILE._04268_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._08995_  (.A1(\u_cpu.REG_FILE.rf[9][28] ),
    .A2(\u_cpu.REG_FILE._03136_ ),
    .B1(\u_cpu.REG_FILE._04268_ ),
    .Y(\u_cpu.REG_FILE._04269_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08996_  (.A(\u_cpu.REG_FILE._03135_ ),
    .B(\u_cpu.REG_FILE._04267_ ),
    .C(\u_cpu.REG_FILE._04269_ ),
    .Y(\u_cpu.REG_FILE._04270_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._08997_  (.A(\u_cpu.REG_FILE._04265_ ),
    .B(\u_cpu.REG_FILE._04270_ ),
    .C(\u_cpu.REG_FILE._03141_ ),
    .Y(\u_cpu.REG_FILE._04271_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._08998_  (.A(\u_cpu.REG_FILE.rf[4][28] ),
    .B(\u_cpu.REG_FILE._03025_ ),
    .Y(\u_cpu.REG_FILE._04272_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._08999_  (.A1(\u_cpu.REG_FILE._02568_ ),
    .A2(\u_cpu.REG_FILE._02968_ ),
    .B1(\u_cpu.REG_FILE._03403_ ),
    .C1(\u_cpu.REG_FILE._04272_ ),
    .Y(\u_cpu.REG_FILE._04273_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._09000_  (.A1(\u_cpu.REG_FILE.rf[6][28] ),
    .A2(\u_cpu.REG_FILE._02797_ ),
    .B1(\u_cpu.REG_FILE._02799_ ),
    .Y(\u_cpu.REG_FILE._04274_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._09001_  (.A_N(\u_cpu.REG_FILE.rf[7][28] ),
    .B(\u_cpu.REG_FILE._02801_ ),
    .X(\u_cpu.REG_FILE._04275_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._09002_  (.A1(\u_cpu.REG_FILE._04274_ ),
    .A2(\u_cpu.REG_FILE._04275_ ),
    .B1(\u_cpu.REG_FILE._02804_ ),
    .Y(\u_cpu.REG_FILE._04276_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._09003_  (.A(\u_cpu.REG_FILE.rf[0][28] ),
    .B(\u_cpu.REG_FILE._02780_ ),
    .Y(\u_cpu.REG_FILE._04277_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._09004_  (.A1(\u_cpu.REG_FILE.rf[1][28] ),
    .A2(\u_cpu.REG_FILE._02845_ ),
    .B1_N(\u_cpu.REG_FILE._02812_ ),
    .Y(\u_cpu.REG_FILE._04278_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._09005_  (.A(\u_cpu.REG_FILE.rf[2][28] ),
    .B(\u_cpu.REG_FILE._02792_ ),
    .X(\u_cpu.REG_FILE._04279_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09006_  (.A1(\u_cpu.REG_FILE.rf[3][28] ),
    .A2(\u_cpu.REG_FILE._03351_ ),
    .B1(\u_cpu.REG_FILE._02818_ ),
    .C1(\u_cpu.REG_FILE._04279_ ),
    .Y(\u_cpu.REG_FILE._04280_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09007_  (.A1(\u_cpu.REG_FILE._04277_ ),
    .A2(\u_cpu.REG_FILE._04278_ ),
    .B1(\u_cpu.REG_FILE._02814_ ),
    .C1(\u_cpu.REG_FILE._04280_ ),
    .Y(\u_cpu.REG_FILE._04281_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09008_  (.A1(\u_cpu.REG_FILE._04273_ ),
    .A2(\u_cpu.REG_FILE._04276_ ),
    .B1(\u_cpu.REG_FILE._02807_ ),
    .C1(\u_cpu.REG_FILE._04281_ ),
    .Y(\u_cpu.REG_FILE._04282_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._09009_  (.A(\u_cpu.REG_FILE._02994_ ),
    .B(\u_cpu.REG_FILE._04271_ ),
    .C(\u_cpu.REG_FILE._04282_ ),
    .Y(\u_cpu.REG_FILE._04283_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._09010_  (.A1(\u_cpu.REG_FILE._04249_ ),
    .A2(\u_cpu.REG_FILE._04260_ ),
    .B1(\u_cpu.REG_FILE._04283_ ),
    .C1(\u_cpu.REG_FILE._03925_ ),
    .X(\u_cpu.ALU.SrcB[28] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._09011_  (.A(\u_cpu.REG_FILE.rf[15][29] ),
    .B_N(\u_cpu.REG_FILE._02748_ ),
    .X(\u_cpu.REG_FILE._04284_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09012_  (.A1(\u_cpu.REG_FILE.rf[14][29] ),
    .A2(\u_cpu.REG_FILE._03418_ ),
    .B1(\u_cpu.REG_FILE._02752_ ),
    .C1(\u_cpu.REG_FILE._04284_ ),
    .Y(\u_cpu.REG_FILE._04285_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._09013_  (.A1(\u_cpu.REG_FILE.rf[12][29] ),
    .A2(\u_cpu.REG_FILE._02974_ ),
    .B1_N(\u_cpu.REG_FILE._02761_ ),
    .X(\u_cpu.REG_FILE._04286_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._09014_  (.A1(\u_cpu.REG_FILE.rf[13][29] ),
    .A2(\u_cpu.REG_FILE._02973_ ),
    .B1(\u_cpu.REG_FILE._04286_ ),
    .Y(\u_cpu.REG_FILE._04287_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._09015_  (.A(\u_cpu.REG_FILE._04285_ ),
    .B(\u_cpu.REG_FILE._04287_ ),
    .C(\u_cpu.REG_FILE._02978_ ),
    .Y(\u_cpu.REG_FILE._04288_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._09016_  (.A_N(\u_cpu.REG_FILE.rf[9][29] ),
    .B(\u_cpu.REG_FILE._02945_ ),
    .X(\u_cpu.REG_FILE._04289_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._09017_  (.A1(\u_cpu.REG_FILE.rf[8][29] ),
    .A2(\u_cpu.REG_FILE._02816_ ),
    .B1_N(\u_cpu.REG_FILE._02947_ ),
    .Y(\u_cpu.REG_FILE._04290_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._09018_  (.A(\u_cpu.REG_FILE.rf[11][29] ),
    .B_N(\u_cpu.REG_FILE._02986_ ),
    .X(\u_cpu.REG_FILE._04291_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09019_  (.A1(\u_cpu.REG_FILE.rf[10][29] ),
    .A2(\u_cpu.REG_FILE._02824_ ),
    .B1(\u_cpu.REG_FILE._02846_ ),
    .C1(\u_cpu.REG_FILE._04291_ ),
    .Y(\u_cpu.REG_FILE._04292_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09020_  (.A1(\u_cpu.REG_FILE._04289_ ),
    .A2(\u_cpu.REG_FILE._04290_ ),
    .B1(\u_cpu.REG_FILE._03062_ ),
    .C1(\u_cpu.REG_FILE._04292_ ),
    .Y(\u_cpu.REG_FILE._04293_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._09021_  (.A(\u_cpu.REG_FILE._04288_ ),
    .B(\u_cpu.REG_FILE._04293_ ),
    .C(\u_cpu.REG_FILE._03218_ ),
    .Y(\u_cpu.REG_FILE._04294_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._09022_  (.A1(\u_cpu.REG_FILE.rf[4][29] ),
    .A2(\u_cpu.REG_FILE._03815_ ),
    .B1_N(\u_cpu.REG_FILE._02954_ ),
    .Y(\u_cpu.REG_FILE._04295_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._09023_  (.A1(\u_cpu.REG_FILE._02616_ ),
    .A2(\u_cpu.REG_FILE._02946_ ),
    .B1(\u_cpu.REG_FILE._04295_ ),
    .Y(\u_cpu.REG_FILE._04296_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._09024_  (.A1(\u_cpu.REG_FILE.rf[6][29] ),
    .A2(\u_cpu.REG_FILE._03331_ ),
    .B1(\u_cpu.REG_FILE._03407_ ),
    .Y(\u_cpu.REG_FILE._04297_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._09025_  (.A_N(\u_cpu.REG_FILE.rf[7][29] ),
    .B(\u_cpu.REG_FILE._02808_ ),
    .X(\u_cpu.REG_FILE._04298_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._09026_  (.A1(\u_cpu.REG_FILE._04297_ ),
    .A2(\u_cpu.REG_FILE._04298_ ),
    .B1(\u_cpu.REG_FILE._03434_ ),
    .Y(\u_cpu.REG_FILE._04299_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._09027_  (.A_N(\u_cpu.REG_FILE.rf[1][29] ),
    .B(\u_cpu.REG_FILE._03530_ ),
    .X(\u_cpu.REG_FILE._04300_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._09028_  (.A1(\u_cpu.REG_FILE.rf[0][29] ),
    .A2(\u_cpu.REG_FILE._03287_ ),
    .B1_N(\u_cpu.REG_FILE._02794_ ),
    .Y(\u_cpu.REG_FILE._04301_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._09029_  (.A(\u_cpu.REG_FILE.rf[3][29] ),
    .B_N(\u_cpu.REG_FILE._03337_ ),
    .X(\u_cpu.REG_FILE._04302_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09030_  (.A1(\u_cpu.REG_FILE.rf[2][29] ),
    .A2(\u_cpu.REG_FILE._02903_ ),
    .B1(\u_cpu.REG_FILE._03026_ ),
    .C1(\u_cpu.REG_FILE._04302_ ),
    .Y(\u_cpu.REG_FILE._04303_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09031_  (.A1(\u_cpu.REG_FILE._04300_ ),
    .A2(\u_cpu.REG_FILE._04301_ ),
    .B1(\u_cpu.REG_FILE._02858_ ),
    .C1(\u_cpu.REG_FILE._04303_ ),
    .Y(\u_cpu.REG_FILE._04304_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09032_  (.A1(\u_cpu.REG_FILE._04296_ ),
    .A2(\u_cpu.REG_FILE._04299_ ),
    .B1(\u_cpu.REG_FILE._02965_ ),
    .C1(\u_cpu.REG_FILE._04304_ ),
    .Y(\u_cpu.REG_FILE._04305_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._09033_  (.A(\u_cpu.REG_FILE._04294_ ),
    .B(\u_cpu.REG_FILE._04305_ ),
    .Y(\u_cpu.REG_FILE._04306_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._09034_  (.A(\u_cpu.REG_FILE.rf[27][29] ),
    .B_N(\u_cpu.REG_FILE._02871_ ),
    .X(\u_cpu.REG_FILE._04307_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._09035_  (.A1(\u_cpu.REG_FILE.rf[26][29] ),
    .A2(\u_cpu.REG_FILE._02982_ ),
    .B1(\u_cpu.REG_FILE._03000_ ),
    .C1(\u_cpu.REG_FILE._04307_ ),
    .X(\u_cpu.REG_FILE._04308_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._09036_  (.A1(\u_cpu.REG_FILE.rf[24][29] ),
    .A2(\u_cpu.REG_FILE._03445_ ),
    .B1_N(\u_cpu.REG_FILE._02865_ ),
    .X(\u_cpu.REG_FILE._04309_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._09037_  (.A(\u_cpu.REG_FILE.rf[25][29] ),
    .B_N(\u_cpu.REG_FILE._02832_ ),
    .X(\u_cpu.REG_FILE._04310_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._09038_  (.A1(\u_cpu.REG_FILE._04309_ ),
    .A2(\u_cpu.REG_FILE._04310_ ),
    .B1(\u_cpu.REG_FILE._02764_ ),
    .X(\u_cpu.REG_FILE._04311_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._09039_  (.A1(\u_cpu.REG_FILE.rf[28][29] ),
    .A2(\u_cpu.REG_FILE._02837_ ),
    .B1_N(\u_cpu.REG_FILE._03201_ ),
    .Y(\u_cpu.REG_FILE._04312_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._09040_  (.A(\u_cpu.REG_FILE.rf[29][29] ),
    .B(\u_cpu.REG_FILE._02841_ ),
    .Y(\u_cpu.REG_FILE._04313_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._09041_  (.A(\u_cpu.REG_FILE.rf[30][29] ),
    .B(\u_cpu.REG_FILE._02916_ ),
    .Y(\u_cpu.REG_FILE._04314_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._09042_  (.A1(\u_cpu.REG_FILE.rf[31][29] ),
    .A2(\u_cpu.REG_FILE._02845_ ),
    .B1(\u_cpu.REG_FILE._02846_ ),
    .Y(\u_cpu.REG_FILE._04315_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._09043_  (.A1(\u_cpu.REG_FILE._04312_ ),
    .A2(\u_cpu.REG_FILE._04313_ ),
    .B1(\u_cpu.REG_FILE._04314_ ),
    .B2(\u_cpu.REG_FILE._04315_ ),
    .C1(\u_cpu.REG_FILE._02919_ ),
    .Y(\u_cpu.REG_FILE._04316_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09044_  (.A1(\u_cpu.REG_FILE._04308_ ),
    .A2(\u_cpu.REG_FILE._04311_ ),
    .B1(\u_cpu.REG_FILE._02992_ ),
    .C1(\u_cpu.REG_FILE._04316_ ),
    .Y(\u_cpu.REG_FILE._04317_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._09045_  (.A1(\u_cpu.REG_FILE.rf[18][29] ),
    .A2(\u_cpu.REG_FILE._03404_ ),
    .B1(\u_cpu.REG_FILE._03249_ ),
    .Y(\u_cpu.REG_FILE._04318_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._09046_  (.A(\u_cpu.REG_FILE.rf[19][29] ),
    .B(\u_cpu.REG_FILE._03037_ ),
    .Y(\u_cpu.REG_FILE._04319_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._09047_  (.A1(\u_cpu.REG_FILE.rf[16][29] ),
    .A2(\u_cpu.REG_FILE._03038_ ),
    .B1_N(\u_cpu.REG_FILE._03039_ ),
    .X(\u_cpu.REG_FILE._04320_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._09048_  (.A1(\u_cpu.REG_FILE.rf[17][29] ),
    .A2(\u_cpu.REG_FILE._03304_ ),
    .B1(\u_cpu.REG_FILE._04320_ ),
    .Y(\u_cpu.REG_FILE._04321_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09049_  (.A1(\u_cpu.REG_FILE._04318_ ),
    .A2(\u_cpu.REG_FILE._04319_ ),
    .B1(\u_cpu.REG_FILE._03292_ ),
    .C1(\u_cpu.REG_FILE._04321_ ),
    .Y(\u_cpu.REG_FILE._04322_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._09050_  (.A(\u_cpu.REG_FILE.rf[22][29] ),
    .B(\u_cpu.REG_FILE._02810_ ),
    .X(\u_cpu.REG_FILE._04323_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09051_  (.A1(\u_cpu.REG_FILE.rf[23][29] ),
    .A2(\u_cpu.REG_FILE._03132_ ),
    .B1(\u_cpu.REG_FILE._02782_ ),
    .C1(\u_cpu.REG_FILE._04323_ ),
    .Y(\u_cpu.REG_FILE._04324_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._09052_  (.A1(\u_cpu.REG_FILE.rf[20][29] ),
    .A2(\u_cpu.REG_FILE._03016_ ),
    .B1_N(\u_cpu.REG_FILE._03017_ ),
    .X(\u_cpu.REG_FILE._04325_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._09053_  (.A1(\u_cpu.REG_FILE.rf[21][29] ),
    .A2(\u_cpu.REG_FILE._03015_ ),
    .B1(\u_cpu.REG_FILE._04325_ ),
    .Y(\u_cpu.REG_FILE._04326_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._09054_  (.A(\u_cpu.REG_FILE._04324_ ),
    .B(\u_cpu.REG_FILE._04326_ ),
    .C(\u_cpu.REG_FILE._03074_ ),
    .Y(\u_cpu.REG_FILE._04327_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._09055_  (.A(\u_cpu.REG_FILE._02807_ ),
    .B(\u_cpu.REG_FILE._04322_ ),
    .C(\u_cpu.REG_FILE._04327_ ),
    .Y(\u_cpu.REG_FILE._04328_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._09056_  (.A(\u_cpu.REG_FILE._04317_ ),
    .B(\u_cpu.REG_FILE._04328_ ),
    .C(\u_cpu.REG_FILE._02745_ ),
    .Y(\u_cpu.REG_FILE._04329_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._09057_  (.A1(\u_cpu.REG_FILE._02878_ ),
    .A2(\u_cpu.REG_FILE._04306_ ),
    .B1(\u_cpu.REG_FILE._04329_ ),
    .C1(\u_cpu.REG_FILE._03925_ ),
    .X(\u_cpu.ALU.SrcB[29] ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._09058_  (.A1(\u_cpu.REG_FILE.rf[18][30] ),
    .A2(\u_cpu.REG_FILE._03653_ ),
    .B1(\u_cpu.REG_FILE._03298_ ),
    .Y(\u_cpu.REG_FILE._04330_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._09059_  (.A1(\u_cpu.REG_FILE._02685_ ),
    .A2(\u_cpu.REG_FILE._02791_ ),
    .B1(\u_cpu.REG_FILE._04330_ ),
    .Y(\u_cpu.REG_FILE._04331_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._09060_  (.A(\u_cpu.REG_FILE.rf[16][30] ),
    .B(\u_cpu.REG_FILE._03371_ ),
    .Y(\u_cpu.REG_FILE._04332_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu.REG_FILE._09061_  (.A1(\u_cpu.REG_FILE._02688_ ),
    .A2(\u_cpu.REG_FILE._02968_ ),
    .B1(\u_cpu.REG_FILE._03057_ ),
    .C1(\u_cpu.REG_FILE._04332_ ),
    .Y(\u_cpu.REG_FILE._04333_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._09062_  (.A1(\u_cpu.REG_FILE.rf[20][30] ),
    .A2(\u_cpu.REG_FILE._02853_ ),
    .B1_N(\u_cpu.REG_FILE._02838_ ),
    .Y(\u_cpu.REG_FILE._04334_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._09063_  (.A(\u_cpu.REG_FILE.rf[21][30] ),
    .B(\u_cpu.REG_FILE._02859_ ),
    .Y(\u_cpu.REG_FILE._04335_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._09064_  (.A(\u_cpu.REG_FILE.rf[22][30] ),
    .B(\u_cpu.REG_FILE._02987_ ),
    .Y(\u_cpu.REG_FILE._04336_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._09065_  (.A1(\u_cpu.REG_FILE.rf[23][30] ),
    .A2(\u_cpu.REG_FILE._03351_ ),
    .B1(\u_cpu.REG_FILE._03377_ ),
    .Y(\u_cpu.REG_FILE._04337_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._09066_  (.A1(\u_cpu.REG_FILE._04334_ ),
    .A2(\u_cpu.REG_FILE._04335_ ),
    .B1(\u_cpu.REG_FILE._04336_ ),
    .B2(\u_cpu.REG_FILE._04337_ ),
    .C1(\u_cpu.REG_FILE._02848_ ),
    .Y(\u_cpu.REG_FILE._04338_ ));
 sky130_fd_sc_hd__o311a_2 \u_cpu.REG_FILE._09067_  (.A1(\u_cpu.REG_FILE._02765_ ),
    .A2(\u_cpu.REG_FILE._04331_ ),
    .A3(\u_cpu.REG_FILE._04333_ ),
    .B1(\u_cpu.REG_FILE._04338_ ),
    .C1(\u_cpu.REG_FILE._03023_ ),
    .X(\u_cpu.REG_FILE._04339_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._09068_  (.A(\u_cpu.REG_FILE.rf[31][30] ),
    .B_N(\u_cpu.REG_FILE._02970_ ),
    .X(\u_cpu.REG_FILE._04340_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09069_  (.A1(\u_cpu.REG_FILE.rf[30][30] ),
    .A2(\u_cpu.REG_FILE._02749_ ),
    .B1(\u_cpu.REG_FILE._02969_ ),
    .C1(\u_cpu.REG_FILE._04340_ ),
    .Y(\u_cpu.REG_FILE._04341_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._09070_  (.A1(\u_cpu.REG_FILE.rf[28][30] ),
    .A2(\u_cpu.REG_FILE._02830_ ),
    .B1_N(\u_cpu.REG_FILE._02975_ ),
    .X(\u_cpu.REG_FILE._04342_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._09071_  (.A1(\u_cpu.REG_FILE.rf[29][30] ),
    .A2(\u_cpu.REG_FILE._03002_ ),
    .B1(\u_cpu.REG_FILE._04342_ ),
    .Y(\u_cpu.REG_FILE._04343_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._09072_  (.A(\u_cpu.REG_FILE._04341_ ),
    .B(\u_cpu.REG_FILE._04343_ ),
    .C(\u_cpu.REG_FILE._03006_ ),
    .Y(\u_cpu.REG_FILE._04344_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._09073_  (.A_N(\u_cpu.REG_FILE.rf[25][30] ),
    .B(\u_cpu.REG_FILE._03069_ ),
    .X(\u_cpu.REG_FILE._04345_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._09074_  (.A1(\u_cpu.REG_FILE.rf[24][30] ),
    .A2(\u_cpu.REG_FILE._03212_ ),
    .B1_N(\u_cpu.REG_FILE._03072_ ),
    .Y(\u_cpu.REG_FILE._04346_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._09075_  (.A(\u_cpu.REG_FILE.rf[27][30] ),
    .B_N(\u_cpu.REG_FILE._03077_ ),
    .X(\u_cpu.REG_FILE._04347_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09076_  (.A1(\u_cpu.REG_FILE.rf[26][30] ),
    .A2(\u_cpu.REG_FILE._03075_ ),
    .B1(\u_cpu.REG_FILE._03137_ ),
    .C1(\u_cpu.REG_FILE._04347_ ),
    .Y(\u_cpu.REG_FILE._04348_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09077_  (.A1(\u_cpu.REG_FILE._04345_ ),
    .A2(\u_cpu.REG_FILE._04346_ ),
    .B1(\u_cpu.REG_FILE._02777_ ),
    .C1(\u_cpu.REG_FILE._04348_ ),
    .Y(\u_cpu.REG_FILE._04349_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu.REG_FILE._09078_  (.A1(\u_cpu.REG_FILE._04344_ ),
    .A2(\u_cpu.REG_FILE._04349_ ),
    .A3(\u_cpu.REG_FILE._03021_ ),
    .B1(\u_cpu.REG_FILE._02996_ ),
    .X(\u_cpu.REG_FILE._04350_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._09079_  (.A(\u_cpu.REG_FILE.rf[12][30] ),
    .B(\u_cpu.REG_FILE._02950_ ),
    .Y(\u_cpu.REG_FILE._04351_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._09080_  (.A1(\u_cpu.REG_FILE.rf[13][30] ),
    .A2(\u_cpu.REG_FILE._03132_ ),
    .B1_N(\u_cpu.REG_FILE._02983_ ),
    .Y(\u_cpu.REG_FILE._04352_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._09081_  (.A(\u_cpu.REG_FILE.rf[14][30] ),
    .B(\u_cpu.REG_FILE._02867_ ),
    .X(\u_cpu.REG_FILE._04353_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09082_  (.A1(\u_cpu.REG_FILE.rf[15][30] ),
    .A2(\u_cpu.REG_FILE._02841_ ),
    .B1(\u_cpu.REG_FILE._03076_ ),
    .C1(\u_cpu.REG_FILE._04353_ ),
    .Y(\u_cpu.REG_FILE._04354_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09083_  (.A1(\u_cpu.REG_FILE._04351_ ),
    .A2(\u_cpu.REG_FILE._04352_ ),
    .B1(\u_cpu.REG_FILE._03042_ ),
    .C1(\u_cpu.REG_FILE._04354_ ),
    .Y(\u_cpu.REG_FILE._04355_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._09084_  (.A(\u_cpu.REG_FILE.rf[8][30] ),
    .B(\u_cpu.REG_FILE._03309_ ),
    .Y(\u_cpu.REG_FILE._04356_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._09085_  (.A_N(\u_cpu.REG_FILE.rf[9][30] ),
    .B(\u_cpu.REG_FILE._03311_ ),
    .X(\u_cpu.REG_FILE._04357_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._09086_  (.A(\u_cpu.REG_FILE.rf[11][30] ),
    .B_N(\u_cpu.REG_FILE._02852_ ),
    .X(\u_cpu.REG_FILE._04358_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09087_  (.A1(\u_cpu.REG_FILE.rf[10][30] ),
    .A2(\u_cpu.REG_FILE._02797_ ),
    .B1(\u_cpu.REG_FILE._03198_ ),
    .C1(\u_cpu.REG_FILE._04358_ ),
    .Y(\u_cpu.REG_FILE._04359_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._09088_  (.A1(\u_cpu.REG_FILE._03308_ ),
    .A2(\u_cpu.REG_FILE._04356_ ),
    .A3(\u_cpu.REG_FILE._04357_ ),
    .B1(\u_cpu.REG_FILE._03008_ ),
    .C1(\u_cpu.REG_FILE._04359_ ),
    .Y(\u_cpu.REG_FILE._04360_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._09089_  (.A(\u_cpu.REG_FILE._04355_ ),
    .B(\u_cpu.REG_FILE._04360_ ),
    .C(\u_cpu.REG_FILE._03141_ ),
    .Y(\u_cpu.REG_FILE._04361_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._09090_  (.A(\u_cpu.REG_FILE.rf[0][30] ),
    .B(\u_cpu.REG_FILE._03309_ ),
    .Y(\u_cpu.REG_FILE._04362_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._09091_  (.A_N(\u_cpu.REG_FILE.rf[1][30] ),
    .B(\u_cpu.REG_FILE._03311_ ),
    .X(\u_cpu.REG_FILE._04363_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._09092_  (.A(\u_cpu.REG_FILE.rf[3][30] ),
    .B_N(\u_cpu.REG_FILE._02852_ ),
    .X(\u_cpu.REG_FILE._04364_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09093_  (.A1(\u_cpu.REG_FILE.rf[2][30] ),
    .A2(\u_cpu.REG_FILE._02837_ ),
    .B1(\u_cpu.REG_FILE._03407_ ),
    .C1(\u_cpu.REG_FILE._04364_ ),
    .Y(\u_cpu.REG_FILE._04365_ ));
 sky130_fd_sc_hd__o311ai_2 \u_cpu.REG_FILE._09094_  (.A1(\u_cpu.REG_FILE._03308_ ),
    .A2(\u_cpu.REG_FILE._04362_ ),
    .A3(\u_cpu.REG_FILE._04363_ ),
    .B1(\u_cpu.REG_FILE._03008_ ),
    .C1(\u_cpu.REG_FILE._04365_ ),
    .Y(\u_cpu.REG_FILE._04366_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._09095_  (.A1(\u_cpu.REG_FILE.rf[4][30] ),
    .A2(\u_cpu.REG_FILE._02748_ ),
    .B1_N(\u_cpu.REG_FILE._02781_ ),
    .X(\u_cpu.REG_FILE._04367_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._09096_  (.A1(\u_cpu.REG_FILE.rf[5][30] ),
    .A2(\u_cpu.REG_FILE._03002_ ),
    .B1(\u_cpu.REG_FILE._04367_ ),
    .Y(\u_cpu.REG_FILE._04368_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu.REG_FILE._09097_  (.A1(\u_cpu.REG_FILE.rf[6][30] ),
    .A2(\u_cpu.REG_FILE._03003_ ),
    .B1(\u_cpu.REG_FILE._02751_ ),
    .X(\u_cpu.REG_FILE._04369_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._09098_  (.A1(\u_cpu.REG_FILE.rf[7][30] ),
    .A2(\u_cpu.REG_FILE._03037_ ),
    .B1(\u_cpu.REG_FILE._04369_ ),
    .Y(\u_cpu.REG_FILE._04370_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._09099_  (.A(\u_cpu.REG_FILE._04368_ ),
    .B(\u_cpu.REG_FILE._02875_ ),
    .C(\u_cpu.REG_FILE._04370_ ),
    .Y(\u_cpu.REG_FILE._04371_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._09100_  (.A(\u_cpu.REG_FILE._02851_ ),
    .B(\u_cpu.REG_FILE._04366_ ),
    .C(\u_cpu.REG_FILE._04371_ ),
    .Y(\u_cpu.REG_FILE._04372_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._09101_  (.A(\u_cpu.REG_FILE._02994_ ),
    .B(\u_cpu.REG_FILE._04361_ ),
    .C(\u_cpu.REG_FILE._04372_ ),
    .Y(\u_cpu.REG_FILE._04373_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._09102_  (.A1(\u_cpu.REG_FILE._04339_ ),
    .A2(\u_cpu.REG_FILE._04350_ ),
    .B1(\u_cpu.REG_FILE._04373_ ),
    .C1(\u_cpu.REG_FILE._02883_ ),
    .X(\u_cpu.ALU.SrcB[30] ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._09103_  (.A(\u_cpu.REG_FILE.rf[15][31] ),
    .B_N(\u_cpu.REG_FILE._02748_ ),
    .X(\u_cpu.REG_FILE._04374_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09104_  (.A1(\u_cpu.REG_FILE.rf[14][31] ),
    .A2(\u_cpu.REG_FILE._03418_ ),
    .B1(\u_cpu.REG_FILE._02752_ ),
    .C1(\u_cpu.REG_FILE._04374_ ),
    .Y(\u_cpu.REG_FILE._04375_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._09105_  (.A1(\u_cpu.REG_FILE.rf[12][31] ),
    .A2(\u_cpu.REG_FILE._02974_ ),
    .B1_N(\u_cpu.REG_FILE._02761_ ),
    .X(\u_cpu.REG_FILE._04376_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._09106_  (.A1(\u_cpu.REG_FILE.rf[13][31] ),
    .A2(\u_cpu.REG_FILE._02973_ ),
    .B1(\u_cpu.REG_FILE._04376_ ),
    .Y(\u_cpu.REG_FILE._04377_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._09107_  (.A(\u_cpu.REG_FILE._04375_ ),
    .B(\u_cpu.REG_FILE._04377_ ),
    .C(\u_cpu.REG_FILE._02978_ ),
    .Y(\u_cpu.REG_FILE._04378_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._09108_  (.A_N(\u_cpu.REG_FILE.rf[9][31] ),
    .B(\u_cpu.REG_FILE._02945_ ),
    .X(\u_cpu.REG_FILE._04379_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._09109_  (.A1(\u_cpu.REG_FILE.rf[8][31] ),
    .A2(\u_cpu.REG_FILE._02816_ ),
    .B1_N(\u_cpu.REG_FILE._02947_ ),
    .Y(\u_cpu.REG_FILE._04380_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._09110_  (.A(\u_cpu.REG_FILE.rf[11][31] ),
    .B_N(\u_cpu.REG_FILE._02986_ ),
    .X(\u_cpu.REG_FILE._04381_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09111_  (.A1(\u_cpu.REG_FILE.rf[10][31] ),
    .A2(\u_cpu.REG_FILE._02824_ ),
    .B1(\u_cpu.REG_FILE._02846_ ),
    .C1(\u_cpu.REG_FILE._04381_ ),
    .Y(\u_cpu.REG_FILE._04382_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09112_  (.A1(\u_cpu.REG_FILE._04379_ ),
    .A2(\u_cpu.REG_FILE._04380_ ),
    .B1(\u_cpu.REG_FILE._03062_ ),
    .C1(\u_cpu.REG_FILE._04382_ ),
    .Y(\u_cpu.REG_FILE._04383_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._09113_  (.A(\u_cpu.REG_FILE._04378_ ),
    .B(\u_cpu.REG_FILE._04383_ ),
    .C(\u_cpu.REG_FILE._03218_ ),
    .Y(\u_cpu.REG_FILE._04384_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._09114_  (.A1(\u_cpu.REG_FILE.rf[4][31] ),
    .A2(\u_cpu.REG_FILE._03815_ ),
    .B1_N(\u_cpu.REG_FILE._02954_ ),
    .Y(\u_cpu.REG_FILE._04385_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu.REG_FILE._09115_  (.A1(\u_cpu.REG_FILE._02709_ ),
    .A2(\u_cpu.REG_FILE._02946_ ),
    .B1(\u_cpu.REG_FILE._04385_ ),
    .Y(\u_cpu.REG_FILE._04386_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._09116_  (.A1(\u_cpu.REG_FILE.rf[6][31] ),
    .A2(\u_cpu.REG_FILE._03331_ ),
    .B1(\u_cpu.REG_FILE._03407_ ),
    .Y(\u_cpu.REG_FILE._04387_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._09117_  (.A_N(\u_cpu.REG_FILE.rf[7][31] ),
    .B(\u_cpu.REG_FILE._02808_ ),
    .X(\u_cpu.REG_FILE._04388_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._09118_  (.A1(\u_cpu.REG_FILE._04387_ ),
    .A2(\u_cpu.REG_FILE._04388_ ),
    .B1(\u_cpu.REG_FILE._03434_ ),
    .Y(\u_cpu.REG_FILE._04389_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu.REG_FILE._09119_  (.A_N(\u_cpu.REG_FILE.rf[1][31] ),
    .B(\u_cpu.REG_FILE._03530_ ),
    .X(\u_cpu.REG_FILE._04390_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._09120_  (.A1(\u_cpu.REG_FILE.rf[0][31] ),
    .A2(\u_cpu.REG_FILE._03287_ ),
    .B1_N(\u_cpu.REG_FILE._02794_ ),
    .Y(\u_cpu.REG_FILE._04391_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._09121_  (.A(\u_cpu.REG_FILE.rf[3][31] ),
    .B_N(\u_cpu.REG_FILE._03337_ ),
    .X(\u_cpu.REG_FILE._04392_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09122_  (.A1(\u_cpu.REG_FILE.rf[2][31] ),
    .A2(\u_cpu.REG_FILE._03025_ ),
    .B1(\u_cpu.REG_FILE._03026_ ),
    .C1(\u_cpu.REG_FILE._04392_ ),
    .Y(\u_cpu.REG_FILE._04393_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09123_  (.A1(\u_cpu.REG_FILE._04390_ ),
    .A2(\u_cpu.REG_FILE._04391_ ),
    .B1(\u_cpu.REG_FILE._02858_ ),
    .C1(\u_cpu.REG_FILE._04393_ ),
    .Y(\u_cpu.REG_FILE._04394_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09124_  (.A1(\u_cpu.REG_FILE._04386_ ),
    .A2(\u_cpu.REG_FILE._04389_ ),
    .B1(\u_cpu.REG_FILE._02965_ ),
    .C1(\u_cpu.REG_FILE._04394_ ),
    .Y(\u_cpu.REG_FILE._04395_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu.REG_FILE._09125_  (.A(\u_cpu.REG_FILE._04384_ ),
    .B(\u_cpu.REG_FILE._04395_ ),
    .Y(\u_cpu.REG_FILE._04396_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._09126_  (.A(\u_cpu.REG_FILE.rf[27][31] ),
    .B_N(\u_cpu.REG_FILE._02871_ ),
    .X(\u_cpu.REG_FILE._04397_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._09127_  (.A1(\u_cpu.REG_FILE.rf[26][31] ),
    .A2(\u_cpu.REG_FILE._02982_ ),
    .B1(\u_cpu.REG_FILE._03000_ ),
    .C1(\u_cpu.REG_FILE._04397_ ),
    .X(\u_cpu.REG_FILE._04398_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._09128_  (.A1(\u_cpu.REG_FILE.rf[24][31] ),
    .A2(\u_cpu.REG_FILE._03445_ ),
    .B1_N(\u_cpu.REG_FILE._02865_ ),
    .X(\u_cpu.REG_FILE._04399_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu.REG_FILE._09129_  (.A(\u_cpu.REG_FILE.rf[25][31] ),
    .B_N(\u_cpu.REG_FILE._03003_ ),
    .X(\u_cpu.REG_FILE._04400_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu.REG_FILE._09130_  (.A1(\u_cpu.REG_FILE._04399_ ),
    .A2(\u_cpu.REG_FILE._04400_ ),
    .B1(\u_cpu.REG_FILE._02764_ ),
    .X(\u_cpu.REG_FILE._04401_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu.REG_FILE._09131_  (.A1(\u_cpu.REG_FILE.rf[28][31] ),
    .A2(\u_cpu.REG_FILE._02837_ ),
    .B1_N(\u_cpu.REG_FILE._03201_ ),
    .Y(\u_cpu.REG_FILE._04402_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._09132_  (.A(\u_cpu.REG_FILE.rf[29][31] ),
    .B(\u_cpu.REG_FILE._02841_ ),
    .Y(\u_cpu.REG_FILE._04403_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._09133_  (.A(\u_cpu.REG_FILE.rf[30][31] ),
    .B(\u_cpu.REG_FILE._02916_ ),
    .Y(\u_cpu.REG_FILE._04404_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._09134_  (.A1(\u_cpu.REG_FILE.rf[31][31] ),
    .A2(\u_cpu.REG_FILE._02845_ ),
    .B1(\u_cpu.REG_FILE._02941_ ),
    .Y(\u_cpu.REG_FILE._04405_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu.REG_FILE._09135_  (.A1(\u_cpu.REG_FILE._04402_ ),
    .A2(\u_cpu.REG_FILE._04403_ ),
    .B1(\u_cpu.REG_FILE._04404_ ),
    .B2(\u_cpu.REG_FILE._04405_ ),
    .C1(\u_cpu.REG_FILE._02919_ ),
    .Y(\u_cpu.REG_FILE._04406_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09136_  (.A1(\u_cpu.REG_FILE._04398_ ),
    .A2(\u_cpu.REG_FILE._04401_ ),
    .B1(\u_cpu.REG_FILE._02992_ ),
    .C1(\u_cpu.REG_FILE._04406_ ),
    .Y(\u_cpu.REG_FILE._04407_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._09137_  (.A1(\u_cpu.REG_FILE.rf[18][31] ),
    .A2(\u_cpu.REG_FILE._03404_ ),
    .B1(\u_cpu.REG_FILE._03470_ ),
    .Y(\u_cpu.REG_FILE._04408_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._09138_  (.A(\u_cpu.REG_FILE.rf[19][31] ),
    .B(\u_cpu.REG_FILE._03037_ ),
    .Y(\u_cpu.REG_FILE._04409_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._09139_  (.A1(\u_cpu.REG_FILE.rf[16][31] ),
    .A2(\u_cpu.REG_FILE._03038_ ),
    .B1_N(\u_cpu.REG_FILE._03039_ ),
    .X(\u_cpu.REG_FILE._04410_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._09140_  (.A1(\u_cpu.REG_FILE.rf[17][31] ),
    .A2(\u_cpu.REG_FILE._03304_ ),
    .B1(\u_cpu.REG_FILE._04410_ ),
    .Y(\u_cpu.REG_FILE._04411_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09141_  (.A1(\u_cpu.REG_FILE._04408_ ),
    .A2(\u_cpu.REG_FILE._04409_ ),
    .B1(\u_cpu.REG_FILE._03292_ ),
    .C1(\u_cpu.REG_FILE._04411_ ),
    .Y(\u_cpu.REG_FILE._04412_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu.REG_FILE._09142_  (.A(\u_cpu.REG_FILE.rf[22][31] ),
    .B(\u_cpu.REG_FILE._02810_ ),
    .X(\u_cpu.REG_FILE._04413_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu.REG_FILE._09143_  (.A1(\u_cpu.REG_FILE.rf[23][31] ),
    .A2(\u_cpu.REG_FILE._03132_ ),
    .B1(\u_cpu.REG_FILE._02782_ ),
    .C1(\u_cpu.REG_FILE._04413_ ),
    .Y(\u_cpu.REG_FILE._04414_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu.REG_FILE._09144_  (.A1(\u_cpu.REG_FILE.rf[20][31] ),
    .A2(\u_cpu.REG_FILE._03016_ ),
    .B1_N(\u_cpu.REG_FILE._03017_ ),
    .X(\u_cpu.REG_FILE._04415_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu.REG_FILE._09145_  (.A1(\u_cpu.REG_FILE.rf[21][31] ),
    .A2(\u_cpu.REG_FILE._03015_ ),
    .B1(\u_cpu.REG_FILE._04415_ ),
    .Y(\u_cpu.REG_FILE._04416_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._09146_  (.A(\u_cpu.REG_FILE._04414_ ),
    .B(\u_cpu.REG_FILE._04416_ ),
    .C(\u_cpu.REG_FILE._03074_ ),
    .Y(\u_cpu.REG_FILE._04417_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._09147_  (.A(\u_cpu.REG_FILE._02807_ ),
    .B(\u_cpu.REG_FILE._04412_ ),
    .C(\u_cpu.REG_FILE._04417_ ),
    .Y(\u_cpu.REG_FILE._04418_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._09148_  (.A(\u_cpu.REG_FILE._04407_ ),
    .B(\u_cpu.REG_FILE._04418_ ),
    .C(\u_cpu.REG_FILE._02745_ ),
    .Y(\u_cpu.REG_FILE._04419_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu.REG_FILE._09149_  (.A1(\u_cpu.REG_FILE._02878_ ),
    .A2(\u_cpu.REG_FILE._04396_ ),
    .B1(\u_cpu.REG_FILE._04419_ ),
    .C1(\u_cpu.REG_FILE._02883_ ),
    .X(\u_cpu.ALU.SrcB[31] ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09150_  (.A(\u_cpu.REG_FILE.wd3[0] ),
    .X(\u_cpu.REG_FILE._04420_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09151_  (.A(\u_cpu.REG_FILE.a3[3] ),
    .X(\u_cpu.REG_FILE._04421_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09152_  (.A(\u_cpu.REG_FILE._04421_ ),
    .X(\u_cpu.REG_FILE._04422_ ));
 sky130_fd_sc_hd__and3b_2 \u_cpu.REG_FILE._09153_  (.A_N(\u_cpu.REG_FILE.a3[1] ),
    .B(\u_cpu.REG_FILE.a3[0] ),
    .C(\u_cpu.REG_FILE.we3 ),
    .X(\u_cpu.REG_FILE._04423_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09154_  (.A(\u_cpu.REG_FILE.a3[4] ),
    .X(\u_cpu.REG_FILE._04424_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09155_  (.A(\u_cpu.REG_FILE.a3[2] ),
    .X(\u_cpu.REG_FILE._04425_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._09156_  (.A(\u_cpu.REG_FILE._04424_ ),
    .B(\u_cpu.REG_FILE._04425_ ),
    .Y(\u_cpu.REG_FILE._04426_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.REG_FILE._09157_  (.A(\u_cpu.REG_FILE._04422_ ),
    .B(\u_cpu.REG_FILE._04423_ ),
    .C(\u_cpu.REG_FILE._04426_ ),
    .X(\u_cpu.REG_FILE._04427_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09158_  (.A(\u_cpu.REG_FILE._04427_ ),
    .X(\u_cpu.REG_FILE._04428_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09159_  (.A0(\u_cpu.REG_FILE.rf[9][0] ),
    .A1(\u_cpu.REG_FILE._04420_ ),
    .S(\u_cpu.REG_FILE._04428_ ),
    .X(\u_cpu.REG_FILE._04429_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09160_  (.A(\u_cpu.REG_FILE._04429_ ),
    .X(\u_cpu.REG_FILE._00000_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09161_  (.A(\u_cpu.REG_FILE.wd3[1] ),
    .X(\u_cpu.REG_FILE._04430_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09162_  (.A0(\u_cpu.REG_FILE.rf[9][1] ),
    .A1(\u_cpu.REG_FILE._04430_ ),
    .S(\u_cpu.REG_FILE._04428_ ),
    .X(\u_cpu.REG_FILE._04431_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09163_  (.A(\u_cpu.REG_FILE._04431_ ),
    .X(\u_cpu.REG_FILE._00001_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09164_  (.A(\u_cpu.REG_FILE.wd3[2] ),
    .X(\u_cpu.REG_FILE._04432_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09165_  (.A0(\u_cpu.REG_FILE.rf[9][2] ),
    .A1(\u_cpu.REG_FILE._04432_ ),
    .S(\u_cpu.REG_FILE._04428_ ),
    .X(\u_cpu.REG_FILE._04433_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09166_  (.A(\u_cpu.REG_FILE._04433_ ),
    .X(\u_cpu.REG_FILE._00002_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09167_  (.A(\u_cpu.REG_FILE.wd3[3] ),
    .X(\u_cpu.REG_FILE._04434_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09168_  (.A0(\u_cpu.REG_FILE.rf[9][3] ),
    .A1(\u_cpu.REG_FILE._04434_ ),
    .S(\u_cpu.REG_FILE._04428_ ),
    .X(\u_cpu.REG_FILE._04435_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09169_  (.A(\u_cpu.REG_FILE._04435_ ),
    .X(\u_cpu.REG_FILE._00003_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09170_  (.A(\u_cpu.REG_FILE.wd3[4] ),
    .X(\u_cpu.REG_FILE._04436_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09171_  (.A0(\u_cpu.REG_FILE.rf[9][4] ),
    .A1(\u_cpu.REG_FILE._04436_ ),
    .S(\u_cpu.REG_FILE._04428_ ),
    .X(\u_cpu.REG_FILE._04437_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09172_  (.A(\u_cpu.REG_FILE._04437_ ),
    .X(\u_cpu.REG_FILE._00004_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09173_  (.A(\u_cpu.REG_FILE.wd3[5] ),
    .X(\u_cpu.REG_FILE._04438_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09174_  (.A0(\u_cpu.REG_FILE.rf[9][5] ),
    .A1(\u_cpu.REG_FILE._04438_ ),
    .S(\u_cpu.REG_FILE._04428_ ),
    .X(\u_cpu.REG_FILE._04439_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09175_  (.A(\u_cpu.REG_FILE._04439_ ),
    .X(\u_cpu.REG_FILE._00005_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09176_  (.A(\u_cpu.REG_FILE.wd3[6] ),
    .X(\u_cpu.REG_FILE._04440_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09177_  (.A0(\u_cpu.REG_FILE.rf[9][6] ),
    .A1(\u_cpu.REG_FILE._04440_ ),
    .S(\u_cpu.REG_FILE._04428_ ),
    .X(\u_cpu.REG_FILE._04441_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09178_  (.A(\u_cpu.REG_FILE._04441_ ),
    .X(\u_cpu.REG_FILE._00006_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09179_  (.A(\u_cpu.REG_FILE.wd3[7] ),
    .X(\u_cpu.REG_FILE._04442_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09180_  (.A0(\u_cpu.REG_FILE.rf[9][7] ),
    .A1(\u_cpu.REG_FILE._04442_ ),
    .S(\u_cpu.REG_FILE._04428_ ),
    .X(\u_cpu.REG_FILE._04443_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09181_  (.A(\u_cpu.REG_FILE._04443_ ),
    .X(\u_cpu.REG_FILE._00007_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09182_  (.A(\u_cpu.REG_FILE.wd3[8] ),
    .X(\u_cpu.REG_FILE._04444_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09183_  (.A0(\u_cpu.REG_FILE.rf[9][8] ),
    .A1(\u_cpu.REG_FILE._04444_ ),
    .S(\u_cpu.REG_FILE._04428_ ),
    .X(\u_cpu.REG_FILE._04445_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09184_  (.A(\u_cpu.REG_FILE._04445_ ),
    .X(\u_cpu.REG_FILE._00008_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09185_  (.A(\u_cpu.REG_FILE.wd3[9] ),
    .X(\u_cpu.REG_FILE._04446_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09186_  (.A0(\u_cpu.REG_FILE.rf[9][9] ),
    .A1(\u_cpu.REG_FILE._04446_ ),
    .S(\u_cpu.REG_FILE._04428_ ),
    .X(\u_cpu.REG_FILE._04447_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09187_  (.A(\u_cpu.REG_FILE._04447_ ),
    .X(\u_cpu.REG_FILE._00009_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09188_  (.A(\u_cpu.REG_FILE.wd3[10] ),
    .X(\u_cpu.REG_FILE._04448_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09189_  (.A(\u_cpu.REG_FILE._04427_ ),
    .X(\u_cpu.REG_FILE._04449_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09190_  (.A0(\u_cpu.REG_FILE.rf[9][10] ),
    .A1(\u_cpu.REG_FILE._04448_ ),
    .S(\u_cpu.REG_FILE._04449_ ),
    .X(\u_cpu.REG_FILE._04450_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09191_  (.A(\u_cpu.REG_FILE._04450_ ),
    .X(\u_cpu.REG_FILE._00010_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09192_  (.A(\u_cpu.REG_FILE.wd3[11] ),
    .X(\u_cpu.REG_FILE._04451_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09193_  (.A0(\u_cpu.REG_FILE.rf[9][11] ),
    .A1(\u_cpu.REG_FILE._04451_ ),
    .S(\u_cpu.REG_FILE._04449_ ),
    .X(\u_cpu.REG_FILE._04452_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09194_  (.A(\u_cpu.REG_FILE._04452_ ),
    .X(\u_cpu.REG_FILE._00011_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09195_  (.A(\u_cpu.REG_FILE.wd3[12] ),
    .X(\u_cpu.REG_FILE._04453_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09196_  (.A0(\u_cpu.REG_FILE.rf[9][12] ),
    .A1(\u_cpu.REG_FILE._04453_ ),
    .S(\u_cpu.REG_FILE._04449_ ),
    .X(\u_cpu.REG_FILE._04454_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09197_  (.A(\u_cpu.REG_FILE._04454_ ),
    .X(\u_cpu.REG_FILE._00012_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09198_  (.A(\u_cpu.REG_FILE.wd3[13] ),
    .X(\u_cpu.REG_FILE._04455_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09199_  (.A0(\u_cpu.REG_FILE.rf[9][13] ),
    .A1(\u_cpu.REG_FILE._04455_ ),
    .S(\u_cpu.REG_FILE._04449_ ),
    .X(\u_cpu.REG_FILE._04456_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09200_  (.A(\u_cpu.REG_FILE._04456_ ),
    .X(\u_cpu.REG_FILE._00013_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09201_  (.A(\u_cpu.REG_FILE.wd3[14] ),
    .X(\u_cpu.REG_FILE._04457_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09202_  (.A0(\u_cpu.REG_FILE.rf[9][14] ),
    .A1(\u_cpu.REG_FILE._04457_ ),
    .S(\u_cpu.REG_FILE._04449_ ),
    .X(\u_cpu.REG_FILE._04458_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09203_  (.A(\u_cpu.REG_FILE._04458_ ),
    .X(\u_cpu.REG_FILE._00014_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09204_  (.A(\u_cpu.REG_FILE.wd3[15] ),
    .X(\u_cpu.REG_FILE._04459_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09205_  (.A0(\u_cpu.REG_FILE.rf[9][15] ),
    .A1(\u_cpu.REG_FILE._04459_ ),
    .S(\u_cpu.REG_FILE._04449_ ),
    .X(\u_cpu.REG_FILE._04460_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09206_  (.A(\u_cpu.REG_FILE._04460_ ),
    .X(\u_cpu.REG_FILE._00015_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09207_  (.A(\u_cpu.REG_FILE.wd3[16] ),
    .X(\u_cpu.REG_FILE._04461_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09208_  (.A0(\u_cpu.REG_FILE.rf[9][16] ),
    .A1(\u_cpu.REG_FILE._04461_ ),
    .S(\u_cpu.REG_FILE._04449_ ),
    .X(\u_cpu.REG_FILE._04462_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09209_  (.A(\u_cpu.REG_FILE._04462_ ),
    .X(\u_cpu.REG_FILE._00016_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09210_  (.A(\u_cpu.REG_FILE.wd3[17] ),
    .X(\u_cpu.REG_FILE._04463_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09211_  (.A0(\u_cpu.REG_FILE.rf[9][17] ),
    .A1(\u_cpu.REG_FILE._04463_ ),
    .S(\u_cpu.REG_FILE._04449_ ),
    .X(\u_cpu.REG_FILE._04464_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09212_  (.A(\u_cpu.REG_FILE._04464_ ),
    .X(\u_cpu.REG_FILE._00017_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09213_  (.A(\u_cpu.REG_FILE.wd3[18] ),
    .X(\u_cpu.REG_FILE._04465_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09214_  (.A0(\u_cpu.REG_FILE.rf[9][18] ),
    .A1(\u_cpu.REG_FILE._04465_ ),
    .S(\u_cpu.REG_FILE._04449_ ),
    .X(\u_cpu.REG_FILE._04466_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09215_  (.A(\u_cpu.REG_FILE._04466_ ),
    .X(\u_cpu.REG_FILE._00018_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09216_  (.A(\u_cpu.REG_FILE.wd3[19] ),
    .X(\u_cpu.REG_FILE._04467_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09217_  (.A0(\u_cpu.REG_FILE.rf[9][19] ),
    .A1(\u_cpu.REG_FILE._04467_ ),
    .S(\u_cpu.REG_FILE._04449_ ),
    .X(\u_cpu.REG_FILE._04468_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09218_  (.A(\u_cpu.REG_FILE._04468_ ),
    .X(\u_cpu.REG_FILE._00019_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09219_  (.A(\u_cpu.REG_FILE.wd3[20] ),
    .X(\u_cpu.REG_FILE._04469_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09220_  (.A(\u_cpu.REG_FILE._04427_ ),
    .X(\u_cpu.REG_FILE._04470_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09221_  (.A0(\u_cpu.REG_FILE.rf[9][20] ),
    .A1(\u_cpu.REG_FILE._04469_ ),
    .S(\u_cpu.REG_FILE._04470_ ),
    .X(\u_cpu.REG_FILE._04471_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09222_  (.A(\u_cpu.REG_FILE._04471_ ),
    .X(\u_cpu.REG_FILE._00020_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09223_  (.A(\u_cpu.REG_FILE.wd3[21] ),
    .X(\u_cpu.REG_FILE._04472_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09224_  (.A0(\u_cpu.REG_FILE.rf[9][21] ),
    .A1(\u_cpu.REG_FILE._04472_ ),
    .S(\u_cpu.REG_FILE._04470_ ),
    .X(\u_cpu.REG_FILE._04473_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09225_  (.A(\u_cpu.REG_FILE._04473_ ),
    .X(\u_cpu.REG_FILE._00021_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09226_  (.A(\u_cpu.REG_FILE.wd3[22] ),
    .X(\u_cpu.REG_FILE._04474_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09227_  (.A0(\u_cpu.REG_FILE.rf[9][22] ),
    .A1(\u_cpu.REG_FILE._04474_ ),
    .S(\u_cpu.REG_FILE._04470_ ),
    .X(\u_cpu.REG_FILE._04475_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09228_  (.A(\u_cpu.REG_FILE._04475_ ),
    .X(\u_cpu.REG_FILE._00022_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09229_  (.A(\u_cpu.REG_FILE.wd3[23] ),
    .X(\u_cpu.REG_FILE._04476_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09230_  (.A0(\u_cpu.REG_FILE.rf[9][23] ),
    .A1(\u_cpu.REG_FILE._04476_ ),
    .S(\u_cpu.REG_FILE._04470_ ),
    .X(\u_cpu.REG_FILE._04477_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09231_  (.A(\u_cpu.REG_FILE._04477_ ),
    .X(\u_cpu.REG_FILE._00023_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09232_  (.A(\u_cpu.REG_FILE.wd3[24] ),
    .X(\u_cpu.REG_FILE._04478_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09233_  (.A0(\u_cpu.REG_FILE.rf[9][24] ),
    .A1(\u_cpu.REG_FILE._04478_ ),
    .S(\u_cpu.REG_FILE._04470_ ),
    .X(\u_cpu.REG_FILE._04479_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09234_  (.A(\u_cpu.REG_FILE._04479_ ),
    .X(\u_cpu.REG_FILE._00024_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09235_  (.A(\u_cpu.REG_FILE.wd3[25] ),
    .X(\u_cpu.REG_FILE._04480_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09236_  (.A0(\u_cpu.REG_FILE.rf[9][25] ),
    .A1(\u_cpu.REG_FILE._04480_ ),
    .S(\u_cpu.REG_FILE._04470_ ),
    .X(\u_cpu.REG_FILE._04481_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09237_  (.A(\u_cpu.REG_FILE._04481_ ),
    .X(\u_cpu.REG_FILE._00025_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09238_  (.A(\u_cpu.REG_FILE.wd3[26] ),
    .X(\u_cpu.REG_FILE._04482_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09239_  (.A0(\u_cpu.REG_FILE.rf[9][26] ),
    .A1(\u_cpu.REG_FILE._04482_ ),
    .S(\u_cpu.REG_FILE._04470_ ),
    .X(\u_cpu.REG_FILE._04483_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09240_  (.A(\u_cpu.REG_FILE._04483_ ),
    .X(\u_cpu.REG_FILE._00026_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09241_  (.A(\u_cpu.REG_FILE.wd3[27] ),
    .X(\u_cpu.REG_FILE._04484_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09242_  (.A0(\u_cpu.REG_FILE.rf[9][27] ),
    .A1(\u_cpu.REG_FILE._04484_ ),
    .S(\u_cpu.REG_FILE._04470_ ),
    .X(\u_cpu.REG_FILE._04485_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09243_  (.A(\u_cpu.REG_FILE._04485_ ),
    .X(\u_cpu.REG_FILE._00027_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09244_  (.A(\u_cpu.REG_FILE.wd3[28] ),
    .X(\u_cpu.REG_FILE._04486_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09245_  (.A0(\u_cpu.REG_FILE.rf[9][28] ),
    .A1(\u_cpu.REG_FILE._04486_ ),
    .S(\u_cpu.REG_FILE._04470_ ),
    .X(\u_cpu.REG_FILE._04487_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09246_  (.A(\u_cpu.REG_FILE._04487_ ),
    .X(\u_cpu.REG_FILE._00028_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09247_  (.A(\u_cpu.REG_FILE.wd3[29] ),
    .X(\u_cpu.REG_FILE._04488_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09248_  (.A0(\u_cpu.REG_FILE.rf[9][29] ),
    .A1(\u_cpu.REG_FILE._04488_ ),
    .S(\u_cpu.REG_FILE._04470_ ),
    .X(\u_cpu.REG_FILE._04489_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09249_  (.A(\u_cpu.REG_FILE._04489_ ),
    .X(\u_cpu.REG_FILE._00029_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09250_  (.A(\u_cpu.REG_FILE.wd3[30] ),
    .X(\u_cpu.REG_FILE._04490_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09251_  (.A0(\u_cpu.REG_FILE.rf[9][30] ),
    .A1(\u_cpu.REG_FILE._04490_ ),
    .S(\u_cpu.REG_FILE._04427_ ),
    .X(\u_cpu.REG_FILE._04491_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09252_  (.A(\u_cpu.REG_FILE._04491_ ),
    .X(\u_cpu.REG_FILE._00030_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09253_  (.A(\u_cpu.REG_FILE.wd3[31] ),
    .X(\u_cpu.REG_FILE._04492_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09254_  (.A0(\u_cpu.REG_FILE.rf[9][31] ),
    .A1(\u_cpu.REG_FILE._04492_ ),
    .S(\u_cpu.REG_FILE._04427_ ),
    .X(\u_cpu.REG_FILE._04493_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09255_  (.A(\u_cpu.REG_FILE._04493_ ),
    .X(\u_cpu.REG_FILE._00031_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09256_  (.A(\u_cpu.REG_FILE.a3[2] ),
    .X(\u_cpu.REG_FILE._04494_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.REG_FILE._09257_  (.A(\u_cpu.REG_FILE.a3[1] ),
    .B(\u_cpu.REG_FILE.a3[0] ),
    .C(\u_cpu.REG_FILE.we3 ),
    .X(\u_cpu.REG_FILE._04495_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09258_  (.A(\u_cpu.REG_FILE._04424_ ),
    .X(\u_cpu.REG_FILE._04496_ ));
 sky130_fd_sc_hd__or4bb_2 \u_cpu.REG_FILE._09259_  (.A(\u_cpu.REG_FILE._04422_ ),
    .B(\u_cpu.REG_FILE._04494_ ),
    .C_N(\u_cpu.REG_FILE._04495_ ),
    .D_N(\u_cpu.REG_FILE._04496_ ),
    .X(\u_cpu.REG_FILE._04497_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09260_  (.A(\u_cpu.REG_FILE._04497_ ),
    .X(\u_cpu.REG_FILE._04498_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09261_  (.A0(\u_cpu.REG_FILE._04420_ ),
    .A1(\u_cpu.REG_FILE.rf[19][0] ),
    .S(\u_cpu.REG_FILE._04498_ ),
    .X(\u_cpu.REG_FILE._04499_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09262_  (.A(\u_cpu.REG_FILE._04499_ ),
    .X(\u_cpu.REG_FILE._00032_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09263_  (.A0(\u_cpu.REG_FILE._04430_ ),
    .A1(\u_cpu.REG_FILE.rf[19][1] ),
    .S(\u_cpu.REG_FILE._04498_ ),
    .X(\u_cpu.REG_FILE._04500_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09264_  (.A(\u_cpu.REG_FILE._04500_ ),
    .X(\u_cpu.REG_FILE._00033_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09265_  (.A0(\u_cpu.REG_FILE._04432_ ),
    .A1(\u_cpu.REG_FILE.rf[19][2] ),
    .S(\u_cpu.REG_FILE._04498_ ),
    .X(\u_cpu.REG_FILE._04501_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09266_  (.A(\u_cpu.REG_FILE._04501_ ),
    .X(\u_cpu.REG_FILE._00034_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09267_  (.A0(\u_cpu.REG_FILE._04434_ ),
    .A1(\u_cpu.REG_FILE.rf[19][3] ),
    .S(\u_cpu.REG_FILE._04498_ ),
    .X(\u_cpu.REG_FILE._04502_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09268_  (.A(\u_cpu.REG_FILE._04502_ ),
    .X(\u_cpu.REG_FILE._00035_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09269_  (.A0(\u_cpu.REG_FILE._04436_ ),
    .A1(\u_cpu.REG_FILE.rf[19][4] ),
    .S(\u_cpu.REG_FILE._04498_ ),
    .X(\u_cpu.REG_FILE._04503_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09270_  (.A(\u_cpu.REG_FILE._04503_ ),
    .X(\u_cpu.REG_FILE._00036_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09271_  (.A0(\u_cpu.REG_FILE._04438_ ),
    .A1(\u_cpu.REG_FILE.rf[19][5] ),
    .S(\u_cpu.REG_FILE._04498_ ),
    .X(\u_cpu.REG_FILE._04504_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09272_  (.A(\u_cpu.REG_FILE._04504_ ),
    .X(\u_cpu.REG_FILE._00037_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09273_  (.A0(\u_cpu.REG_FILE._04440_ ),
    .A1(\u_cpu.REG_FILE.rf[19][6] ),
    .S(\u_cpu.REG_FILE._04498_ ),
    .X(\u_cpu.REG_FILE._04505_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09274_  (.A(\u_cpu.REG_FILE._04505_ ),
    .X(\u_cpu.REG_FILE._00038_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09275_  (.A0(\u_cpu.REG_FILE._04442_ ),
    .A1(\u_cpu.REG_FILE.rf[19][7] ),
    .S(\u_cpu.REG_FILE._04498_ ),
    .X(\u_cpu.REG_FILE._04506_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09276_  (.A(\u_cpu.REG_FILE._04506_ ),
    .X(\u_cpu.REG_FILE._00039_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09277_  (.A0(\u_cpu.REG_FILE._04444_ ),
    .A1(\u_cpu.REG_FILE.rf[19][8] ),
    .S(\u_cpu.REG_FILE._04498_ ),
    .X(\u_cpu.REG_FILE._04507_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09278_  (.A(\u_cpu.REG_FILE._04507_ ),
    .X(\u_cpu.REG_FILE._00040_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09279_  (.A0(\u_cpu.REG_FILE._04446_ ),
    .A1(\u_cpu.REG_FILE.rf[19][9] ),
    .S(\u_cpu.REG_FILE._04498_ ),
    .X(\u_cpu.REG_FILE._04508_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09280_  (.A(\u_cpu.REG_FILE._04508_ ),
    .X(\u_cpu.REG_FILE._00041_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09281_  (.A(\u_cpu.REG_FILE._04497_ ),
    .X(\u_cpu.REG_FILE._04509_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09282_  (.A0(\u_cpu.REG_FILE._04448_ ),
    .A1(\u_cpu.REG_FILE.rf[19][10] ),
    .S(\u_cpu.REG_FILE._04509_ ),
    .X(\u_cpu.REG_FILE._04510_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09283_  (.A(\u_cpu.REG_FILE._04510_ ),
    .X(\u_cpu.REG_FILE._00042_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09284_  (.A0(\u_cpu.REG_FILE._04451_ ),
    .A1(\u_cpu.REG_FILE.rf[19][11] ),
    .S(\u_cpu.REG_FILE._04509_ ),
    .X(\u_cpu.REG_FILE._04511_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09285_  (.A(\u_cpu.REG_FILE._04511_ ),
    .X(\u_cpu.REG_FILE._00043_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09286_  (.A0(\u_cpu.REG_FILE._04453_ ),
    .A1(\u_cpu.REG_FILE.rf[19][12] ),
    .S(\u_cpu.REG_FILE._04509_ ),
    .X(\u_cpu.REG_FILE._04512_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09287_  (.A(\u_cpu.REG_FILE._04512_ ),
    .X(\u_cpu.REG_FILE._00044_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09288_  (.A0(\u_cpu.REG_FILE._04455_ ),
    .A1(\u_cpu.REG_FILE.rf[19][13] ),
    .S(\u_cpu.REG_FILE._04509_ ),
    .X(\u_cpu.REG_FILE._04513_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09289_  (.A(\u_cpu.REG_FILE._04513_ ),
    .X(\u_cpu.REG_FILE._00045_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09290_  (.A0(\u_cpu.REG_FILE._04457_ ),
    .A1(\u_cpu.REG_FILE.rf[19][14] ),
    .S(\u_cpu.REG_FILE._04509_ ),
    .X(\u_cpu.REG_FILE._04514_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09291_  (.A(\u_cpu.REG_FILE._04514_ ),
    .X(\u_cpu.REG_FILE._00046_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09292_  (.A0(\u_cpu.REG_FILE._04459_ ),
    .A1(\u_cpu.REG_FILE.rf[19][15] ),
    .S(\u_cpu.REG_FILE._04509_ ),
    .X(\u_cpu.REG_FILE._04515_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09293_  (.A(\u_cpu.REG_FILE._04515_ ),
    .X(\u_cpu.REG_FILE._00047_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09294_  (.A0(\u_cpu.REG_FILE._04461_ ),
    .A1(\u_cpu.REG_FILE.rf[19][16] ),
    .S(\u_cpu.REG_FILE._04509_ ),
    .X(\u_cpu.REG_FILE._04516_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09295_  (.A(\u_cpu.REG_FILE._04516_ ),
    .X(\u_cpu.REG_FILE._00048_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09296_  (.A0(\u_cpu.REG_FILE._04463_ ),
    .A1(\u_cpu.REG_FILE.rf[19][17] ),
    .S(\u_cpu.REG_FILE._04509_ ),
    .X(\u_cpu.REG_FILE._04517_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09297_  (.A(\u_cpu.REG_FILE._04517_ ),
    .X(\u_cpu.REG_FILE._00049_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09298_  (.A0(\u_cpu.REG_FILE._04465_ ),
    .A1(\u_cpu.REG_FILE.rf[19][18] ),
    .S(\u_cpu.REG_FILE._04509_ ),
    .X(\u_cpu.REG_FILE._04518_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09299_  (.A(\u_cpu.REG_FILE._04518_ ),
    .X(\u_cpu.REG_FILE._00050_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09300_  (.A0(\u_cpu.REG_FILE._04467_ ),
    .A1(\u_cpu.REG_FILE.rf[19][19] ),
    .S(\u_cpu.REG_FILE._04509_ ),
    .X(\u_cpu.REG_FILE._04519_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09301_  (.A(\u_cpu.REG_FILE._04519_ ),
    .X(\u_cpu.REG_FILE._00051_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09302_  (.A(\u_cpu.REG_FILE._04497_ ),
    .X(\u_cpu.REG_FILE._04520_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09303_  (.A0(\u_cpu.REG_FILE._04469_ ),
    .A1(\u_cpu.REG_FILE.rf[19][20] ),
    .S(\u_cpu.REG_FILE._04520_ ),
    .X(\u_cpu.REG_FILE._04521_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09304_  (.A(\u_cpu.REG_FILE._04521_ ),
    .X(\u_cpu.REG_FILE._00052_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09305_  (.A0(\u_cpu.REG_FILE._04472_ ),
    .A1(\u_cpu.REG_FILE.rf[19][21] ),
    .S(\u_cpu.REG_FILE._04520_ ),
    .X(\u_cpu.REG_FILE._04522_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09306_  (.A(\u_cpu.REG_FILE._04522_ ),
    .X(\u_cpu.REG_FILE._00053_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09307_  (.A0(\u_cpu.REG_FILE._04474_ ),
    .A1(\u_cpu.REG_FILE.rf[19][22] ),
    .S(\u_cpu.REG_FILE._04520_ ),
    .X(\u_cpu.REG_FILE._04523_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09308_  (.A(\u_cpu.REG_FILE._04523_ ),
    .X(\u_cpu.REG_FILE._00054_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09309_  (.A0(\u_cpu.REG_FILE._04476_ ),
    .A1(\u_cpu.REG_FILE.rf[19][23] ),
    .S(\u_cpu.REG_FILE._04520_ ),
    .X(\u_cpu.REG_FILE._04524_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09310_  (.A(\u_cpu.REG_FILE._04524_ ),
    .X(\u_cpu.REG_FILE._00055_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09311_  (.A0(\u_cpu.REG_FILE._04478_ ),
    .A1(\u_cpu.REG_FILE.rf[19][24] ),
    .S(\u_cpu.REG_FILE._04520_ ),
    .X(\u_cpu.REG_FILE._04525_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09312_  (.A(\u_cpu.REG_FILE._04525_ ),
    .X(\u_cpu.REG_FILE._00056_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09313_  (.A0(\u_cpu.REG_FILE._04480_ ),
    .A1(\u_cpu.REG_FILE.rf[19][25] ),
    .S(\u_cpu.REG_FILE._04520_ ),
    .X(\u_cpu.REG_FILE._04526_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09314_  (.A(\u_cpu.REG_FILE._04526_ ),
    .X(\u_cpu.REG_FILE._00057_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09315_  (.A0(\u_cpu.REG_FILE._04482_ ),
    .A1(\u_cpu.REG_FILE.rf[19][26] ),
    .S(\u_cpu.REG_FILE._04520_ ),
    .X(\u_cpu.REG_FILE._04527_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09316_  (.A(\u_cpu.REG_FILE._04527_ ),
    .X(\u_cpu.REG_FILE._00058_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09317_  (.A0(\u_cpu.REG_FILE._04484_ ),
    .A1(\u_cpu.REG_FILE.rf[19][27] ),
    .S(\u_cpu.REG_FILE._04520_ ),
    .X(\u_cpu.REG_FILE._04528_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09318_  (.A(\u_cpu.REG_FILE._04528_ ),
    .X(\u_cpu.REG_FILE._00059_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09319_  (.A0(\u_cpu.REG_FILE._04486_ ),
    .A1(\u_cpu.REG_FILE.rf[19][28] ),
    .S(\u_cpu.REG_FILE._04520_ ),
    .X(\u_cpu.REG_FILE._04529_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09320_  (.A(\u_cpu.REG_FILE._04529_ ),
    .X(\u_cpu.REG_FILE._00060_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09321_  (.A0(\u_cpu.REG_FILE._04488_ ),
    .A1(\u_cpu.REG_FILE.rf[19][29] ),
    .S(\u_cpu.REG_FILE._04520_ ),
    .X(\u_cpu.REG_FILE._04530_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09322_  (.A(\u_cpu.REG_FILE._04530_ ),
    .X(\u_cpu.REG_FILE._00061_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09323_  (.A0(\u_cpu.REG_FILE._04490_ ),
    .A1(\u_cpu.REG_FILE.rf[19][30] ),
    .S(\u_cpu.REG_FILE._04497_ ),
    .X(\u_cpu.REG_FILE._04531_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09324_  (.A(\u_cpu.REG_FILE._04531_ ),
    .X(\u_cpu.REG_FILE._00062_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09325_  (.A0(\u_cpu.REG_FILE._04492_ ),
    .A1(\u_cpu.REG_FILE.rf[19][31] ),
    .S(\u_cpu.REG_FILE._04497_ ),
    .X(\u_cpu.REG_FILE._04532_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09326_  (.A(\u_cpu.REG_FILE._04532_ ),
    .X(\u_cpu.REG_FILE._00063_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.REG_FILE._09327_  (.A(\u_cpu.REG_FILE._04496_ ),
    .B(\u_cpu.REG_FILE._04422_ ),
    .C(\u_cpu.REG_FILE._04494_ ),
    .D(\u_cpu.REG_FILE._04423_ ),
    .X(\u_cpu.REG_FILE._04533_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09328_  (.A(\u_cpu.REG_FILE._04533_ ),
    .X(\u_cpu.REG_FILE._04534_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09329_  (.A0(\u_cpu.REG_FILE.rf[29][0] ),
    .A1(\u_cpu.REG_FILE._04420_ ),
    .S(\u_cpu.REG_FILE._04534_ ),
    .X(\u_cpu.REG_FILE._04535_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09330_  (.A(\u_cpu.REG_FILE._04535_ ),
    .X(\u_cpu.REG_FILE._00064_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09331_  (.A0(\u_cpu.REG_FILE.rf[29][1] ),
    .A1(\u_cpu.REG_FILE._04430_ ),
    .S(\u_cpu.REG_FILE._04534_ ),
    .X(\u_cpu.REG_FILE._04536_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09332_  (.A(\u_cpu.REG_FILE._04536_ ),
    .X(\u_cpu.REG_FILE._00065_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09333_  (.A0(\u_cpu.REG_FILE.rf[29][2] ),
    .A1(\u_cpu.REG_FILE._04432_ ),
    .S(\u_cpu.REG_FILE._04534_ ),
    .X(\u_cpu.REG_FILE._04537_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09334_  (.A(\u_cpu.REG_FILE._04537_ ),
    .X(\u_cpu.REG_FILE._00066_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09335_  (.A0(\u_cpu.REG_FILE.rf[29][3] ),
    .A1(\u_cpu.REG_FILE._04434_ ),
    .S(\u_cpu.REG_FILE._04534_ ),
    .X(\u_cpu.REG_FILE._04538_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09336_  (.A(\u_cpu.REG_FILE._04538_ ),
    .X(\u_cpu.REG_FILE._00067_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09337_  (.A0(\u_cpu.REG_FILE.rf[29][4] ),
    .A1(\u_cpu.REG_FILE._04436_ ),
    .S(\u_cpu.REG_FILE._04534_ ),
    .X(\u_cpu.REG_FILE._04539_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09338_  (.A(\u_cpu.REG_FILE._04539_ ),
    .X(\u_cpu.REG_FILE._00068_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09339_  (.A0(\u_cpu.REG_FILE.rf[29][5] ),
    .A1(\u_cpu.REG_FILE._04438_ ),
    .S(\u_cpu.REG_FILE._04534_ ),
    .X(\u_cpu.REG_FILE._04540_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09340_  (.A(\u_cpu.REG_FILE._04540_ ),
    .X(\u_cpu.REG_FILE._00069_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09341_  (.A0(\u_cpu.REG_FILE.rf[29][6] ),
    .A1(\u_cpu.REG_FILE._04440_ ),
    .S(\u_cpu.REG_FILE._04534_ ),
    .X(\u_cpu.REG_FILE._04541_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09342_  (.A(\u_cpu.REG_FILE._04541_ ),
    .X(\u_cpu.REG_FILE._00070_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09343_  (.A0(\u_cpu.REG_FILE.rf[29][7] ),
    .A1(\u_cpu.REG_FILE._04442_ ),
    .S(\u_cpu.REG_FILE._04534_ ),
    .X(\u_cpu.REG_FILE._04542_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09344_  (.A(\u_cpu.REG_FILE._04542_ ),
    .X(\u_cpu.REG_FILE._00071_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09345_  (.A0(\u_cpu.REG_FILE.rf[29][8] ),
    .A1(\u_cpu.REG_FILE._04444_ ),
    .S(\u_cpu.REG_FILE._04534_ ),
    .X(\u_cpu.REG_FILE._04543_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09346_  (.A(\u_cpu.REG_FILE._04543_ ),
    .X(\u_cpu.REG_FILE._00072_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09347_  (.A0(\u_cpu.REG_FILE.rf[29][9] ),
    .A1(\u_cpu.REG_FILE._04446_ ),
    .S(\u_cpu.REG_FILE._04534_ ),
    .X(\u_cpu.REG_FILE._04544_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09348_  (.A(\u_cpu.REG_FILE._04544_ ),
    .X(\u_cpu.REG_FILE._00073_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09349_  (.A(\u_cpu.REG_FILE._04533_ ),
    .X(\u_cpu.REG_FILE._04545_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09350_  (.A0(\u_cpu.REG_FILE.rf[29][10] ),
    .A1(\u_cpu.REG_FILE._04448_ ),
    .S(\u_cpu.REG_FILE._04545_ ),
    .X(\u_cpu.REG_FILE._04546_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09351_  (.A(\u_cpu.REG_FILE._04546_ ),
    .X(\u_cpu.REG_FILE._00074_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09352_  (.A0(\u_cpu.REG_FILE.rf[29][11] ),
    .A1(\u_cpu.REG_FILE._04451_ ),
    .S(\u_cpu.REG_FILE._04545_ ),
    .X(\u_cpu.REG_FILE._04547_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09353_  (.A(\u_cpu.REG_FILE._04547_ ),
    .X(\u_cpu.REG_FILE._00075_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09354_  (.A0(\u_cpu.REG_FILE.rf[29][12] ),
    .A1(\u_cpu.REG_FILE._04453_ ),
    .S(\u_cpu.REG_FILE._04545_ ),
    .X(\u_cpu.REG_FILE._04548_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09355_  (.A(\u_cpu.REG_FILE._04548_ ),
    .X(\u_cpu.REG_FILE._00076_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09356_  (.A0(\u_cpu.REG_FILE.rf[29][13] ),
    .A1(\u_cpu.REG_FILE._04455_ ),
    .S(\u_cpu.REG_FILE._04545_ ),
    .X(\u_cpu.REG_FILE._04549_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09357_  (.A(\u_cpu.REG_FILE._04549_ ),
    .X(\u_cpu.REG_FILE._00077_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09358_  (.A0(\u_cpu.REG_FILE.rf[29][14] ),
    .A1(\u_cpu.REG_FILE._04457_ ),
    .S(\u_cpu.REG_FILE._04545_ ),
    .X(\u_cpu.REG_FILE._04550_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09359_  (.A(\u_cpu.REG_FILE._04550_ ),
    .X(\u_cpu.REG_FILE._00078_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09360_  (.A0(\u_cpu.REG_FILE.rf[29][15] ),
    .A1(\u_cpu.REG_FILE._04459_ ),
    .S(\u_cpu.REG_FILE._04545_ ),
    .X(\u_cpu.REG_FILE._04551_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09361_  (.A(\u_cpu.REG_FILE._04551_ ),
    .X(\u_cpu.REG_FILE._00079_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09362_  (.A0(\u_cpu.REG_FILE.rf[29][16] ),
    .A1(\u_cpu.REG_FILE._04461_ ),
    .S(\u_cpu.REG_FILE._04545_ ),
    .X(\u_cpu.REG_FILE._04552_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09363_  (.A(\u_cpu.REG_FILE._04552_ ),
    .X(\u_cpu.REG_FILE._00080_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09364_  (.A0(\u_cpu.REG_FILE.rf[29][17] ),
    .A1(\u_cpu.REG_FILE._04463_ ),
    .S(\u_cpu.REG_FILE._04545_ ),
    .X(\u_cpu.REG_FILE._04553_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09365_  (.A(\u_cpu.REG_FILE._04553_ ),
    .X(\u_cpu.REG_FILE._00081_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09366_  (.A0(\u_cpu.REG_FILE.rf[29][18] ),
    .A1(\u_cpu.REG_FILE._04465_ ),
    .S(\u_cpu.REG_FILE._04545_ ),
    .X(\u_cpu.REG_FILE._04554_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09367_  (.A(\u_cpu.REG_FILE._04554_ ),
    .X(\u_cpu.REG_FILE._00082_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09368_  (.A0(\u_cpu.REG_FILE.rf[29][19] ),
    .A1(\u_cpu.REG_FILE._04467_ ),
    .S(\u_cpu.REG_FILE._04545_ ),
    .X(\u_cpu.REG_FILE._04555_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09369_  (.A(\u_cpu.REG_FILE._04555_ ),
    .X(\u_cpu.REG_FILE._00083_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09370_  (.A(\u_cpu.REG_FILE._04533_ ),
    .X(\u_cpu.REG_FILE._04556_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09371_  (.A0(\u_cpu.REG_FILE.rf[29][20] ),
    .A1(\u_cpu.REG_FILE._04469_ ),
    .S(\u_cpu.REG_FILE._04556_ ),
    .X(\u_cpu.REG_FILE._04557_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09372_  (.A(\u_cpu.REG_FILE._04557_ ),
    .X(\u_cpu.REG_FILE._00084_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09373_  (.A0(\u_cpu.REG_FILE.rf[29][21] ),
    .A1(\u_cpu.REG_FILE._04472_ ),
    .S(\u_cpu.REG_FILE._04556_ ),
    .X(\u_cpu.REG_FILE._04558_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09374_  (.A(\u_cpu.REG_FILE._04558_ ),
    .X(\u_cpu.REG_FILE._00085_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09375_  (.A0(\u_cpu.REG_FILE.rf[29][22] ),
    .A1(\u_cpu.REG_FILE._04474_ ),
    .S(\u_cpu.REG_FILE._04556_ ),
    .X(\u_cpu.REG_FILE._04559_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09376_  (.A(\u_cpu.REG_FILE._04559_ ),
    .X(\u_cpu.REG_FILE._00086_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09377_  (.A0(\u_cpu.REG_FILE.rf[29][23] ),
    .A1(\u_cpu.REG_FILE._04476_ ),
    .S(\u_cpu.REG_FILE._04556_ ),
    .X(\u_cpu.REG_FILE._04560_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09378_  (.A(\u_cpu.REG_FILE._04560_ ),
    .X(\u_cpu.REG_FILE._00087_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09379_  (.A0(\u_cpu.REG_FILE.rf[29][24] ),
    .A1(\u_cpu.REG_FILE._04478_ ),
    .S(\u_cpu.REG_FILE._04556_ ),
    .X(\u_cpu.REG_FILE._04561_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09380_  (.A(\u_cpu.REG_FILE._04561_ ),
    .X(\u_cpu.REG_FILE._00088_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09381_  (.A0(\u_cpu.REG_FILE.rf[29][25] ),
    .A1(\u_cpu.REG_FILE._04480_ ),
    .S(\u_cpu.REG_FILE._04556_ ),
    .X(\u_cpu.REG_FILE._04562_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09382_  (.A(\u_cpu.REG_FILE._04562_ ),
    .X(\u_cpu.REG_FILE._00089_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09383_  (.A0(\u_cpu.REG_FILE.rf[29][26] ),
    .A1(\u_cpu.REG_FILE._04482_ ),
    .S(\u_cpu.REG_FILE._04556_ ),
    .X(\u_cpu.REG_FILE._04563_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09384_  (.A(\u_cpu.REG_FILE._04563_ ),
    .X(\u_cpu.REG_FILE._00090_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09385_  (.A0(\u_cpu.REG_FILE.rf[29][27] ),
    .A1(\u_cpu.REG_FILE._04484_ ),
    .S(\u_cpu.REG_FILE._04556_ ),
    .X(\u_cpu.REG_FILE._04564_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09386_  (.A(\u_cpu.REG_FILE._04564_ ),
    .X(\u_cpu.REG_FILE._00091_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09387_  (.A0(\u_cpu.REG_FILE.rf[29][28] ),
    .A1(\u_cpu.REG_FILE._04486_ ),
    .S(\u_cpu.REG_FILE._04556_ ),
    .X(\u_cpu.REG_FILE._04565_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09388_  (.A(\u_cpu.REG_FILE._04565_ ),
    .X(\u_cpu.REG_FILE._00092_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09389_  (.A0(\u_cpu.REG_FILE.rf[29][29] ),
    .A1(\u_cpu.REG_FILE._04488_ ),
    .S(\u_cpu.REG_FILE._04556_ ),
    .X(\u_cpu.REG_FILE._04566_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09390_  (.A(\u_cpu.REG_FILE._04566_ ),
    .X(\u_cpu.REG_FILE._00093_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09391_  (.A0(\u_cpu.REG_FILE.rf[29][30] ),
    .A1(\u_cpu.REG_FILE._04490_ ),
    .S(\u_cpu.REG_FILE._04533_ ),
    .X(\u_cpu.REG_FILE._04567_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09392_  (.A(\u_cpu.REG_FILE._04567_ ),
    .X(\u_cpu.REG_FILE._00094_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09393_  (.A0(\u_cpu.REG_FILE.rf[29][31] ),
    .A1(\u_cpu.REG_FILE._04492_ ),
    .S(\u_cpu.REG_FILE._04533_ ),
    .X(\u_cpu.REG_FILE._04568_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09394_  (.A(\u_cpu.REG_FILE._04568_ ),
    .X(\u_cpu.REG_FILE._00095_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.REG_FILE._09395_  (.A(\u_cpu.REG_FILE._04496_ ),
    .B(\u_cpu.REG_FILE._04422_ ),
    .C(\u_cpu.REG_FILE._04494_ ),
    .D(\u_cpu.REG_FILE._04495_ ),
    .Y(\u_cpu.REG_FILE._04569_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09396_  (.A(\u_cpu.REG_FILE._04569_ ),
    .X(\u_cpu.REG_FILE._04570_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09397_  (.A0(\u_cpu.REG_FILE._04420_ ),
    .A1(\u_cpu.REG_FILE.rf[31][0] ),
    .S(\u_cpu.REG_FILE._04570_ ),
    .X(\u_cpu.REG_FILE._04571_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09398_  (.A(\u_cpu.REG_FILE._04571_ ),
    .X(\u_cpu.REG_FILE._00096_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09399_  (.A0(\u_cpu.REG_FILE._04430_ ),
    .A1(\u_cpu.REG_FILE.rf[31][1] ),
    .S(\u_cpu.REG_FILE._04570_ ),
    .X(\u_cpu.REG_FILE._04572_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09400_  (.A(\u_cpu.REG_FILE._04572_ ),
    .X(\u_cpu.REG_FILE._00097_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09401_  (.A0(\u_cpu.REG_FILE._04432_ ),
    .A1(\u_cpu.REG_FILE.rf[31][2] ),
    .S(\u_cpu.REG_FILE._04570_ ),
    .X(\u_cpu.REG_FILE._04573_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09402_  (.A(\u_cpu.REG_FILE._04573_ ),
    .X(\u_cpu.REG_FILE._00098_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09403_  (.A0(\u_cpu.REG_FILE._04434_ ),
    .A1(\u_cpu.REG_FILE.rf[31][3] ),
    .S(\u_cpu.REG_FILE._04570_ ),
    .X(\u_cpu.REG_FILE._04574_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09404_  (.A(\u_cpu.REG_FILE._04574_ ),
    .X(\u_cpu.REG_FILE._00099_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09405_  (.A0(\u_cpu.REG_FILE._04436_ ),
    .A1(\u_cpu.REG_FILE.rf[31][4] ),
    .S(\u_cpu.REG_FILE._04570_ ),
    .X(\u_cpu.REG_FILE._04575_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09406_  (.A(\u_cpu.REG_FILE._04575_ ),
    .X(\u_cpu.REG_FILE._00100_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09407_  (.A0(\u_cpu.REG_FILE._04438_ ),
    .A1(\u_cpu.REG_FILE.rf[31][5] ),
    .S(\u_cpu.REG_FILE._04570_ ),
    .X(\u_cpu.REG_FILE._04576_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09408_  (.A(\u_cpu.REG_FILE._04576_ ),
    .X(\u_cpu.REG_FILE._00101_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09409_  (.A0(\u_cpu.REG_FILE._04440_ ),
    .A1(\u_cpu.REG_FILE.rf[31][6] ),
    .S(\u_cpu.REG_FILE._04570_ ),
    .X(\u_cpu.REG_FILE._04577_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09410_  (.A(\u_cpu.REG_FILE._04577_ ),
    .X(\u_cpu.REG_FILE._00102_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09411_  (.A0(\u_cpu.REG_FILE._04442_ ),
    .A1(\u_cpu.REG_FILE.rf[31][7] ),
    .S(\u_cpu.REG_FILE._04570_ ),
    .X(\u_cpu.REG_FILE._04578_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09412_  (.A(\u_cpu.REG_FILE._04578_ ),
    .X(\u_cpu.REG_FILE._00103_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09413_  (.A0(\u_cpu.REG_FILE._04444_ ),
    .A1(\u_cpu.REG_FILE.rf[31][8] ),
    .S(\u_cpu.REG_FILE._04570_ ),
    .X(\u_cpu.REG_FILE._04579_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09414_  (.A(\u_cpu.REG_FILE._04579_ ),
    .X(\u_cpu.REG_FILE._00104_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09415_  (.A0(\u_cpu.REG_FILE._04446_ ),
    .A1(\u_cpu.REG_FILE.rf[31][9] ),
    .S(\u_cpu.REG_FILE._04570_ ),
    .X(\u_cpu.REG_FILE._04580_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09416_  (.A(\u_cpu.REG_FILE._04580_ ),
    .X(\u_cpu.REG_FILE._00105_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09417_  (.A(\u_cpu.REG_FILE._04569_ ),
    .X(\u_cpu.REG_FILE._04581_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09418_  (.A0(\u_cpu.REG_FILE._04448_ ),
    .A1(\u_cpu.REG_FILE.rf[31][10] ),
    .S(\u_cpu.REG_FILE._04581_ ),
    .X(\u_cpu.REG_FILE._04582_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09419_  (.A(\u_cpu.REG_FILE._04582_ ),
    .X(\u_cpu.REG_FILE._00106_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09420_  (.A0(\u_cpu.REG_FILE._04451_ ),
    .A1(\u_cpu.REG_FILE.rf[31][11] ),
    .S(\u_cpu.REG_FILE._04581_ ),
    .X(\u_cpu.REG_FILE._04583_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09421_  (.A(\u_cpu.REG_FILE._04583_ ),
    .X(\u_cpu.REG_FILE._00107_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09422_  (.A0(\u_cpu.REG_FILE._04453_ ),
    .A1(\u_cpu.REG_FILE.rf[31][12] ),
    .S(\u_cpu.REG_FILE._04581_ ),
    .X(\u_cpu.REG_FILE._04584_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09423_  (.A(\u_cpu.REG_FILE._04584_ ),
    .X(\u_cpu.REG_FILE._00108_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09424_  (.A0(\u_cpu.REG_FILE._04455_ ),
    .A1(\u_cpu.REG_FILE.rf[31][13] ),
    .S(\u_cpu.REG_FILE._04581_ ),
    .X(\u_cpu.REG_FILE._04585_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09425_  (.A(\u_cpu.REG_FILE._04585_ ),
    .X(\u_cpu.REG_FILE._00109_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09426_  (.A0(\u_cpu.REG_FILE._04457_ ),
    .A1(\u_cpu.REG_FILE.rf[31][14] ),
    .S(\u_cpu.REG_FILE._04581_ ),
    .X(\u_cpu.REG_FILE._04586_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09427_  (.A(\u_cpu.REG_FILE._04586_ ),
    .X(\u_cpu.REG_FILE._00110_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09428_  (.A0(\u_cpu.REG_FILE._04459_ ),
    .A1(\u_cpu.REG_FILE.rf[31][15] ),
    .S(\u_cpu.REG_FILE._04581_ ),
    .X(\u_cpu.REG_FILE._04587_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09429_  (.A(\u_cpu.REG_FILE._04587_ ),
    .X(\u_cpu.REG_FILE._00111_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09430_  (.A0(\u_cpu.REG_FILE._04461_ ),
    .A1(\u_cpu.REG_FILE.rf[31][16] ),
    .S(\u_cpu.REG_FILE._04581_ ),
    .X(\u_cpu.REG_FILE._04588_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09431_  (.A(\u_cpu.REG_FILE._04588_ ),
    .X(\u_cpu.REG_FILE._00112_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09432_  (.A0(\u_cpu.REG_FILE._04463_ ),
    .A1(\u_cpu.REG_FILE.rf[31][17] ),
    .S(\u_cpu.REG_FILE._04581_ ),
    .X(\u_cpu.REG_FILE._04589_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09433_  (.A(\u_cpu.REG_FILE._04589_ ),
    .X(\u_cpu.REG_FILE._00113_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09434_  (.A0(\u_cpu.REG_FILE._04465_ ),
    .A1(\u_cpu.REG_FILE.rf[31][18] ),
    .S(\u_cpu.REG_FILE._04581_ ),
    .X(\u_cpu.REG_FILE._04590_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09435_  (.A(\u_cpu.REG_FILE._04590_ ),
    .X(\u_cpu.REG_FILE._00114_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09436_  (.A0(\u_cpu.REG_FILE._04467_ ),
    .A1(\u_cpu.REG_FILE.rf[31][19] ),
    .S(\u_cpu.REG_FILE._04581_ ),
    .X(\u_cpu.REG_FILE._04591_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09437_  (.A(\u_cpu.REG_FILE._04591_ ),
    .X(\u_cpu.REG_FILE._00115_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09438_  (.A(\u_cpu.REG_FILE._04569_ ),
    .X(\u_cpu.REG_FILE._04592_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09439_  (.A0(\u_cpu.REG_FILE._04469_ ),
    .A1(\u_cpu.REG_FILE.rf[31][20] ),
    .S(\u_cpu.REG_FILE._04592_ ),
    .X(\u_cpu.REG_FILE._04593_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09440_  (.A(\u_cpu.REG_FILE._04593_ ),
    .X(\u_cpu.REG_FILE._00116_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09441_  (.A0(\u_cpu.REG_FILE._04472_ ),
    .A1(\u_cpu.REG_FILE.rf[31][21] ),
    .S(\u_cpu.REG_FILE._04592_ ),
    .X(\u_cpu.REG_FILE._04594_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09442_  (.A(\u_cpu.REG_FILE._04594_ ),
    .X(\u_cpu.REG_FILE._00117_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09443_  (.A0(\u_cpu.REG_FILE._04474_ ),
    .A1(\u_cpu.REG_FILE.rf[31][22] ),
    .S(\u_cpu.REG_FILE._04592_ ),
    .X(\u_cpu.REG_FILE._04595_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09444_  (.A(\u_cpu.REG_FILE._04595_ ),
    .X(\u_cpu.REG_FILE._00118_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09445_  (.A0(\u_cpu.REG_FILE._04476_ ),
    .A1(\u_cpu.REG_FILE.rf[31][23] ),
    .S(\u_cpu.REG_FILE._04592_ ),
    .X(\u_cpu.REG_FILE._04596_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09446_  (.A(\u_cpu.REG_FILE._04596_ ),
    .X(\u_cpu.REG_FILE._00119_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09447_  (.A0(\u_cpu.REG_FILE._04478_ ),
    .A1(\u_cpu.REG_FILE.rf[31][24] ),
    .S(\u_cpu.REG_FILE._04592_ ),
    .X(\u_cpu.REG_FILE._04597_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09448_  (.A(\u_cpu.REG_FILE._04597_ ),
    .X(\u_cpu.REG_FILE._00120_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09449_  (.A0(\u_cpu.REG_FILE._04480_ ),
    .A1(\u_cpu.REG_FILE.rf[31][25] ),
    .S(\u_cpu.REG_FILE._04592_ ),
    .X(\u_cpu.REG_FILE._04598_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09450_  (.A(\u_cpu.REG_FILE._04598_ ),
    .X(\u_cpu.REG_FILE._00121_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09451_  (.A0(\u_cpu.REG_FILE._04482_ ),
    .A1(\u_cpu.REG_FILE.rf[31][26] ),
    .S(\u_cpu.REG_FILE._04592_ ),
    .X(\u_cpu.REG_FILE._04599_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09452_  (.A(\u_cpu.REG_FILE._04599_ ),
    .X(\u_cpu.REG_FILE._00122_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09453_  (.A0(\u_cpu.REG_FILE._04484_ ),
    .A1(\u_cpu.REG_FILE.rf[31][27] ),
    .S(\u_cpu.REG_FILE._04592_ ),
    .X(\u_cpu.REG_FILE._04600_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09454_  (.A(\u_cpu.REG_FILE._04600_ ),
    .X(\u_cpu.REG_FILE._00123_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09455_  (.A0(\u_cpu.REG_FILE._04486_ ),
    .A1(\u_cpu.REG_FILE.rf[31][28] ),
    .S(\u_cpu.REG_FILE._04592_ ),
    .X(\u_cpu.REG_FILE._04601_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09456_  (.A(\u_cpu.REG_FILE._04601_ ),
    .X(\u_cpu.REG_FILE._00124_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09457_  (.A0(\u_cpu.REG_FILE._04488_ ),
    .A1(\u_cpu.REG_FILE.rf[31][29] ),
    .S(\u_cpu.REG_FILE._04592_ ),
    .X(\u_cpu.REG_FILE._04602_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09458_  (.A(\u_cpu.REG_FILE._04602_ ),
    .X(\u_cpu.REG_FILE._00125_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09459_  (.A0(\u_cpu.REG_FILE._04490_ ),
    .A1(\u_cpu.REG_FILE.rf[31][30] ),
    .S(\u_cpu.REG_FILE._04569_ ),
    .X(\u_cpu.REG_FILE._04603_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09460_  (.A(\u_cpu.REG_FILE._04603_ ),
    .X(\u_cpu.REG_FILE._00126_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09461_  (.A0(\u_cpu.REG_FILE._04492_ ),
    .A1(\u_cpu.REG_FILE.rf[31][31] ),
    .S(\u_cpu.REG_FILE._04569_ ),
    .X(\u_cpu.REG_FILE._04604_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09462_  (.A(\u_cpu.REG_FILE._04604_ ),
    .X(\u_cpu.REG_FILE._00127_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu.REG_FILE._09463_  (.A(\u_cpu.REG_FILE.a3[4] ),
    .B(\u_cpu.REG_FILE.a3[3] ),
    .C(\u_cpu.REG_FILE.a3[2] ),
    .Y(\u_cpu.REG_FILE._04605_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.REG_FILE._09464_  (.A(\u_cpu.REG_FILE.a3[1] ),
    .B(\u_cpu.REG_FILE.a3[0] ),
    .C(\u_cpu.REG_FILE.we3 ),
    .D(\u_cpu.REG_FILE._04605_ ),
    .X(\u_cpu.REG_FILE._04606_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09465_  (.A(\u_cpu.REG_FILE._04606_ ),
    .X(\u_cpu.REG_FILE._04607_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09466_  (.A0(\u_cpu.REG_FILE.rf[3][0] ),
    .A1(\u_cpu.REG_FILE._04420_ ),
    .S(\u_cpu.REG_FILE._04607_ ),
    .X(\u_cpu.REG_FILE._04608_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09467_  (.A(\u_cpu.REG_FILE._04608_ ),
    .X(\u_cpu.REG_FILE._00128_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09468_  (.A0(\u_cpu.REG_FILE.rf[3][1] ),
    .A1(\u_cpu.REG_FILE._04430_ ),
    .S(\u_cpu.REG_FILE._04607_ ),
    .X(\u_cpu.REG_FILE._04609_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09469_  (.A(\u_cpu.REG_FILE._04609_ ),
    .X(\u_cpu.REG_FILE._00129_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09470_  (.A0(\u_cpu.REG_FILE.rf[3][2] ),
    .A1(\u_cpu.REG_FILE._04432_ ),
    .S(\u_cpu.REG_FILE._04607_ ),
    .X(\u_cpu.REG_FILE._04610_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09471_  (.A(\u_cpu.REG_FILE._04610_ ),
    .X(\u_cpu.REG_FILE._00130_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09472_  (.A0(\u_cpu.REG_FILE.rf[3][3] ),
    .A1(\u_cpu.REG_FILE._04434_ ),
    .S(\u_cpu.REG_FILE._04607_ ),
    .X(\u_cpu.REG_FILE._04611_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09473_  (.A(\u_cpu.REG_FILE._04611_ ),
    .X(\u_cpu.REG_FILE._00131_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09474_  (.A0(\u_cpu.REG_FILE.rf[3][4] ),
    .A1(\u_cpu.REG_FILE._04436_ ),
    .S(\u_cpu.REG_FILE._04607_ ),
    .X(\u_cpu.REG_FILE._04612_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09475_  (.A(\u_cpu.REG_FILE._04612_ ),
    .X(\u_cpu.REG_FILE._00132_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09476_  (.A0(\u_cpu.REG_FILE.rf[3][5] ),
    .A1(\u_cpu.REG_FILE._04438_ ),
    .S(\u_cpu.REG_FILE._04607_ ),
    .X(\u_cpu.REG_FILE._04613_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09477_  (.A(\u_cpu.REG_FILE._04613_ ),
    .X(\u_cpu.REG_FILE._00133_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09478_  (.A0(\u_cpu.REG_FILE.rf[3][6] ),
    .A1(\u_cpu.REG_FILE._04440_ ),
    .S(\u_cpu.REG_FILE._04607_ ),
    .X(\u_cpu.REG_FILE._04614_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09479_  (.A(\u_cpu.REG_FILE._04614_ ),
    .X(\u_cpu.REG_FILE._00134_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09480_  (.A0(\u_cpu.REG_FILE.rf[3][7] ),
    .A1(\u_cpu.REG_FILE._04442_ ),
    .S(\u_cpu.REG_FILE._04607_ ),
    .X(\u_cpu.REG_FILE._04615_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09481_  (.A(\u_cpu.REG_FILE._04615_ ),
    .X(\u_cpu.REG_FILE._00135_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09482_  (.A0(\u_cpu.REG_FILE.rf[3][8] ),
    .A1(\u_cpu.REG_FILE._04444_ ),
    .S(\u_cpu.REG_FILE._04607_ ),
    .X(\u_cpu.REG_FILE._04616_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09483_  (.A(\u_cpu.REG_FILE._04616_ ),
    .X(\u_cpu.REG_FILE._00136_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09484_  (.A0(\u_cpu.REG_FILE.rf[3][9] ),
    .A1(\u_cpu.REG_FILE._04446_ ),
    .S(\u_cpu.REG_FILE._04607_ ),
    .X(\u_cpu.REG_FILE._04617_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09485_  (.A(\u_cpu.REG_FILE._04617_ ),
    .X(\u_cpu.REG_FILE._00137_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09486_  (.A(\u_cpu.REG_FILE._04606_ ),
    .X(\u_cpu.REG_FILE._04618_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09487_  (.A0(\u_cpu.REG_FILE.rf[3][10] ),
    .A1(\u_cpu.REG_FILE._04448_ ),
    .S(\u_cpu.REG_FILE._04618_ ),
    .X(\u_cpu.REG_FILE._04619_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09488_  (.A(\u_cpu.REG_FILE._04619_ ),
    .X(\u_cpu.REG_FILE._00138_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09489_  (.A0(\u_cpu.REG_FILE.rf[3][11] ),
    .A1(\u_cpu.REG_FILE._04451_ ),
    .S(\u_cpu.REG_FILE._04618_ ),
    .X(\u_cpu.REG_FILE._04620_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09490_  (.A(\u_cpu.REG_FILE._04620_ ),
    .X(\u_cpu.REG_FILE._00139_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09491_  (.A0(\u_cpu.REG_FILE.rf[3][12] ),
    .A1(\u_cpu.REG_FILE._04453_ ),
    .S(\u_cpu.REG_FILE._04618_ ),
    .X(\u_cpu.REG_FILE._04621_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09492_  (.A(\u_cpu.REG_FILE._04621_ ),
    .X(\u_cpu.REG_FILE._00140_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09493_  (.A0(\u_cpu.REG_FILE.rf[3][13] ),
    .A1(\u_cpu.REG_FILE._04455_ ),
    .S(\u_cpu.REG_FILE._04618_ ),
    .X(\u_cpu.REG_FILE._04622_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09494_  (.A(\u_cpu.REG_FILE._04622_ ),
    .X(\u_cpu.REG_FILE._00141_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09495_  (.A0(\u_cpu.REG_FILE.rf[3][14] ),
    .A1(\u_cpu.REG_FILE._04457_ ),
    .S(\u_cpu.REG_FILE._04618_ ),
    .X(\u_cpu.REG_FILE._04623_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09496_  (.A(\u_cpu.REG_FILE._04623_ ),
    .X(\u_cpu.REG_FILE._00142_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09497_  (.A0(\u_cpu.REG_FILE.rf[3][15] ),
    .A1(\u_cpu.REG_FILE._04459_ ),
    .S(\u_cpu.REG_FILE._04618_ ),
    .X(\u_cpu.REG_FILE._04624_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09498_  (.A(\u_cpu.REG_FILE._04624_ ),
    .X(\u_cpu.REG_FILE._00143_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09499_  (.A0(\u_cpu.REG_FILE.rf[3][16] ),
    .A1(\u_cpu.REG_FILE._04461_ ),
    .S(\u_cpu.REG_FILE._04618_ ),
    .X(\u_cpu.REG_FILE._04625_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09500_  (.A(\u_cpu.REG_FILE._04625_ ),
    .X(\u_cpu.REG_FILE._00144_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09501_  (.A0(\u_cpu.REG_FILE.rf[3][17] ),
    .A1(\u_cpu.REG_FILE._04463_ ),
    .S(\u_cpu.REG_FILE._04618_ ),
    .X(\u_cpu.REG_FILE._04626_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09502_  (.A(\u_cpu.REG_FILE._04626_ ),
    .X(\u_cpu.REG_FILE._00145_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09503_  (.A0(\u_cpu.REG_FILE.rf[3][18] ),
    .A1(\u_cpu.REG_FILE._04465_ ),
    .S(\u_cpu.REG_FILE._04618_ ),
    .X(\u_cpu.REG_FILE._04627_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09504_  (.A(\u_cpu.REG_FILE._04627_ ),
    .X(\u_cpu.REG_FILE._00146_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09505_  (.A0(\u_cpu.REG_FILE.rf[3][19] ),
    .A1(\u_cpu.REG_FILE._04467_ ),
    .S(\u_cpu.REG_FILE._04618_ ),
    .X(\u_cpu.REG_FILE._04628_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09506_  (.A(\u_cpu.REG_FILE._04628_ ),
    .X(\u_cpu.REG_FILE._00147_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09507_  (.A(\u_cpu.REG_FILE._04606_ ),
    .X(\u_cpu.REG_FILE._04629_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09508_  (.A0(\u_cpu.REG_FILE.rf[3][20] ),
    .A1(\u_cpu.REG_FILE._04469_ ),
    .S(\u_cpu.REG_FILE._04629_ ),
    .X(\u_cpu.REG_FILE._04630_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09509_  (.A(\u_cpu.REG_FILE._04630_ ),
    .X(\u_cpu.REG_FILE._00148_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09510_  (.A0(\u_cpu.REG_FILE.rf[3][21] ),
    .A1(\u_cpu.REG_FILE._04472_ ),
    .S(\u_cpu.REG_FILE._04629_ ),
    .X(\u_cpu.REG_FILE._04631_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09511_  (.A(\u_cpu.REG_FILE._04631_ ),
    .X(\u_cpu.REG_FILE._00149_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09512_  (.A0(\u_cpu.REG_FILE.rf[3][22] ),
    .A1(\u_cpu.REG_FILE._04474_ ),
    .S(\u_cpu.REG_FILE._04629_ ),
    .X(\u_cpu.REG_FILE._04632_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09513_  (.A(\u_cpu.REG_FILE._04632_ ),
    .X(\u_cpu.REG_FILE._00150_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09514_  (.A0(\u_cpu.REG_FILE.rf[3][23] ),
    .A1(\u_cpu.REG_FILE._04476_ ),
    .S(\u_cpu.REG_FILE._04629_ ),
    .X(\u_cpu.REG_FILE._04633_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09515_  (.A(\u_cpu.REG_FILE._04633_ ),
    .X(\u_cpu.REG_FILE._00151_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09516_  (.A0(\u_cpu.REG_FILE.rf[3][24] ),
    .A1(\u_cpu.REG_FILE._04478_ ),
    .S(\u_cpu.REG_FILE._04629_ ),
    .X(\u_cpu.REG_FILE._04634_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09517_  (.A(\u_cpu.REG_FILE._04634_ ),
    .X(\u_cpu.REG_FILE._00152_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09518_  (.A0(\u_cpu.REG_FILE.rf[3][25] ),
    .A1(\u_cpu.REG_FILE._04480_ ),
    .S(\u_cpu.REG_FILE._04629_ ),
    .X(\u_cpu.REG_FILE._04635_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09519_  (.A(\u_cpu.REG_FILE._04635_ ),
    .X(\u_cpu.REG_FILE._00153_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09520_  (.A0(\u_cpu.REG_FILE.rf[3][26] ),
    .A1(\u_cpu.REG_FILE._04482_ ),
    .S(\u_cpu.REG_FILE._04629_ ),
    .X(\u_cpu.REG_FILE._04636_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09521_  (.A(\u_cpu.REG_FILE._04636_ ),
    .X(\u_cpu.REG_FILE._00154_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09522_  (.A0(\u_cpu.REG_FILE.rf[3][27] ),
    .A1(\u_cpu.REG_FILE._04484_ ),
    .S(\u_cpu.REG_FILE._04629_ ),
    .X(\u_cpu.REG_FILE._04637_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09523_  (.A(\u_cpu.REG_FILE._04637_ ),
    .X(\u_cpu.REG_FILE._00155_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09524_  (.A0(\u_cpu.REG_FILE.rf[3][28] ),
    .A1(\u_cpu.REG_FILE._04486_ ),
    .S(\u_cpu.REG_FILE._04629_ ),
    .X(\u_cpu.REG_FILE._04638_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09525_  (.A(\u_cpu.REG_FILE._04638_ ),
    .X(\u_cpu.REG_FILE._00156_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09526_  (.A0(\u_cpu.REG_FILE.rf[3][29] ),
    .A1(\u_cpu.REG_FILE._04488_ ),
    .S(\u_cpu.REG_FILE._04629_ ),
    .X(\u_cpu.REG_FILE._04639_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09527_  (.A(\u_cpu.REG_FILE._04639_ ),
    .X(\u_cpu.REG_FILE._00157_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09528_  (.A0(\u_cpu.REG_FILE.rf[3][30] ),
    .A1(\u_cpu.REG_FILE._04490_ ),
    .S(\u_cpu.REG_FILE._04606_ ),
    .X(\u_cpu.REG_FILE._04640_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09529_  (.A(\u_cpu.REG_FILE._04640_ ),
    .X(\u_cpu.REG_FILE._00158_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09530_  (.A0(\u_cpu.REG_FILE.rf[3][31] ),
    .A1(\u_cpu.REG_FILE._04492_ ),
    .S(\u_cpu.REG_FILE._04606_ ),
    .X(\u_cpu.REG_FILE._04641_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09531_  (.A(\u_cpu.REG_FILE._04641_ ),
    .X(\u_cpu.REG_FILE._00159_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09532_  (.A(\u_cpu.REG_FILE.wd3[0] ),
    .X(\u_cpu.REG_FILE._04642_ ));
 sky130_fd_sc_hd__nor3b_2 \u_cpu.REG_FILE._09533_  (.A(\u_cpu.REG_FILE.a3[1] ),
    .B(\u_cpu.REG_FILE.a3[0] ),
    .C_N(\u_cpu.REG_FILE.we3 ),
    .Y(\u_cpu.REG_FILE._04643_ ));
 sky130_fd_sc_hd__and4bb_2 \u_cpu.REG_FILE._09534_  (.A_N(\u_cpu.REG_FILE._04424_ ),
    .B_N(\u_cpu.REG_FILE._04421_ ),
    .C(\u_cpu.REG_FILE._04494_ ),
    .D(\u_cpu.REG_FILE._04643_ ),
    .X(\u_cpu.REG_FILE._04644_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09535_  (.A(\u_cpu.REG_FILE._04644_ ),
    .X(\u_cpu.REG_FILE._04645_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09536_  (.A0(\u_cpu.REG_FILE.rf[4][0] ),
    .A1(\u_cpu.REG_FILE._04642_ ),
    .S(\u_cpu.REG_FILE._04645_ ),
    .X(\u_cpu.REG_FILE._04646_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09537_  (.A(\u_cpu.REG_FILE._04646_ ),
    .X(\u_cpu.REG_FILE._00160_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09538_  (.A(\u_cpu.REG_FILE.wd3[1] ),
    .X(\u_cpu.REG_FILE._04647_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09539_  (.A0(\u_cpu.REG_FILE.rf[4][1] ),
    .A1(\u_cpu.REG_FILE._04647_ ),
    .S(\u_cpu.REG_FILE._04645_ ),
    .X(\u_cpu.REG_FILE._04648_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09540_  (.A(\u_cpu.REG_FILE._04648_ ),
    .X(\u_cpu.REG_FILE._00161_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09541_  (.A(\u_cpu.REG_FILE.wd3[2] ),
    .X(\u_cpu.REG_FILE._04649_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09542_  (.A0(\u_cpu.REG_FILE.rf[4][2] ),
    .A1(\u_cpu.REG_FILE._04649_ ),
    .S(\u_cpu.REG_FILE._04645_ ),
    .X(\u_cpu.REG_FILE._04650_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09543_  (.A(\u_cpu.REG_FILE._04650_ ),
    .X(\u_cpu.REG_FILE._00162_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09544_  (.A(\u_cpu.REG_FILE.wd3[3] ),
    .X(\u_cpu.REG_FILE._04651_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09545_  (.A0(\u_cpu.REG_FILE.rf[4][3] ),
    .A1(\u_cpu.REG_FILE._04651_ ),
    .S(\u_cpu.REG_FILE._04645_ ),
    .X(\u_cpu.REG_FILE._04652_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09546_  (.A(\u_cpu.REG_FILE._04652_ ),
    .X(\u_cpu.REG_FILE._00163_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09547_  (.A(\u_cpu.REG_FILE.wd3[4] ),
    .X(\u_cpu.REG_FILE._04653_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09548_  (.A0(\u_cpu.REG_FILE.rf[4][4] ),
    .A1(\u_cpu.REG_FILE._04653_ ),
    .S(\u_cpu.REG_FILE._04645_ ),
    .X(\u_cpu.REG_FILE._04654_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09549_  (.A(\u_cpu.REG_FILE._04654_ ),
    .X(\u_cpu.REG_FILE._00164_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09550_  (.A(\u_cpu.REG_FILE.wd3[5] ),
    .X(\u_cpu.REG_FILE._04655_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09551_  (.A0(\u_cpu.REG_FILE.rf[4][5] ),
    .A1(\u_cpu.REG_FILE._04655_ ),
    .S(\u_cpu.REG_FILE._04645_ ),
    .X(\u_cpu.REG_FILE._04656_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09552_  (.A(\u_cpu.REG_FILE._04656_ ),
    .X(\u_cpu.REG_FILE._00165_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09553_  (.A(\u_cpu.REG_FILE.wd3[6] ),
    .X(\u_cpu.REG_FILE._04657_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09554_  (.A0(\u_cpu.REG_FILE.rf[4][6] ),
    .A1(\u_cpu.REG_FILE._04657_ ),
    .S(\u_cpu.REG_FILE._04645_ ),
    .X(\u_cpu.REG_FILE._04658_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09555_  (.A(\u_cpu.REG_FILE._04658_ ),
    .X(\u_cpu.REG_FILE._00166_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09556_  (.A(\u_cpu.REG_FILE.wd3[7] ),
    .X(\u_cpu.REG_FILE._04659_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09557_  (.A0(\u_cpu.REG_FILE.rf[4][7] ),
    .A1(\u_cpu.REG_FILE._04659_ ),
    .S(\u_cpu.REG_FILE._04645_ ),
    .X(\u_cpu.REG_FILE._04660_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09558_  (.A(\u_cpu.REG_FILE._04660_ ),
    .X(\u_cpu.REG_FILE._00167_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09559_  (.A(\u_cpu.REG_FILE.wd3[8] ),
    .X(\u_cpu.REG_FILE._04661_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09560_  (.A0(\u_cpu.REG_FILE.rf[4][8] ),
    .A1(\u_cpu.REG_FILE._04661_ ),
    .S(\u_cpu.REG_FILE._04645_ ),
    .X(\u_cpu.REG_FILE._04662_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09561_  (.A(\u_cpu.REG_FILE._04662_ ),
    .X(\u_cpu.REG_FILE._00168_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09562_  (.A(\u_cpu.REG_FILE.wd3[9] ),
    .X(\u_cpu.REG_FILE._04663_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09563_  (.A0(\u_cpu.REG_FILE.rf[4][9] ),
    .A1(\u_cpu.REG_FILE._04663_ ),
    .S(\u_cpu.REG_FILE._04645_ ),
    .X(\u_cpu.REG_FILE._04664_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09564_  (.A(\u_cpu.REG_FILE._04664_ ),
    .X(\u_cpu.REG_FILE._00169_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09565_  (.A(\u_cpu.REG_FILE.wd3[10] ),
    .X(\u_cpu.REG_FILE._04665_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09566_  (.A(\u_cpu.REG_FILE._04644_ ),
    .X(\u_cpu.REG_FILE._04666_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09567_  (.A0(\u_cpu.REG_FILE.rf[4][10] ),
    .A1(\u_cpu.REG_FILE._04665_ ),
    .S(\u_cpu.REG_FILE._04666_ ),
    .X(\u_cpu.REG_FILE._04667_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09568_  (.A(\u_cpu.REG_FILE._04667_ ),
    .X(\u_cpu.REG_FILE._00170_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09569_  (.A(\u_cpu.REG_FILE.wd3[11] ),
    .X(\u_cpu.REG_FILE._04668_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09570_  (.A0(\u_cpu.REG_FILE.rf[4][11] ),
    .A1(\u_cpu.REG_FILE._04668_ ),
    .S(\u_cpu.REG_FILE._04666_ ),
    .X(\u_cpu.REG_FILE._04669_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09571_  (.A(\u_cpu.REG_FILE._04669_ ),
    .X(\u_cpu.REG_FILE._00171_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09572_  (.A(\u_cpu.REG_FILE.wd3[12] ),
    .X(\u_cpu.REG_FILE._04670_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09573_  (.A0(\u_cpu.REG_FILE.rf[4][12] ),
    .A1(\u_cpu.REG_FILE._04670_ ),
    .S(\u_cpu.REG_FILE._04666_ ),
    .X(\u_cpu.REG_FILE._04671_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09574_  (.A(\u_cpu.REG_FILE._04671_ ),
    .X(\u_cpu.REG_FILE._00172_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09575_  (.A(\u_cpu.REG_FILE.wd3[13] ),
    .X(\u_cpu.REG_FILE._04672_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09576_  (.A0(\u_cpu.REG_FILE.rf[4][13] ),
    .A1(\u_cpu.REG_FILE._04672_ ),
    .S(\u_cpu.REG_FILE._04666_ ),
    .X(\u_cpu.REG_FILE._04673_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09577_  (.A(\u_cpu.REG_FILE._04673_ ),
    .X(\u_cpu.REG_FILE._00173_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09578_  (.A(\u_cpu.REG_FILE.wd3[14] ),
    .X(\u_cpu.REG_FILE._04674_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09579_  (.A0(\u_cpu.REG_FILE.rf[4][14] ),
    .A1(\u_cpu.REG_FILE._04674_ ),
    .S(\u_cpu.REG_FILE._04666_ ),
    .X(\u_cpu.REG_FILE._04675_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09580_  (.A(\u_cpu.REG_FILE._04675_ ),
    .X(\u_cpu.REG_FILE._00174_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09581_  (.A(\u_cpu.REG_FILE.wd3[15] ),
    .X(\u_cpu.REG_FILE._04676_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09582_  (.A0(\u_cpu.REG_FILE.rf[4][15] ),
    .A1(\u_cpu.REG_FILE._04676_ ),
    .S(\u_cpu.REG_FILE._04666_ ),
    .X(\u_cpu.REG_FILE._04677_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09583_  (.A(\u_cpu.REG_FILE._04677_ ),
    .X(\u_cpu.REG_FILE._00175_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09584_  (.A(\u_cpu.REG_FILE.wd3[16] ),
    .X(\u_cpu.REG_FILE._04678_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09585_  (.A0(\u_cpu.REG_FILE.rf[4][16] ),
    .A1(\u_cpu.REG_FILE._04678_ ),
    .S(\u_cpu.REG_FILE._04666_ ),
    .X(\u_cpu.REG_FILE._04679_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09586_  (.A(\u_cpu.REG_FILE._04679_ ),
    .X(\u_cpu.REG_FILE._00176_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09587_  (.A(\u_cpu.REG_FILE.wd3[17] ),
    .X(\u_cpu.REG_FILE._04680_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09588_  (.A0(\u_cpu.REG_FILE.rf[4][17] ),
    .A1(\u_cpu.REG_FILE._04680_ ),
    .S(\u_cpu.REG_FILE._04666_ ),
    .X(\u_cpu.REG_FILE._04681_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09589_  (.A(\u_cpu.REG_FILE._04681_ ),
    .X(\u_cpu.REG_FILE._00177_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09590_  (.A(\u_cpu.REG_FILE.wd3[18] ),
    .X(\u_cpu.REG_FILE._04682_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09591_  (.A0(\u_cpu.REG_FILE.rf[4][18] ),
    .A1(\u_cpu.REG_FILE._04682_ ),
    .S(\u_cpu.REG_FILE._04666_ ),
    .X(\u_cpu.REG_FILE._04683_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09592_  (.A(\u_cpu.REG_FILE._04683_ ),
    .X(\u_cpu.REG_FILE._00178_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09593_  (.A(\u_cpu.REG_FILE.wd3[19] ),
    .X(\u_cpu.REG_FILE._04684_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09594_  (.A0(\u_cpu.REG_FILE.rf[4][19] ),
    .A1(\u_cpu.REG_FILE._04684_ ),
    .S(\u_cpu.REG_FILE._04666_ ),
    .X(\u_cpu.REG_FILE._04685_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09595_  (.A(\u_cpu.REG_FILE._04685_ ),
    .X(\u_cpu.REG_FILE._00179_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09596_  (.A(\u_cpu.REG_FILE.wd3[20] ),
    .X(\u_cpu.REG_FILE._04686_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09597_  (.A(\u_cpu.REG_FILE._04644_ ),
    .X(\u_cpu.REG_FILE._04687_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09598_  (.A0(\u_cpu.REG_FILE.rf[4][20] ),
    .A1(\u_cpu.REG_FILE._04686_ ),
    .S(\u_cpu.REG_FILE._04687_ ),
    .X(\u_cpu.REG_FILE._04688_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09599_  (.A(\u_cpu.REG_FILE._04688_ ),
    .X(\u_cpu.REG_FILE._00180_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09600_  (.A(\u_cpu.REG_FILE.wd3[21] ),
    .X(\u_cpu.REG_FILE._04689_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09601_  (.A0(\u_cpu.REG_FILE.rf[4][21] ),
    .A1(\u_cpu.REG_FILE._04689_ ),
    .S(\u_cpu.REG_FILE._04687_ ),
    .X(\u_cpu.REG_FILE._04690_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09602_  (.A(\u_cpu.REG_FILE._04690_ ),
    .X(\u_cpu.REG_FILE._00181_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09603_  (.A(\u_cpu.REG_FILE.wd3[22] ),
    .X(\u_cpu.REG_FILE._04691_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09604_  (.A0(\u_cpu.REG_FILE.rf[4][22] ),
    .A1(\u_cpu.REG_FILE._04691_ ),
    .S(\u_cpu.REG_FILE._04687_ ),
    .X(\u_cpu.REG_FILE._04692_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09605_  (.A(\u_cpu.REG_FILE._04692_ ),
    .X(\u_cpu.REG_FILE._00182_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09606_  (.A(\u_cpu.REG_FILE.wd3[23] ),
    .X(\u_cpu.REG_FILE._04693_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09607_  (.A0(\u_cpu.REG_FILE.rf[4][23] ),
    .A1(\u_cpu.REG_FILE._04693_ ),
    .S(\u_cpu.REG_FILE._04687_ ),
    .X(\u_cpu.REG_FILE._04694_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09608_  (.A(\u_cpu.REG_FILE._04694_ ),
    .X(\u_cpu.REG_FILE._00183_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09609_  (.A(\u_cpu.REG_FILE.wd3[24] ),
    .X(\u_cpu.REG_FILE._04695_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09610_  (.A0(\u_cpu.REG_FILE.rf[4][24] ),
    .A1(\u_cpu.REG_FILE._04695_ ),
    .S(\u_cpu.REG_FILE._04687_ ),
    .X(\u_cpu.REG_FILE._04696_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09611_  (.A(\u_cpu.REG_FILE._04696_ ),
    .X(\u_cpu.REG_FILE._00184_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09612_  (.A(\u_cpu.REG_FILE.wd3[25] ),
    .X(\u_cpu.REG_FILE._04697_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09613_  (.A0(\u_cpu.REG_FILE.rf[4][25] ),
    .A1(\u_cpu.REG_FILE._04697_ ),
    .S(\u_cpu.REG_FILE._04687_ ),
    .X(\u_cpu.REG_FILE._04698_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09614_  (.A(\u_cpu.REG_FILE._04698_ ),
    .X(\u_cpu.REG_FILE._00185_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09615_  (.A(\u_cpu.REG_FILE.wd3[26] ),
    .X(\u_cpu.REG_FILE._04699_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09616_  (.A0(\u_cpu.REG_FILE.rf[4][26] ),
    .A1(\u_cpu.REG_FILE._04699_ ),
    .S(\u_cpu.REG_FILE._04687_ ),
    .X(\u_cpu.REG_FILE._04700_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09617_  (.A(\u_cpu.REG_FILE._04700_ ),
    .X(\u_cpu.REG_FILE._00186_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09618_  (.A(\u_cpu.REG_FILE.wd3[27] ),
    .X(\u_cpu.REG_FILE._04701_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09619_  (.A0(\u_cpu.REG_FILE.rf[4][27] ),
    .A1(\u_cpu.REG_FILE._04701_ ),
    .S(\u_cpu.REG_FILE._04687_ ),
    .X(\u_cpu.REG_FILE._04702_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09620_  (.A(\u_cpu.REG_FILE._04702_ ),
    .X(\u_cpu.REG_FILE._00187_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09621_  (.A(\u_cpu.REG_FILE.wd3[28] ),
    .X(\u_cpu.REG_FILE._04703_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09622_  (.A0(\u_cpu.REG_FILE.rf[4][28] ),
    .A1(\u_cpu.REG_FILE._04703_ ),
    .S(\u_cpu.REG_FILE._04687_ ),
    .X(\u_cpu.REG_FILE._04704_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09623_  (.A(\u_cpu.REG_FILE._04704_ ),
    .X(\u_cpu.REG_FILE._00188_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09624_  (.A(\u_cpu.REG_FILE.wd3[29] ),
    .X(\u_cpu.REG_FILE._04705_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09625_  (.A0(\u_cpu.REG_FILE.rf[4][29] ),
    .A1(\u_cpu.REG_FILE._04705_ ),
    .S(\u_cpu.REG_FILE._04687_ ),
    .X(\u_cpu.REG_FILE._04706_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09626_  (.A(\u_cpu.REG_FILE._04706_ ),
    .X(\u_cpu.REG_FILE._00189_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09627_  (.A(\u_cpu.REG_FILE.wd3[30] ),
    .X(\u_cpu.REG_FILE._04707_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09628_  (.A0(\u_cpu.REG_FILE.rf[4][30] ),
    .A1(\u_cpu.REG_FILE._04707_ ),
    .S(\u_cpu.REG_FILE._04644_ ),
    .X(\u_cpu.REG_FILE._04708_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09629_  (.A(\u_cpu.REG_FILE._04708_ ),
    .X(\u_cpu.REG_FILE._00190_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09630_  (.A(\u_cpu.REG_FILE.wd3[31] ),
    .X(\u_cpu.REG_FILE._04709_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09631_  (.A0(\u_cpu.REG_FILE.rf[4][31] ),
    .A1(\u_cpu.REG_FILE._04709_ ),
    .S(\u_cpu.REG_FILE._04644_ ),
    .X(\u_cpu.REG_FILE._04710_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09632_  (.A(\u_cpu.REG_FILE._04710_ ),
    .X(\u_cpu.REG_FILE._00191_ ));
 sky130_fd_sc_hd__or4bb_2 \u_cpu.REG_FILE._09633_  (.A(\u_cpu.REG_FILE._04496_ ),
    .B(\u_cpu.REG_FILE._04421_ ),
    .C_N(\u_cpu.REG_FILE._04494_ ),
    .D_N(\u_cpu.REG_FILE._04423_ ),
    .X(\u_cpu.REG_FILE._04711_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09634_  (.A(\u_cpu.REG_FILE._04711_ ),
    .X(\u_cpu.REG_FILE._04712_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09635_  (.A0(\u_cpu.REG_FILE._04420_ ),
    .A1(\u_cpu.REG_FILE.rf[5][0] ),
    .S(\u_cpu.REG_FILE._04712_ ),
    .X(\u_cpu.REG_FILE._04713_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09636_  (.A(\u_cpu.REG_FILE._04713_ ),
    .X(\u_cpu.REG_FILE._00192_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09637_  (.A0(\u_cpu.REG_FILE._04430_ ),
    .A1(\u_cpu.REG_FILE.rf[5][1] ),
    .S(\u_cpu.REG_FILE._04712_ ),
    .X(\u_cpu.REG_FILE._04714_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09638_  (.A(\u_cpu.REG_FILE._04714_ ),
    .X(\u_cpu.REG_FILE._00193_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09639_  (.A0(\u_cpu.REG_FILE._04432_ ),
    .A1(\u_cpu.REG_FILE.rf[5][2] ),
    .S(\u_cpu.REG_FILE._04712_ ),
    .X(\u_cpu.REG_FILE._04715_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09640_  (.A(\u_cpu.REG_FILE._04715_ ),
    .X(\u_cpu.REG_FILE._00194_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09641_  (.A0(\u_cpu.REG_FILE._04434_ ),
    .A1(\u_cpu.REG_FILE.rf[5][3] ),
    .S(\u_cpu.REG_FILE._04712_ ),
    .X(\u_cpu.REG_FILE._04716_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09642_  (.A(\u_cpu.REG_FILE._04716_ ),
    .X(\u_cpu.REG_FILE._00195_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09643_  (.A0(\u_cpu.REG_FILE._04436_ ),
    .A1(\u_cpu.REG_FILE.rf[5][4] ),
    .S(\u_cpu.REG_FILE._04712_ ),
    .X(\u_cpu.REG_FILE._04717_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09644_  (.A(\u_cpu.REG_FILE._04717_ ),
    .X(\u_cpu.REG_FILE._00196_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09645_  (.A0(\u_cpu.REG_FILE._04438_ ),
    .A1(\u_cpu.REG_FILE.rf[5][5] ),
    .S(\u_cpu.REG_FILE._04712_ ),
    .X(\u_cpu.REG_FILE._04718_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09646_  (.A(\u_cpu.REG_FILE._04718_ ),
    .X(\u_cpu.REG_FILE._00197_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09647_  (.A0(\u_cpu.REG_FILE._04440_ ),
    .A1(\u_cpu.REG_FILE.rf[5][6] ),
    .S(\u_cpu.REG_FILE._04712_ ),
    .X(\u_cpu.REG_FILE._04719_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09648_  (.A(\u_cpu.REG_FILE._04719_ ),
    .X(\u_cpu.REG_FILE._00198_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09649_  (.A0(\u_cpu.REG_FILE._04442_ ),
    .A1(\u_cpu.REG_FILE.rf[5][7] ),
    .S(\u_cpu.REG_FILE._04712_ ),
    .X(\u_cpu.REG_FILE._04720_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09650_  (.A(\u_cpu.REG_FILE._04720_ ),
    .X(\u_cpu.REG_FILE._00199_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09651_  (.A0(\u_cpu.REG_FILE._04444_ ),
    .A1(\u_cpu.REG_FILE.rf[5][8] ),
    .S(\u_cpu.REG_FILE._04712_ ),
    .X(\u_cpu.REG_FILE._04721_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09652_  (.A(\u_cpu.REG_FILE._04721_ ),
    .X(\u_cpu.REG_FILE._00200_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09653_  (.A0(\u_cpu.REG_FILE._04446_ ),
    .A1(\u_cpu.REG_FILE.rf[5][9] ),
    .S(\u_cpu.REG_FILE._04712_ ),
    .X(\u_cpu.REG_FILE._04722_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09654_  (.A(\u_cpu.REG_FILE._04722_ ),
    .X(\u_cpu.REG_FILE._00201_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09655_  (.A(\u_cpu.REG_FILE._04711_ ),
    .X(\u_cpu.REG_FILE._04723_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09656_  (.A0(\u_cpu.REG_FILE._04448_ ),
    .A1(\u_cpu.REG_FILE.rf[5][10] ),
    .S(\u_cpu.REG_FILE._04723_ ),
    .X(\u_cpu.REG_FILE._04724_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09657_  (.A(\u_cpu.REG_FILE._04724_ ),
    .X(\u_cpu.REG_FILE._00202_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09658_  (.A0(\u_cpu.REG_FILE._04451_ ),
    .A1(\u_cpu.REG_FILE.rf[5][11] ),
    .S(\u_cpu.REG_FILE._04723_ ),
    .X(\u_cpu.REG_FILE._04725_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09659_  (.A(\u_cpu.REG_FILE._04725_ ),
    .X(\u_cpu.REG_FILE._00203_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09660_  (.A0(\u_cpu.REG_FILE._04453_ ),
    .A1(\u_cpu.REG_FILE.rf[5][12] ),
    .S(\u_cpu.REG_FILE._04723_ ),
    .X(\u_cpu.REG_FILE._04726_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09661_  (.A(\u_cpu.REG_FILE._04726_ ),
    .X(\u_cpu.REG_FILE._00204_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09662_  (.A0(\u_cpu.REG_FILE._04455_ ),
    .A1(\u_cpu.REG_FILE.rf[5][13] ),
    .S(\u_cpu.REG_FILE._04723_ ),
    .X(\u_cpu.REG_FILE._04727_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09663_  (.A(\u_cpu.REG_FILE._04727_ ),
    .X(\u_cpu.REG_FILE._00205_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09664_  (.A0(\u_cpu.REG_FILE._04457_ ),
    .A1(\u_cpu.REG_FILE.rf[5][14] ),
    .S(\u_cpu.REG_FILE._04723_ ),
    .X(\u_cpu.REG_FILE._04728_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09665_  (.A(\u_cpu.REG_FILE._04728_ ),
    .X(\u_cpu.REG_FILE._00206_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09666_  (.A0(\u_cpu.REG_FILE._04459_ ),
    .A1(\u_cpu.REG_FILE.rf[5][15] ),
    .S(\u_cpu.REG_FILE._04723_ ),
    .X(\u_cpu.REG_FILE._04729_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09667_  (.A(\u_cpu.REG_FILE._04729_ ),
    .X(\u_cpu.REG_FILE._00207_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09668_  (.A0(\u_cpu.REG_FILE._04461_ ),
    .A1(\u_cpu.REG_FILE.rf[5][16] ),
    .S(\u_cpu.REG_FILE._04723_ ),
    .X(\u_cpu.REG_FILE._04730_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09669_  (.A(\u_cpu.REG_FILE._04730_ ),
    .X(\u_cpu.REG_FILE._00208_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09670_  (.A0(\u_cpu.REG_FILE._04463_ ),
    .A1(\u_cpu.REG_FILE.rf[5][17] ),
    .S(\u_cpu.REG_FILE._04723_ ),
    .X(\u_cpu.REG_FILE._04731_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09671_  (.A(\u_cpu.REG_FILE._04731_ ),
    .X(\u_cpu.REG_FILE._00209_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09672_  (.A0(\u_cpu.REG_FILE._04465_ ),
    .A1(\u_cpu.REG_FILE.rf[5][18] ),
    .S(\u_cpu.REG_FILE._04723_ ),
    .X(\u_cpu.REG_FILE._04732_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09673_  (.A(\u_cpu.REG_FILE._04732_ ),
    .X(\u_cpu.REG_FILE._00210_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09674_  (.A0(\u_cpu.REG_FILE._04467_ ),
    .A1(\u_cpu.REG_FILE.rf[5][19] ),
    .S(\u_cpu.REG_FILE._04723_ ),
    .X(\u_cpu.REG_FILE._04733_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09675_  (.A(\u_cpu.REG_FILE._04733_ ),
    .X(\u_cpu.REG_FILE._00211_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09676_  (.A(\u_cpu.REG_FILE._04711_ ),
    .X(\u_cpu.REG_FILE._04734_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09677_  (.A0(\u_cpu.REG_FILE._04469_ ),
    .A1(\u_cpu.REG_FILE.rf[5][20] ),
    .S(\u_cpu.REG_FILE._04734_ ),
    .X(\u_cpu.REG_FILE._04735_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09678_  (.A(\u_cpu.REG_FILE._04735_ ),
    .X(\u_cpu.REG_FILE._00212_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09679_  (.A0(\u_cpu.REG_FILE._04472_ ),
    .A1(\u_cpu.REG_FILE.rf[5][21] ),
    .S(\u_cpu.REG_FILE._04734_ ),
    .X(\u_cpu.REG_FILE._04736_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09680_  (.A(\u_cpu.REG_FILE._04736_ ),
    .X(\u_cpu.REG_FILE._00213_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09681_  (.A0(\u_cpu.REG_FILE._04474_ ),
    .A1(\u_cpu.REG_FILE.rf[5][22] ),
    .S(\u_cpu.REG_FILE._04734_ ),
    .X(\u_cpu.REG_FILE._04737_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09682_  (.A(\u_cpu.REG_FILE._04737_ ),
    .X(\u_cpu.REG_FILE._00214_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09683_  (.A0(\u_cpu.REG_FILE._04476_ ),
    .A1(\u_cpu.REG_FILE.rf[5][23] ),
    .S(\u_cpu.REG_FILE._04734_ ),
    .X(\u_cpu.REG_FILE._04738_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09684_  (.A(\u_cpu.REG_FILE._04738_ ),
    .X(\u_cpu.REG_FILE._00215_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09685_  (.A0(\u_cpu.REG_FILE._04478_ ),
    .A1(\u_cpu.REG_FILE.rf[5][24] ),
    .S(\u_cpu.REG_FILE._04734_ ),
    .X(\u_cpu.REG_FILE._04739_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09686_  (.A(\u_cpu.REG_FILE._04739_ ),
    .X(\u_cpu.REG_FILE._00216_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09687_  (.A0(\u_cpu.REG_FILE._04480_ ),
    .A1(\u_cpu.REG_FILE.rf[5][25] ),
    .S(\u_cpu.REG_FILE._04734_ ),
    .X(\u_cpu.REG_FILE._04740_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09688_  (.A(\u_cpu.REG_FILE._04740_ ),
    .X(\u_cpu.REG_FILE._00217_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09689_  (.A0(\u_cpu.REG_FILE._04482_ ),
    .A1(\u_cpu.REG_FILE.rf[5][26] ),
    .S(\u_cpu.REG_FILE._04734_ ),
    .X(\u_cpu.REG_FILE._04741_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09690_  (.A(\u_cpu.REG_FILE._04741_ ),
    .X(\u_cpu.REG_FILE._00218_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09691_  (.A0(\u_cpu.REG_FILE._04484_ ),
    .A1(\u_cpu.REG_FILE.rf[5][27] ),
    .S(\u_cpu.REG_FILE._04734_ ),
    .X(\u_cpu.REG_FILE._04742_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09692_  (.A(\u_cpu.REG_FILE._04742_ ),
    .X(\u_cpu.REG_FILE._00219_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09693_  (.A0(\u_cpu.REG_FILE._04486_ ),
    .A1(\u_cpu.REG_FILE.rf[5][28] ),
    .S(\u_cpu.REG_FILE._04734_ ),
    .X(\u_cpu.REG_FILE._04743_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09694_  (.A(\u_cpu.REG_FILE._04743_ ),
    .X(\u_cpu.REG_FILE._00220_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09695_  (.A0(\u_cpu.REG_FILE._04488_ ),
    .A1(\u_cpu.REG_FILE.rf[5][29] ),
    .S(\u_cpu.REG_FILE._04734_ ),
    .X(\u_cpu.REG_FILE._04744_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09696_  (.A(\u_cpu.REG_FILE._04744_ ),
    .X(\u_cpu.REG_FILE._00221_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09697_  (.A0(\u_cpu.REG_FILE._04490_ ),
    .A1(\u_cpu.REG_FILE.rf[5][30] ),
    .S(\u_cpu.REG_FILE._04711_ ),
    .X(\u_cpu.REG_FILE._04745_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09698_  (.A(\u_cpu.REG_FILE._04745_ ),
    .X(\u_cpu.REG_FILE._00222_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09699_  (.A0(\u_cpu.REG_FILE._04492_ ),
    .A1(\u_cpu.REG_FILE.rf[5][31] ),
    .S(\u_cpu.REG_FILE._04711_ ),
    .X(\u_cpu.REG_FILE._04746_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09700_  (.A(\u_cpu.REG_FILE._04746_ ),
    .X(\u_cpu.REG_FILE._00223_ ));
 sky130_fd_sc_hd__and3b_2 \u_cpu.REG_FILE._09701_  (.A_N(\u_cpu.REG_FILE.a3[0] ),
    .B(\u_cpu.REG_FILE.we3 ),
    .C(\u_cpu.REG_FILE.a3[1] ),
    .X(\u_cpu.REG_FILE._04747_ ));
 sky130_fd_sc_hd__and4bb_2 \u_cpu.REG_FILE._09702_  (.A_N(\u_cpu.REG_FILE._04424_ ),
    .B_N(\u_cpu.REG_FILE._04421_ ),
    .C(\u_cpu.REG_FILE._04494_ ),
    .D(\u_cpu.REG_FILE._04747_ ),
    .X(\u_cpu.REG_FILE._04748_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09703_  (.A(\u_cpu.REG_FILE._04748_ ),
    .X(\u_cpu.REG_FILE._04749_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09704_  (.A0(\u_cpu.REG_FILE.rf[6][0] ),
    .A1(\u_cpu.REG_FILE._04642_ ),
    .S(\u_cpu.REG_FILE._04749_ ),
    .X(\u_cpu.REG_FILE._04750_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09705_  (.A(\u_cpu.REG_FILE._04750_ ),
    .X(\u_cpu.REG_FILE._00224_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09706_  (.A0(\u_cpu.REG_FILE.rf[6][1] ),
    .A1(\u_cpu.REG_FILE._04647_ ),
    .S(\u_cpu.REG_FILE._04749_ ),
    .X(\u_cpu.REG_FILE._04751_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09707_  (.A(\u_cpu.REG_FILE._04751_ ),
    .X(\u_cpu.REG_FILE._00225_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09708_  (.A0(\u_cpu.REG_FILE.rf[6][2] ),
    .A1(\u_cpu.REG_FILE._04649_ ),
    .S(\u_cpu.REG_FILE._04749_ ),
    .X(\u_cpu.REG_FILE._04752_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09709_  (.A(\u_cpu.REG_FILE._04752_ ),
    .X(\u_cpu.REG_FILE._00226_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09710_  (.A0(\u_cpu.REG_FILE.rf[6][3] ),
    .A1(\u_cpu.REG_FILE._04651_ ),
    .S(\u_cpu.REG_FILE._04749_ ),
    .X(\u_cpu.REG_FILE._04753_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09711_  (.A(\u_cpu.REG_FILE._04753_ ),
    .X(\u_cpu.REG_FILE._00227_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09712_  (.A0(\u_cpu.REG_FILE.rf[6][4] ),
    .A1(\u_cpu.REG_FILE._04653_ ),
    .S(\u_cpu.REG_FILE._04749_ ),
    .X(\u_cpu.REG_FILE._04754_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09713_  (.A(\u_cpu.REG_FILE._04754_ ),
    .X(\u_cpu.REG_FILE._00228_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09714_  (.A0(\u_cpu.REG_FILE.rf[6][5] ),
    .A1(\u_cpu.REG_FILE._04655_ ),
    .S(\u_cpu.REG_FILE._04749_ ),
    .X(\u_cpu.REG_FILE._04755_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09715_  (.A(\u_cpu.REG_FILE._04755_ ),
    .X(\u_cpu.REG_FILE._00229_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09716_  (.A0(\u_cpu.REG_FILE.rf[6][6] ),
    .A1(\u_cpu.REG_FILE._04657_ ),
    .S(\u_cpu.REG_FILE._04749_ ),
    .X(\u_cpu.REG_FILE._04756_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09717_  (.A(\u_cpu.REG_FILE._04756_ ),
    .X(\u_cpu.REG_FILE._00230_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09718_  (.A0(\u_cpu.REG_FILE.rf[6][7] ),
    .A1(\u_cpu.REG_FILE._04659_ ),
    .S(\u_cpu.REG_FILE._04749_ ),
    .X(\u_cpu.REG_FILE._04757_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09719_  (.A(\u_cpu.REG_FILE._04757_ ),
    .X(\u_cpu.REG_FILE._00231_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09720_  (.A0(\u_cpu.REG_FILE.rf[6][8] ),
    .A1(\u_cpu.REG_FILE._04661_ ),
    .S(\u_cpu.REG_FILE._04749_ ),
    .X(\u_cpu.REG_FILE._04758_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09721_  (.A(\u_cpu.REG_FILE._04758_ ),
    .X(\u_cpu.REG_FILE._00232_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09722_  (.A0(\u_cpu.REG_FILE.rf[6][9] ),
    .A1(\u_cpu.REG_FILE._04663_ ),
    .S(\u_cpu.REG_FILE._04749_ ),
    .X(\u_cpu.REG_FILE._04759_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09723_  (.A(\u_cpu.REG_FILE._04759_ ),
    .X(\u_cpu.REG_FILE._00233_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09724_  (.A(\u_cpu.REG_FILE._04748_ ),
    .X(\u_cpu.REG_FILE._04760_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09725_  (.A0(\u_cpu.REG_FILE.rf[6][10] ),
    .A1(\u_cpu.REG_FILE._04665_ ),
    .S(\u_cpu.REG_FILE._04760_ ),
    .X(\u_cpu.REG_FILE._04761_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09726_  (.A(\u_cpu.REG_FILE._04761_ ),
    .X(\u_cpu.REG_FILE._00234_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09727_  (.A0(\u_cpu.REG_FILE.rf[6][11] ),
    .A1(\u_cpu.REG_FILE._04668_ ),
    .S(\u_cpu.REG_FILE._04760_ ),
    .X(\u_cpu.REG_FILE._04762_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09728_  (.A(\u_cpu.REG_FILE._04762_ ),
    .X(\u_cpu.REG_FILE._00235_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09729_  (.A0(\u_cpu.REG_FILE.rf[6][12] ),
    .A1(\u_cpu.REG_FILE._04670_ ),
    .S(\u_cpu.REG_FILE._04760_ ),
    .X(\u_cpu.REG_FILE._04763_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09730_  (.A(\u_cpu.REG_FILE._04763_ ),
    .X(\u_cpu.REG_FILE._00236_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09731_  (.A0(\u_cpu.REG_FILE.rf[6][13] ),
    .A1(\u_cpu.REG_FILE._04672_ ),
    .S(\u_cpu.REG_FILE._04760_ ),
    .X(\u_cpu.REG_FILE._04764_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09732_  (.A(\u_cpu.REG_FILE._04764_ ),
    .X(\u_cpu.REG_FILE._00237_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09733_  (.A0(\u_cpu.REG_FILE.rf[6][14] ),
    .A1(\u_cpu.REG_FILE._04674_ ),
    .S(\u_cpu.REG_FILE._04760_ ),
    .X(\u_cpu.REG_FILE._04765_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09734_  (.A(\u_cpu.REG_FILE._04765_ ),
    .X(\u_cpu.REG_FILE._00238_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09735_  (.A0(\u_cpu.REG_FILE.rf[6][15] ),
    .A1(\u_cpu.REG_FILE._04676_ ),
    .S(\u_cpu.REG_FILE._04760_ ),
    .X(\u_cpu.REG_FILE._04766_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09736_  (.A(\u_cpu.REG_FILE._04766_ ),
    .X(\u_cpu.REG_FILE._00239_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09737_  (.A0(\u_cpu.REG_FILE.rf[6][16] ),
    .A1(\u_cpu.REG_FILE._04678_ ),
    .S(\u_cpu.REG_FILE._04760_ ),
    .X(\u_cpu.REG_FILE._04767_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09738_  (.A(\u_cpu.REG_FILE._04767_ ),
    .X(\u_cpu.REG_FILE._00240_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09739_  (.A0(\u_cpu.REG_FILE.rf[6][17] ),
    .A1(\u_cpu.REG_FILE._04680_ ),
    .S(\u_cpu.REG_FILE._04760_ ),
    .X(\u_cpu.REG_FILE._04768_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09740_  (.A(\u_cpu.REG_FILE._04768_ ),
    .X(\u_cpu.REG_FILE._00241_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09741_  (.A0(\u_cpu.REG_FILE.rf[6][18] ),
    .A1(\u_cpu.REG_FILE._04682_ ),
    .S(\u_cpu.REG_FILE._04760_ ),
    .X(\u_cpu.REG_FILE._04769_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09742_  (.A(\u_cpu.REG_FILE._04769_ ),
    .X(\u_cpu.REG_FILE._00242_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09743_  (.A0(\u_cpu.REG_FILE.rf[6][19] ),
    .A1(\u_cpu.REG_FILE._04684_ ),
    .S(\u_cpu.REG_FILE._04760_ ),
    .X(\u_cpu.REG_FILE._04770_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09744_  (.A(\u_cpu.REG_FILE._04770_ ),
    .X(\u_cpu.REG_FILE._00243_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09745_  (.A(\u_cpu.REG_FILE._04748_ ),
    .X(\u_cpu.REG_FILE._04771_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09746_  (.A0(\u_cpu.REG_FILE.rf[6][20] ),
    .A1(\u_cpu.REG_FILE._04686_ ),
    .S(\u_cpu.REG_FILE._04771_ ),
    .X(\u_cpu.REG_FILE._04772_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09747_  (.A(\u_cpu.REG_FILE._04772_ ),
    .X(\u_cpu.REG_FILE._00244_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09748_  (.A0(\u_cpu.REG_FILE.rf[6][21] ),
    .A1(\u_cpu.REG_FILE._04689_ ),
    .S(\u_cpu.REG_FILE._04771_ ),
    .X(\u_cpu.REG_FILE._04773_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09749_  (.A(\u_cpu.REG_FILE._04773_ ),
    .X(\u_cpu.REG_FILE._00245_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09750_  (.A0(\u_cpu.REG_FILE.rf[6][22] ),
    .A1(\u_cpu.REG_FILE._04691_ ),
    .S(\u_cpu.REG_FILE._04771_ ),
    .X(\u_cpu.REG_FILE._04774_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09751_  (.A(\u_cpu.REG_FILE._04774_ ),
    .X(\u_cpu.REG_FILE._00246_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09752_  (.A0(\u_cpu.REG_FILE.rf[6][23] ),
    .A1(\u_cpu.REG_FILE._04693_ ),
    .S(\u_cpu.REG_FILE._04771_ ),
    .X(\u_cpu.REG_FILE._04775_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09753_  (.A(\u_cpu.REG_FILE._04775_ ),
    .X(\u_cpu.REG_FILE._00247_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09754_  (.A0(\u_cpu.REG_FILE.rf[6][24] ),
    .A1(\u_cpu.REG_FILE._04695_ ),
    .S(\u_cpu.REG_FILE._04771_ ),
    .X(\u_cpu.REG_FILE._04776_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09755_  (.A(\u_cpu.REG_FILE._04776_ ),
    .X(\u_cpu.REG_FILE._00248_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09756_  (.A0(\u_cpu.REG_FILE.rf[6][25] ),
    .A1(\u_cpu.REG_FILE._04697_ ),
    .S(\u_cpu.REG_FILE._04771_ ),
    .X(\u_cpu.REG_FILE._04777_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09757_  (.A(\u_cpu.REG_FILE._04777_ ),
    .X(\u_cpu.REG_FILE._00249_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09758_  (.A0(\u_cpu.REG_FILE.rf[6][26] ),
    .A1(\u_cpu.REG_FILE._04699_ ),
    .S(\u_cpu.REG_FILE._04771_ ),
    .X(\u_cpu.REG_FILE._04778_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09759_  (.A(\u_cpu.REG_FILE._04778_ ),
    .X(\u_cpu.REG_FILE._00250_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09760_  (.A0(\u_cpu.REG_FILE.rf[6][27] ),
    .A1(\u_cpu.REG_FILE._04701_ ),
    .S(\u_cpu.REG_FILE._04771_ ),
    .X(\u_cpu.REG_FILE._04779_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09761_  (.A(\u_cpu.REG_FILE._04779_ ),
    .X(\u_cpu.REG_FILE._00251_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09762_  (.A0(\u_cpu.REG_FILE.rf[6][28] ),
    .A1(\u_cpu.REG_FILE._04703_ ),
    .S(\u_cpu.REG_FILE._04771_ ),
    .X(\u_cpu.REG_FILE._04780_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09763_  (.A(\u_cpu.REG_FILE._04780_ ),
    .X(\u_cpu.REG_FILE._00252_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09764_  (.A0(\u_cpu.REG_FILE.rf[6][29] ),
    .A1(\u_cpu.REG_FILE._04705_ ),
    .S(\u_cpu.REG_FILE._04771_ ),
    .X(\u_cpu.REG_FILE._04781_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09765_  (.A(\u_cpu.REG_FILE._04781_ ),
    .X(\u_cpu.REG_FILE._00253_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09766_  (.A0(\u_cpu.REG_FILE.rf[6][30] ),
    .A1(\u_cpu.REG_FILE._04707_ ),
    .S(\u_cpu.REG_FILE._04748_ ),
    .X(\u_cpu.REG_FILE._04782_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09767_  (.A(\u_cpu.REG_FILE._04782_ ),
    .X(\u_cpu.REG_FILE._00254_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09768_  (.A0(\u_cpu.REG_FILE.rf[6][31] ),
    .A1(\u_cpu.REG_FILE._04709_ ),
    .S(\u_cpu.REG_FILE._04748_ ),
    .X(\u_cpu.REG_FILE._04783_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09769_  (.A(\u_cpu.REG_FILE._04783_ ),
    .X(\u_cpu.REG_FILE._00255_ ));
 sky130_fd_sc_hd__and4bb_2 \u_cpu.REG_FILE._09770_  (.A_N(\u_cpu.REG_FILE._04424_ ),
    .B_N(\u_cpu.REG_FILE._04421_ ),
    .C(\u_cpu.REG_FILE._04425_ ),
    .D(\u_cpu.REG_FILE._04495_ ),
    .X(\u_cpu.REG_FILE._04784_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09771_  (.A(\u_cpu.REG_FILE._04784_ ),
    .X(\u_cpu.REG_FILE._04785_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09772_  (.A0(\u_cpu.REG_FILE.rf[7][0] ),
    .A1(\u_cpu.REG_FILE._04642_ ),
    .S(\u_cpu.REG_FILE._04785_ ),
    .X(\u_cpu.REG_FILE._04786_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09773_  (.A(\u_cpu.REG_FILE._04786_ ),
    .X(\u_cpu.REG_FILE._00256_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09774_  (.A0(\u_cpu.REG_FILE.rf[7][1] ),
    .A1(\u_cpu.REG_FILE._04647_ ),
    .S(\u_cpu.REG_FILE._04785_ ),
    .X(\u_cpu.REG_FILE._04787_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09775_  (.A(\u_cpu.REG_FILE._04787_ ),
    .X(\u_cpu.REG_FILE._00257_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09776_  (.A0(\u_cpu.REG_FILE.rf[7][2] ),
    .A1(\u_cpu.REG_FILE._04649_ ),
    .S(\u_cpu.REG_FILE._04785_ ),
    .X(\u_cpu.REG_FILE._04788_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09777_  (.A(\u_cpu.REG_FILE._04788_ ),
    .X(\u_cpu.REG_FILE._00258_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09778_  (.A0(\u_cpu.REG_FILE.rf[7][3] ),
    .A1(\u_cpu.REG_FILE._04651_ ),
    .S(\u_cpu.REG_FILE._04785_ ),
    .X(\u_cpu.REG_FILE._04789_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09779_  (.A(\u_cpu.REG_FILE._04789_ ),
    .X(\u_cpu.REG_FILE._00259_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09780_  (.A0(\u_cpu.REG_FILE.rf[7][4] ),
    .A1(\u_cpu.REG_FILE._04653_ ),
    .S(\u_cpu.REG_FILE._04785_ ),
    .X(\u_cpu.REG_FILE._04790_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09781_  (.A(\u_cpu.REG_FILE._04790_ ),
    .X(\u_cpu.REG_FILE._00260_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09782_  (.A0(\u_cpu.REG_FILE.rf[7][5] ),
    .A1(\u_cpu.REG_FILE._04655_ ),
    .S(\u_cpu.REG_FILE._04785_ ),
    .X(\u_cpu.REG_FILE._04791_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09783_  (.A(\u_cpu.REG_FILE._04791_ ),
    .X(\u_cpu.REG_FILE._00261_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09784_  (.A0(\u_cpu.REG_FILE.rf[7][6] ),
    .A1(\u_cpu.REG_FILE._04657_ ),
    .S(\u_cpu.REG_FILE._04785_ ),
    .X(\u_cpu.REG_FILE._04792_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09785_  (.A(\u_cpu.REG_FILE._04792_ ),
    .X(\u_cpu.REG_FILE._00262_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09786_  (.A0(\u_cpu.REG_FILE.rf[7][7] ),
    .A1(\u_cpu.REG_FILE._04659_ ),
    .S(\u_cpu.REG_FILE._04785_ ),
    .X(\u_cpu.REG_FILE._04793_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09787_  (.A(\u_cpu.REG_FILE._04793_ ),
    .X(\u_cpu.REG_FILE._00263_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09788_  (.A0(\u_cpu.REG_FILE.rf[7][8] ),
    .A1(\u_cpu.REG_FILE._04661_ ),
    .S(\u_cpu.REG_FILE._04785_ ),
    .X(\u_cpu.REG_FILE._04794_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09789_  (.A(\u_cpu.REG_FILE._04794_ ),
    .X(\u_cpu.REG_FILE._00264_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09790_  (.A0(\u_cpu.REG_FILE.rf[7][9] ),
    .A1(\u_cpu.REG_FILE._04663_ ),
    .S(\u_cpu.REG_FILE._04785_ ),
    .X(\u_cpu.REG_FILE._04795_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09791_  (.A(\u_cpu.REG_FILE._04795_ ),
    .X(\u_cpu.REG_FILE._00265_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09792_  (.A(\u_cpu.REG_FILE._04784_ ),
    .X(\u_cpu.REG_FILE._04796_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09793_  (.A0(\u_cpu.REG_FILE.rf[7][10] ),
    .A1(\u_cpu.REG_FILE._04665_ ),
    .S(\u_cpu.REG_FILE._04796_ ),
    .X(\u_cpu.REG_FILE._04797_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09794_  (.A(\u_cpu.REG_FILE._04797_ ),
    .X(\u_cpu.REG_FILE._00266_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09795_  (.A0(\u_cpu.REG_FILE.rf[7][11] ),
    .A1(\u_cpu.REG_FILE._04668_ ),
    .S(\u_cpu.REG_FILE._04796_ ),
    .X(\u_cpu.REG_FILE._04798_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09796_  (.A(\u_cpu.REG_FILE._04798_ ),
    .X(\u_cpu.REG_FILE._00267_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09797_  (.A0(\u_cpu.REG_FILE.rf[7][12] ),
    .A1(\u_cpu.REG_FILE._04670_ ),
    .S(\u_cpu.REG_FILE._04796_ ),
    .X(\u_cpu.REG_FILE._04799_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09798_  (.A(\u_cpu.REG_FILE._04799_ ),
    .X(\u_cpu.REG_FILE._00268_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09799_  (.A0(\u_cpu.REG_FILE.rf[7][13] ),
    .A1(\u_cpu.REG_FILE._04672_ ),
    .S(\u_cpu.REG_FILE._04796_ ),
    .X(\u_cpu.REG_FILE._04800_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09800_  (.A(\u_cpu.REG_FILE._04800_ ),
    .X(\u_cpu.REG_FILE._00269_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09801_  (.A0(\u_cpu.REG_FILE.rf[7][14] ),
    .A1(\u_cpu.REG_FILE._04674_ ),
    .S(\u_cpu.REG_FILE._04796_ ),
    .X(\u_cpu.REG_FILE._04801_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09802_  (.A(\u_cpu.REG_FILE._04801_ ),
    .X(\u_cpu.REG_FILE._00270_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09803_  (.A0(\u_cpu.REG_FILE.rf[7][15] ),
    .A1(\u_cpu.REG_FILE._04676_ ),
    .S(\u_cpu.REG_FILE._04796_ ),
    .X(\u_cpu.REG_FILE._04802_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09804_  (.A(\u_cpu.REG_FILE._04802_ ),
    .X(\u_cpu.REG_FILE._00271_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09805_  (.A0(\u_cpu.REG_FILE.rf[7][16] ),
    .A1(\u_cpu.REG_FILE._04678_ ),
    .S(\u_cpu.REG_FILE._04796_ ),
    .X(\u_cpu.REG_FILE._04803_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09806_  (.A(\u_cpu.REG_FILE._04803_ ),
    .X(\u_cpu.REG_FILE._00272_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09807_  (.A0(\u_cpu.REG_FILE.rf[7][17] ),
    .A1(\u_cpu.REG_FILE._04680_ ),
    .S(\u_cpu.REG_FILE._04796_ ),
    .X(\u_cpu.REG_FILE._04804_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09808_  (.A(\u_cpu.REG_FILE._04804_ ),
    .X(\u_cpu.REG_FILE._00273_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09809_  (.A0(\u_cpu.REG_FILE.rf[7][18] ),
    .A1(\u_cpu.REG_FILE._04682_ ),
    .S(\u_cpu.REG_FILE._04796_ ),
    .X(\u_cpu.REG_FILE._04805_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09810_  (.A(\u_cpu.REG_FILE._04805_ ),
    .X(\u_cpu.REG_FILE._00274_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09811_  (.A0(\u_cpu.REG_FILE.rf[7][19] ),
    .A1(\u_cpu.REG_FILE._04684_ ),
    .S(\u_cpu.REG_FILE._04796_ ),
    .X(\u_cpu.REG_FILE._04806_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09812_  (.A(\u_cpu.REG_FILE._04806_ ),
    .X(\u_cpu.REG_FILE._00275_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09813_  (.A(\u_cpu.REG_FILE._04784_ ),
    .X(\u_cpu.REG_FILE._04807_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09814_  (.A0(\u_cpu.REG_FILE.rf[7][20] ),
    .A1(\u_cpu.REG_FILE._04686_ ),
    .S(\u_cpu.REG_FILE._04807_ ),
    .X(\u_cpu.REG_FILE._04808_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09815_  (.A(\u_cpu.REG_FILE._04808_ ),
    .X(\u_cpu.REG_FILE._00276_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09816_  (.A0(\u_cpu.REG_FILE.rf[7][21] ),
    .A1(\u_cpu.REG_FILE._04689_ ),
    .S(\u_cpu.REG_FILE._04807_ ),
    .X(\u_cpu.REG_FILE._04809_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09817_  (.A(\u_cpu.REG_FILE._04809_ ),
    .X(\u_cpu.REG_FILE._00277_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09818_  (.A0(\u_cpu.REG_FILE.rf[7][22] ),
    .A1(\u_cpu.REG_FILE._04691_ ),
    .S(\u_cpu.REG_FILE._04807_ ),
    .X(\u_cpu.REG_FILE._04810_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09819_  (.A(\u_cpu.REG_FILE._04810_ ),
    .X(\u_cpu.REG_FILE._00278_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09820_  (.A0(\u_cpu.REG_FILE.rf[7][23] ),
    .A1(\u_cpu.REG_FILE._04693_ ),
    .S(\u_cpu.REG_FILE._04807_ ),
    .X(\u_cpu.REG_FILE._04811_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09821_  (.A(\u_cpu.REG_FILE._04811_ ),
    .X(\u_cpu.REG_FILE._00279_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09822_  (.A0(\u_cpu.REG_FILE.rf[7][24] ),
    .A1(\u_cpu.REG_FILE._04695_ ),
    .S(\u_cpu.REG_FILE._04807_ ),
    .X(\u_cpu.REG_FILE._04812_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09823_  (.A(\u_cpu.REG_FILE._04812_ ),
    .X(\u_cpu.REG_FILE._00280_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09824_  (.A0(\u_cpu.REG_FILE.rf[7][25] ),
    .A1(\u_cpu.REG_FILE._04697_ ),
    .S(\u_cpu.REG_FILE._04807_ ),
    .X(\u_cpu.REG_FILE._04813_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09825_  (.A(\u_cpu.REG_FILE._04813_ ),
    .X(\u_cpu.REG_FILE._00281_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09826_  (.A0(\u_cpu.REG_FILE.rf[7][26] ),
    .A1(\u_cpu.REG_FILE._04699_ ),
    .S(\u_cpu.REG_FILE._04807_ ),
    .X(\u_cpu.REG_FILE._04814_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09827_  (.A(\u_cpu.REG_FILE._04814_ ),
    .X(\u_cpu.REG_FILE._00282_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09828_  (.A0(\u_cpu.REG_FILE.rf[7][27] ),
    .A1(\u_cpu.REG_FILE._04701_ ),
    .S(\u_cpu.REG_FILE._04807_ ),
    .X(\u_cpu.REG_FILE._04815_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09829_  (.A(\u_cpu.REG_FILE._04815_ ),
    .X(\u_cpu.REG_FILE._00283_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09830_  (.A0(\u_cpu.REG_FILE.rf[7][28] ),
    .A1(\u_cpu.REG_FILE._04703_ ),
    .S(\u_cpu.REG_FILE._04807_ ),
    .X(\u_cpu.REG_FILE._04816_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09831_  (.A(\u_cpu.REG_FILE._04816_ ),
    .X(\u_cpu.REG_FILE._00284_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09832_  (.A0(\u_cpu.REG_FILE.rf[7][29] ),
    .A1(\u_cpu.REG_FILE._04705_ ),
    .S(\u_cpu.REG_FILE._04807_ ),
    .X(\u_cpu.REG_FILE._04817_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09833_  (.A(\u_cpu.REG_FILE._04817_ ),
    .X(\u_cpu.REG_FILE._00285_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09834_  (.A0(\u_cpu.REG_FILE.rf[7][30] ),
    .A1(\u_cpu.REG_FILE._04707_ ),
    .S(\u_cpu.REG_FILE._04784_ ),
    .X(\u_cpu.REG_FILE._04818_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09835_  (.A(\u_cpu.REG_FILE._04818_ ),
    .X(\u_cpu.REG_FILE._00286_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09836_  (.A0(\u_cpu.REG_FILE.rf[7][31] ),
    .A1(\u_cpu.REG_FILE._04709_ ),
    .S(\u_cpu.REG_FILE._04784_ ),
    .X(\u_cpu.REG_FILE._04819_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09837_  (.A(\u_cpu.REG_FILE._04819_ ),
    .X(\u_cpu.REG_FILE._00287_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.REG_FILE._09838_  (.A(\u_cpu.REG_FILE._04422_ ),
    .B(\u_cpu.REG_FILE._04426_ ),
    .C(\u_cpu.REG_FILE._04643_ ),
    .X(\u_cpu.REG_FILE._04820_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09839_  (.A(\u_cpu.REG_FILE._04820_ ),
    .X(\u_cpu.REG_FILE._04821_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09840_  (.A0(\u_cpu.REG_FILE.rf[8][0] ),
    .A1(\u_cpu.REG_FILE._04642_ ),
    .S(\u_cpu.REG_FILE._04821_ ),
    .X(\u_cpu.REG_FILE._04822_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09841_  (.A(\u_cpu.REG_FILE._04822_ ),
    .X(\u_cpu.REG_FILE._00288_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09842_  (.A0(\u_cpu.REG_FILE.rf[8][1] ),
    .A1(\u_cpu.REG_FILE._04647_ ),
    .S(\u_cpu.REG_FILE._04821_ ),
    .X(\u_cpu.REG_FILE._04823_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09843_  (.A(\u_cpu.REG_FILE._04823_ ),
    .X(\u_cpu.REG_FILE._00289_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09844_  (.A0(\u_cpu.REG_FILE.rf[8][2] ),
    .A1(\u_cpu.REG_FILE._04649_ ),
    .S(\u_cpu.REG_FILE._04821_ ),
    .X(\u_cpu.REG_FILE._04824_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09845_  (.A(\u_cpu.REG_FILE._04824_ ),
    .X(\u_cpu.REG_FILE._00290_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09846_  (.A0(\u_cpu.REG_FILE.rf[8][3] ),
    .A1(\u_cpu.REG_FILE._04651_ ),
    .S(\u_cpu.REG_FILE._04821_ ),
    .X(\u_cpu.REG_FILE._04825_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09847_  (.A(\u_cpu.REG_FILE._04825_ ),
    .X(\u_cpu.REG_FILE._00291_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09848_  (.A0(\u_cpu.REG_FILE.rf[8][4] ),
    .A1(\u_cpu.REG_FILE._04653_ ),
    .S(\u_cpu.REG_FILE._04821_ ),
    .X(\u_cpu.REG_FILE._04826_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09849_  (.A(\u_cpu.REG_FILE._04826_ ),
    .X(\u_cpu.REG_FILE._00292_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09850_  (.A0(\u_cpu.REG_FILE.rf[8][5] ),
    .A1(\u_cpu.REG_FILE._04655_ ),
    .S(\u_cpu.REG_FILE._04821_ ),
    .X(\u_cpu.REG_FILE._04827_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09851_  (.A(\u_cpu.REG_FILE._04827_ ),
    .X(\u_cpu.REG_FILE._00293_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09852_  (.A0(\u_cpu.REG_FILE.rf[8][6] ),
    .A1(\u_cpu.REG_FILE._04657_ ),
    .S(\u_cpu.REG_FILE._04821_ ),
    .X(\u_cpu.REG_FILE._04828_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09853_  (.A(\u_cpu.REG_FILE._04828_ ),
    .X(\u_cpu.REG_FILE._00294_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09854_  (.A0(\u_cpu.REG_FILE.rf[8][7] ),
    .A1(\u_cpu.REG_FILE._04659_ ),
    .S(\u_cpu.REG_FILE._04821_ ),
    .X(\u_cpu.REG_FILE._04829_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09855_  (.A(\u_cpu.REG_FILE._04829_ ),
    .X(\u_cpu.REG_FILE._00295_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09856_  (.A0(\u_cpu.REG_FILE.rf[8][8] ),
    .A1(\u_cpu.REG_FILE._04661_ ),
    .S(\u_cpu.REG_FILE._04821_ ),
    .X(\u_cpu.REG_FILE._04830_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09857_  (.A(\u_cpu.REG_FILE._04830_ ),
    .X(\u_cpu.REG_FILE._00296_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09858_  (.A0(\u_cpu.REG_FILE.rf[8][9] ),
    .A1(\u_cpu.REG_FILE._04663_ ),
    .S(\u_cpu.REG_FILE._04821_ ),
    .X(\u_cpu.REG_FILE._04831_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09859_  (.A(\u_cpu.REG_FILE._04831_ ),
    .X(\u_cpu.REG_FILE._00297_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09860_  (.A(\u_cpu.REG_FILE._04820_ ),
    .X(\u_cpu.REG_FILE._04832_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09861_  (.A0(\u_cpu.REG_FILE.rf[8][10] ),
    .A1(\u_cpu.REG_FILE._04665_ ),
    .S(\u_cpu.REG_FILE._04832_ ),
    .X(\u_cpu.REG_FILE._04833_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09862_  (.A(\u_cpu.REG_FILE._04833_ ),
    .X(\u_cpu.REG_FILE._00298_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09863_  (.A0(\u_cpu.REG_FILE.rf[8][11] ),
    .A1(\u_cpu.REG_FILE._04668_ ),
    .S(\u_cpu.REG_FILE._04832_ ),
    .X(\u_cpu.REG_FILE._04834_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09864_  (.A(\u_cpu.REG_FILE._04834_ ),
    .X(\u_cpu.REG_FILE._00299_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09865_  (.A0(\u_cpu.REG_FILE.rf[8][12] ),
    .A1(\u_cpu.REG_FILE._04670_ ),
    .S(\u_cpu.REG_FILE._04832_ ),
    .X(\u_cpu.REG_FILE._04835_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09866_  (.A(\u_cpu.REG_FILE._04835_ ),
    .X(\u_cpu.REG_FILE._00300_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09867_  (.A0(\u_cpu.REG_FILE.rf[8][13] ),
    .A1(\u_cpu.REG_FILE._04672_ ),
    .S(\u_cpu.REG_FILE._04832_ ),
    .X(\u_cpu.REG_FILE._04836_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09868_  (.A(\u_cpu.REG_FILE._04836_ ),
    .X(\u_cpu.REG_FILE._00301_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09869_  (.A0(\u_cpu.REG_FILE.rf[8][14] ),
    .A1(\u_cpu.REG_FILE._04674_ ),
    .S(\u_cpu.REG_FILE._04832_ ),
    .X(\u_cpu.REG_FILE._04837_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09870_  (.A(\u_cpu.REG_FILE._04837_ ),
    .X(\u_cpu.REG_FILE._00302_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09871_  (.A0(\u_cpu.REG_FILE.rf[8][15] ),
    .A1(\u_cpu.REG_FILE._04676_ ),
    .S(\u_cpu.REG_FILE._04832_ ),
    .X(\u_cpu.REG_FILE._04838_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09872_  (.A(\u_cpu.REG_FILE._04838_ ),
    .X(\u_cpu.REG_FILE._00303_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09873_  (.A0(\u_cpu.REG_FILE.rf[8][16] ),
    .A1(\u_cpu.REG_FILE._04678_ ),
    .S(\u_cpu.REG_FILE._04832_ ),
    .X(\u_cpu.REG_FILE._04839_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09874_  (.A(\u_cpu.REG_FILE._04839_ ),
    .X(\u_cpu.REG_FILE._00304_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09875_  (.A0(\u_cpu.REG_FILE.rf[8][17] ),
    .A1(\u_cpu.REG_FILE._04680_ ),
    .S(\u_cpu.REG_FILE._04832_ ),
    .X(\u_cpu.REG_FILE._04840_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09876_  (.A(\u_cpu.REG_FILE._04840_ ),
    .X(\u_cpu.REG_FILE._00305_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09877_  (.A0(\u_cpu.REG_FILE.rf[8][18] ),
    .A1(\u_cpu.REG_FILE._04682_ ),
    .S(\u_cpu.REG_FILE._04832_ ),
    .X(\u_cpu.REG_FILE._04841_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09878_  (.A(\u_cpu.REG_FILE._04841_ ),
    .X(\u_cpu.REG_FILE._00306_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09879_  (.A0(\u_cpu.REG_FILE.rf[8][19] ),
    .A1(\u_cpu.REG_FILE._04684_ ),
    .S(\u_cpu.REG_FILE._04832_ ),
    .X(\u_cpu.REG_FILE._04842_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09880_  (.A(\u_cpu.REG_FILE._04842_ ),
    .X(\u_cpu.REG_FILE._00307_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09881_  (.A(\u_cpu.REG_FILE._04820_ ),
    .X(\u_cpu.REG_FILE._04843_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09882_  (.A0(\u_cpu.REG_FILE.rf[8][20] ),
    .A1(\u_cpu.REG_FILE._04686_ ),
    .S(\u_cpu.REG_FILE._04843_ ),
    .X(\u_cpu.REG_FILE._04844_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09883_  (.A(\u_cpu.REG_FILE._04844_ ),
    .X(\u_cpu.REG_FILE._00308_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09884_  (.A0(\u_cpu.REG_FILE.rf[8][21] ),
    .A1(\u_cpu.REG_FILE._04689_ ),
    .S(\u_cpu.REG_FILE._04843_ ),
    .X(\u_cpu.REG_FILE._04845_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09885_  (.A(\u_cpu.REG_FILE._04845_ ),
    .X(\u_cpu.REG_FILE._00309_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09886_  (.A0(\u_cpu.REG_FILE.rf[8][22] ),
    .A1(\u_cpu.REG_FILE._04691_ ),
    .S(\u_cpu.REG_FILE._04843_ ),
    .X(\u_cpu.REG_FILE._04846_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09887_  (.A(\u_cpu.REG_FILE._04846_ ),
    .X(\u_cpu.REG_FILE._00310_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09888_  (.A0(\u_cpu.REG_FILE.rf[8][23] ),
    .A1(\u_cpu.REG_FILE._04693_ ),
    .S(\u_cpu.REG_FILE._04843_ ),
    .X(\u_cpu.REG_FILE._04847_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09889_  (.A(\u_cpu.REG_FILE._04847_ ),
    .X(\u_cpu.REG_FILE._00311_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09890_  (.A0(\u_cpu.REG_FILE.rf[8][24] ),
    .A1(\u_cpu.REG_FILE._04695_ ),
    .S(\u_cpu.REG_FILE._04843_ ),
    .X(\u_cpu.REG_FILE._04848_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09891_  (.A(\u_cpu.REG_FILE._04848_ ),
    .X(\u_cpu.REG_FILE._00312_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09892_  (.A0(\u_cpu.REG_FILE.rf[8][25] ),
    .A1(\u_cpu.REG_FILE._04697_ ),
    .S(\u_cpu.REG_FILE._04843_ ),
    .X(\u_cpu.REG_FILE._04849_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09893_  (.A(\u_cpu.REG_FILE._04849_ ),
    .X(\u_cpu.REG_FILE._00313_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09894_  (.A0(\u_cpu.REG_FILE.rf[8][26] ),
    .A1(\u_cpu.REG_FILE._04699_ ),
    .S(\u_cpu.REG_FILE._04843_ ),
    .X(\u_cpu.REG_FILE._04850_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09895_  (.A(\u_cpu.REG_FILE._04850_ ),
    .X(\u_cpu.REG_FILE._00314_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09896_  (.A0(\u_cpu.REG_FILE.rf[8][27] ),
    .A1(\u_cpu.REG_FILE._04701_ ),
    .S(\u_cpu.REG_FILE._04843_ ),
    .X(\u_cpu.REG_FILE._04851_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09897_  (.A(\u_cpu.REG_FILE._04851_ ),
    .X(\u_cpu.REG_FILE._00315_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09898_  (.A0(\u_cpu.REG_FILE.rf[8][28] ),
    .A1(\u_cpu.REG_FILE._04703_ ),
    .S(\u_cpu.REG_FILE._04843_ ),
    .X(\u_cpu.REG_FILE._04852_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09899_  (.A(\u_cpu.REG_FILE._04852_ ),
    .X(\u_cpu.REG_FILE._00316_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09900_  (.A0(\u_cpu.REG_FILE.rf[8][29] ),
    .A1(\u_cpu.REG_FILE._04705_ ),
    .S(\u_cpu.REG_FILE._04843_ ),
    .X(\u_cpu.REG_FILE._04853_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09901_  (.A(\u_cpu.REG_FILE._04853_ ),
    .X(\u_cpu.REG_FILE._00317_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09902_  (.A0(\u_cpu.REG_FILE.rf[8][30] ),
    .A1(\u_cpu.REG_FILE._04707_ ),
    .S(\u_cpu.REG_FILE._04820_ ),
    .X(\u_cpu.REG_FILE._04854_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09903_  (.A(\u_cpu.REG_FILE._04854_ ),
    .X(\u_cpu.REG_FILE._00318_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09904_  (.A0(\u_cpu.REG_FILE.rf[8][31] ),
    .A1(\u_cpu.REG_FILE._04709_ ),
    .S(\u_cpu.REG_FILE._04820_ ),
    .X(\u_cpu.REG_FILE._04855_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09905_  (.A(\u_cpu.REG_FILE._04855_ ),
    .X(\u_cpu.REG_FILE._00319_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09906_  (.A(\u_cpu.REG_FILE.rf[0][0] ),
    .X(\u_cpu.REG_FILE._04856_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09907_  (.A(\u_cpu.REG_FILE._04856_ ),
    .X(\u_cpu.REG_FILE._00320_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09908_  (.A(\u_cpu.REG_FILE.rf[0][1] ),
    .X(\u_cpu.REG_FILE._04857_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09909_  (.A(\u_cpu.REG_FILE._04857_ ),
    .X(\u_cpu.REG_FILE._00321_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09910_  (.A(\u_cpu.REG_FILE.rf[0][2] ),
    .X(\u_cpu.REG_FILE._04858_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09911_  (.A(\u_cpu.REG_FILE._04858_ ),
    .X(\u_cpu.REG_FILE._00322_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09912_  (.A(\u_cpu.REG_FILE.rf[0][3] ),
    .X(\u_cpu.REG_FILE._04859_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09913_  (.A(\u_cpu.REG_FILE._04859_ ),
    .X(\u_cpu.REG_FILE._00323_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09914_  (.A(\u_cpu.REG_FILE.rf[0][4] ),
    .X(\u_cpu.REG_FILE._04860_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09915_  (.A(\u_cpu.REG_FILE._04860_ ),
    .X(\u_cpu.REG_FILE._00324_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09916_  (.A(\u_cpu.REG_FILE.rf[0][5] ),
    .X(\u_cpu.REG_FILE._04861_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09917_  (.A(\u_cpu.REG_FILE._04861_ ),
    .X(\u_cpu.REG_FILE._00325_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09918_  (.A(\u_cpu.REG_FILE.rf[0][6] ),
    .X(\u_cpu.REG_FILE._04862_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09919_  (.A(\u_cpu.REG_FILE._04862_ ),
    .X(\u_cpu.REG_FILE._00326_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09920_  (.A(\u_cpu.REG_FILE.rf[0][7] ),
    .X(\u_cpu.REG_FILE._04863_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09921_  (.A(\u_cpu.REG_FILE._04863_ ),
    .X(\u_cpu.REG_FILE._00327_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09922_  (.A(\u_cpu.REG_FILE.rf[0][8] ),
    .X(\u_cpu.REG_FILE._04864_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09923_  (.A(\u_cpu.REG_FILE._04864_ ),
    .X(\u_cpu.REG_FILE._00328_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09924_  (.A(\u_cpu.REG_FILE.rf[0][9] ),
    .X(\u_cpu.REG_FILE._04865_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09925_  (.A(\u_cpu.REG_FILE._04865_ ),
    .X(\u_cpu.REG_FILE._00329_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09926_  (.A(\u_cpu.REG_FILE.rf[0][10] ),
    .X(\u_cpu.REG_FILE._04866_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09927_  (.A(\u_cpu.REG_FILE._04866_ ),
    .X(\u_cpu.REG_FILE._00330_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09928_  (.A(\u_cpu.REG_FILE.rf[0][11] ),
    .X(\u_cpu.REG_FILE._04867_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09929_  (.A(\u_cpu.REG_FILE._04867_ ),
    .X(\u_cpu.REG_FILE._00331_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09930_  (.A(\u_cpu.REG_FILE.rf[0][12] ),
    .X(\u_cpu.REG_FILE._04868_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09931_  (.A(\u_cpu.REG_FILE._04868_ ),
    .X(\u_cpu.REG_FILE._00332_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09932_  (.A(\u_cpu.REG_FILE.rf[0][13] ),
    .X(\u_cpu.REG_FILE._04869_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09933_  (.A(\u_cpu.REG_FILE._04869_ ),
    .X(\u_cpu.REG_FILE._00333_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09934_  (.A(\u_cpu.REG_FILE.rf[0][14] ),
    .X(\u_cpu.REG_FILE._04870_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09935_  (.A(\u_cpu.REG_FILE._04870_ ),
    .X(\u_cpu.REG_FILE._00334_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09936_  (.A(\u_cpu.REG_FILE.rf[0][15] ),
    .X(\u_cpu.REG_FILE._04871_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09937_  (.A(\u_cpu.REG_FILE._04871_ ),
    .X(\u_cpu.REG_FILE._00335_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09938_  (.A(\u_cpu.REG_FILE.rf[0][16] ),
    .X(\u_cpu.REG_FILE._04872_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09939_  (.A(\u_cpu.REG_FILE._04872_ ),
    .X(\u_cpu.REG_FILE._00336_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09940_  (.A(\u_cpu.REG_FILE.rf[0][17] ),
    .X(\u_cpu.REG_FILE._04873_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09941_  (.A(\u_cpu.REG_FILE._04873_ ),
    .X(\u_cpu.REG_FILE._00337_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09942_  (.A(\u_cpu.REG_FILE.rf[0][18] ),
    .X(\u_cpu.REG_FILE._04874_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09943_  (.A(\u_cpu.REG_FILE._04874_ ),
    .X(\u_cpu.REG_FILE._00338_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09944_  (.A(\u_cpu.REG_FILE.rf[0][19] ),
    .X(\u_cpu.REG_FILE._04875_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09945_  (.A(\u_cpu.REG_FILE._04875_ ),
    .X(\u_cpu.REG_FILE._00339_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09946_  (.A(\u_cpu.REG_FILE.rf[0][20] ),
    .X(\u_cpu.REG_FILE._04876_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09947_  (.A(\u_cpu.REG_FILE._04876_ ),
    .X(\u_cpu.REG_FILE._00340_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09948_  (.A(\u_cpu.REG_FILE.rf[0][21] ),
    .X(\u_cpu.REG_FILE._04877_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09949_  (.A(\u_cpu.REG_FILE._04877_ ),
    .X(\u_cpu.REG_FILE._00341_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09950_  (.A(\u_cpu.REG_FILE.rf[0][22] ),
    .X(\u_cpu.REG_FILE._04878_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09951_  (.A(\u_cpu.REG_FILE._04878_ ),
    .X(\u_cpu.REG_FILE._00342_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09952_  (.A(\u_cpu.REG_FILE.rf[0][23] ),
    .X(\u_cpu.REG_FILE._04879_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09953_  (.A(\u_cpu.REG_FILE._04879_ ),
    .X(\u_cpu.REG_FILE._00343_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09954_  (.A(\u_cpu.REG_FILE.rf[0][24] ),
    .X(\u_cpu.REG_FILE._04880_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09955_  (.A(\u_cpu.REG_FILE._04880_ ),
    .X(\u_cpu.REG_FILE._00344_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09956_  (.A(\u_cpu.REG_FILE.rf[0][25] ),
    .X(\u_cpu.REG_FILE._04881_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09957_  (.A(\u_cpu.REG_FILE._04881_ ),
    .X(\u_cpu.REG_FILE._00345_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09958_  (.A(\u_cpu.REG_FILE.rf[0][26] ),
    .X(\u_cpu.REG_FILE._04882_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09959_  (.A(\u_cpu.REG_FILE._04882_ ),
    .X(\u_cpu.REG_FILE._00346_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09960_  (.A(\u_cpu.REG_FILE.rf[0][27] ),
    .X(\u_cpu.REG_FILE._04883_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09961_  (.A(\u_cpu.REG_FILE._04883_ ),
    .X(\u_cpu.REG_FILE._00347_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09962_  (.A(\u_cpu.REG_FILE.rf[0][28] ),
    .X(\u_cpu.REG_FILE._04884_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09963_  (.A(\u_cpu.REG_FILE._04884_ ),
    .X(\u_cpu.REG_FILE._00348_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09964_  (.A(\u_cpu.REG_FILE.rf[0][29] ),
    .X(\u_cpu.REG_FILE._04885_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09965_  (.A(\u_cpu.REG_FILE._04885_ ),
    .X(\u_cpu.REG_FILE._00349_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09966_  (.A(\u_cpu.REG_FILE.rf[0][30] ),
    .X(\u_cpu.REG_FILE._04886_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09967_  (.A(\u_cpu.REG_FILE._04886_ ),
    .X(\u_cpu.REG_FILE._00350_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09968_  (.A(\u_cpu.REG_FILE.rf[0][31] ),
    .X(\u_cpu.REG_FILE._04887_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09969_  (.A(\u_cpu.REG_FILE._04887_ ),
    .X(\u_cpu.REG_FILE._00351_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.REG_FILE._09970_  (.A(\u_cpu.REG_FILE._04422_ ),
    .B(\u_cpu.REG_FILE._04426_ ),
    .C(\u_cpu.REG_FILE._04747_ ),
    .X(\u_cpu.REG_FILE._04888_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09971_  (.A(\u_cpu.REG_FILE._04888_ ),
    .X(\u_cpu.REG_FILE._04889_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09972_  (.A0(\u_cpu.REG_FILE.rf[10][0] ),
    .A1(\u_cpu.REG_FILE._04642_ ),
    .S(\u_cpu.REG_FILE._04889_ ),
    .X(\u_cpu.REG_FILE._04890_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09973_  (.A(\u_cpu.REG_FILE._04890_ ),
    .X(\u_cpu.REG_FILE._00352_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09974_  (.A0(\u_cpu.REG_FILE.rf[10][1] ),
    .A1(\u_cpu.REG_FILE._04647_ ),
    .S(\u_cpu.REG_FILE._04889_ ),
    .X(\u_cpu.REG_FILE._04891_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09975_  (.A(\u_cpu.REG_FILE._04891_ ),
    .X(\u_cpu.REG_FILE._00353_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09976_  (.A0(\u_cpu.REG_FILE.rf[10][2] ),
    .A1(\u_cpu.REG_FILE._04649_ ),
    .S(\u_cpu.REG_FILE._04889_ ),
    .X(\u_cpu.REG_FILE._04892_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09977_  (.A(\u_cpu.REG_FILE._04892_ ),
    .X(\u_cpu.REG_FILE._00354_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09978_  (.A0(\u_cpu.REG_FILE.rf[10][3] ),
    .A1(\u_cpu.REG_FILE._04651_ ),
    .S(\u_cpu.REG_FILE._04889_ ),
    .X(\u_cpu.REG_FILE._04893_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09979_  (.A(\u_cpu.REG_FILE._04893_ ),
    .X(\u_cpu.REG_FILE._00355_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09980_  (.A0(\u_cpu.REG_FILE.rf[10][4] ),
    .A1(\u_cpu.REG_FILE._04653_ ),
    .S(\u_cpu.REG_FILE._04889_ ),
    .X(\u_cpu.REG_FILE._04894_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09981_  (.A(\u_cpu.REG_FILE._04894_ ),
    .X(\u_cpu.REG_FILE._00356_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09982_  (.A0(\u_cpu.REG_FILE.rf[10][5] ),
    .A1(\u_cpu.REG_FILE._04655_ ),
    .S(\u_cpu.REG_FILE._04889_ ),
    .X(\u_cpu.REG_FILE._04895_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09983_  (.A(\u_cpu.REG_FILE._04895_ ),
    .X(\u_cpu.REG_FILE._00357_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09984_  (.A0(\u_cpu.REG_FILE.rf[10][6] ),
    .A1(\u_cpu.REG_FILE._04657_ ),
    .S(\u_cpu.REG_FILE._04889_ ),
    .X(\u_cpu.REG_FILE._04896_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09985_  (.A(\u_cpu.REG_FILE._04896_ ),
    .X(\u_cpu.REG_FILE._00358_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09986_  (.A0(\u_cpu.REG_FILE.rf[10][7] ),
    .A1(\u_cpu.REG_FILE._04659_ ),
    .S(\u_cpu.REG_FILE._04889_ ),
    .X(\u_cpu.REG_FILE._04897_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09987_  (.A(\u_cpu.REG_FILE._04897_ ),
    .X(\u_cpu.REG_FILE._00359_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09988_  (.A0(\u_cpu.REG_FILE.rf[10][8] ),
    .A1(\u_cpu.REG_FILE._04661_ ),
    .S(\u_cpu.REG_FILE._04889_ ),
    .X(\u_cpu.REG_FILE._04898_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09989_  (.A(\u_cpu.REG_FILE._04898_ ),
    .X(\u_cpu.REG_FILE._00360_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09990_  (.A0(\u_cpu.REG_FILE.rf[10][9] ),
    .A1(\u_cpu.REG_FILE._04663_ ),
    .S(\u_cpu.REG_FILE._04889_ ),
    .X(\u_cpu.REG_FILE._04899_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09991_  (.A(\u_cpu.REG_FILE._04899_ ),
    .X(\u_cpu.REG_FILE._00361_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09992_  (.A(\u_cpu.REG_FILE._04888_ ),
    .X(\u_cpu.REG_FILE._04900_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09993_  (.A0(\u_cpu.REG_FILE.rf[10][10] ),
    .A1(\u_cpu.REG_FILE._04665_ ),
    .S(\u_cpu.REG_FILE._04900_ ),
    .X(\u_cpu.REG_FILE._04901_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09994_  (.A(\u_cpu.REG_FILE._04901_ ),
    .X(\u_cpu.REG_FILE._00362_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09995_  (.A0(\u_cpu.REG_FILE.rf[10][11] ),
    .A1(\u_cpu.REG_FILE._04668_ ),
    .S(\u_cpu.REG_FILE._04900_ ),
    .X(\u_cpu.REG_FILE._04902_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09996_  (.A(\u_cpu.REG_FILE._04902_ ),
    .X(\u_cpu.REG_FILE._00363_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09997_  (.A0(\u_cpu.REG_FILE.rf[10][12] ),
    .A1(\u_cpu.REG_FILE._04670_ ),
    .S(\u_cpu.REG_FILE._04900_ ),
    .X(\u_cpu.REG_FILE._04903_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._09998_  (.A(\u_cpu.REG_FILE._04903_ ),
    .X(\u_cpu.REG_FILE._00364_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._09999_  (.A0(\u_cpu.REG_FILE.rf[10][13] ),
    .A1(\u_cpu.REG_FILE._04672_ ),
    .S(\u_cpu.REG_FILE._04900_ ),
    .X(\u_cpu.REG_FILE._04904_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10000_  (.A(\u_cpu.REG_FILE._04904_ ),
    .X(\u_cpu.REG_FILE._00365_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10001_  (.A0(\u_cpu.REG_FILE.rf[10][14] ),
    .A1(\u_cpu.REG_FILE._04674_ ),
    .S(\u_cpu.REG_FILE._04900_ ),
    .X(\u_cpu.REG_FILE._04905_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10002_  (.A(\u_cpu.REG_FILE._04905_ ),
    .X(\u_cpu.REG_FILE._00366_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10003_  (.A0(\u_cpu.REG_FILE.rf[10][15] ),
    .A1(\u_cpu.REG_FILE._04676_ ),
    .S(\u_cpu.REG_FILE._04900_ ),
    .X(\u_cpu.REG_FILE._04906_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10004_  (.A(\u_cpu.REG_FILE._04906_ ),
    .X(\u_cpu.REG_FILE._00367_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10005_  (.A0(\u_cpu.REG_FILE.rf[10][16] ),
    .A1(\u_cpu.REG_FILE._04678_ ),
    .S(\u_cpu.REG_FILE._04900_ ),
    .X(\u_cpu.REG_FILE._04907_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10006_  (.A(\u_cpu.REG_FILE._04907_ ),
    .X(\u_cpu.REG_FILE._00368_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10007_  (.A0(\u_cpu.REG_FILE.rf[10][17] ),
    .A1(\u_cpu.REG_FILE._04680_ ),
    .S(\u_cpu.REG_FILE._04900_ ),
    .X(\u_cpu.REG_FILE._04908_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10008_  (.A(\u_cpu.REG_FILE._04908_ ),
    .X(\u_cpu.REG_FILE._00369_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10009_  (.A0(\u_cpu.REG_FILE.rf[10][18] ),
    .A1(\u_cpu.REG_FILE._04682_ ),
    .S(\u_cpu.REG_FILE._04900_ ),
    .X(\u_cpu.REG_FILE._04909_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10010_  (.A(\u_cpu.REG_FILE._04909_ ),
    .X(\u_cpu.REG_FILE._00370_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10011_  (.A0(\u_cpu.REG_FILE.rf[10][19] ),
    .A1(\u_cpu.REG_FILE._04684_ ),
    .S(\u_cpu.REG_FILE._04900_ ),
    .X(\u_cpu.REG_FILE._04910_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10012_  (.A(\u_cpu.REG_FILE._04910_ ),
    .X(\u_cpu.REG_FILE._00371_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10013_  (.A(\u_cpu.REG_FILE._04888_ ),
    .X(\u_cpu.REG_FILE._04911_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10014_  (.A0(\u_cpu.REG_FILE.rf[10][20] ),
    .A1(\u_cpu.REG_FILE._04686_ ),
    .S(\u_cpu.REG_FILE._04911_ ),
    .X(\u_cpu.REG_FILE._04912_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10015_  (.A(\u_cpu.REG_FILE._04912_ ),
    .X(\u_cpu.REG_FILE._00372_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10016_  (.A0(\u_cpu.REG_FILE.rf[10][21] ),
    .A1(\u_cpu.REG_FILE._04689_ ),
    .S(\u_cpu.REG_FILE._04911_ ),
    .X(\u_cpu.REG_FILE._04913_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10017_  (.A(\u_cpu.REG_FILE._04913_ ),
    .X(\u_cpu.REG_FILE._00373_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10018_  (.A0(\u_cpu.REG_FILE.rf[10][22] ),
    .A1(\u_cpu.REG_FILE._04691_ ),
    .S(\u_cpu.REG_FILE._04911_ ),
    .X(\u_cpu.REG_FILE._04914_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10019_  (.A(\u_cpu.REG_FILE._04914_ ),
    .X(\u_cpu.REG_FILE._00374_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10020_  (.A0(\u_cpu.REG_FILE.rf[10][23] ),
    .A1(\u_cpu.REG_FILE._04693_ ),
    .S(\u_cpu.REG_FILE._04911_ ),
    .X(\u_cpu.REG_FILE._04915_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10021_  (.A(\u_cpu.REG_FILE._04915_ ),
    .X(\u_cpu.REG_FILE._00375_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10022_  (.A0(\u_cpu.REG_FILE.rf[10][24] ),
    .A1(\u_cpu.REG_FILE._04695_ ),
    .S(\u_cpu.REG_FILE._04911_ ),
    .X(\u_cpu.REG_FILE._04916_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10023_  (.A(\u_cpu.REG_FILE._04916_ ),
    .X(\u_cpu.REG_FILE._00376_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10024_  (.A0(\u_cpu.REG_FILE.rf[10][25] ),
    .A1(\u_cpu.REG_FILE._04697_ ),
    .S(\u_cpu.REG_FILE._04911_ ),
    .X(\u_cpu.REG_FILE._04917_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10025_  (.A(\u_cpu.REG_FILE._04917_ ),
    .X(\u_cpu.REG_FILE._00377_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10026_  (.A0(\u_cpu.REG_FILE.rf[10][26] ),
    .A1(\u_cpu.REG_FILE._04699_ ),
    .S(\u_cpu.REG_FILE._04911_ ),
    .X(\u_cpu.REG_FILE._04918_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10027_  (.A(\u_cpu.REG_FILE._04918_ ),
    .X(\u_cpu.REG_FILE._00378_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10028_  (.A0(\u_cpu.REG_FILE.rf[10][27] ),
    .A1(\u_cpu.REG_FILE._04701_ ),
    .S(\u_cpu.REG_FILE._04911_ ),
    .X(\u_cpu.REG_FILE._04919_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10029_  (.A(\u_cpu.REG_FILE._04919_ ),
    .X(\u_cpu.REG_FILE._00379_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10030_  (.A0(\u_cpu.REG_FILE.rf[10][28] ),
    .A1(\u_cpu.REG_FILE._04703_ ),
    .S(\u_cpu.REG_FILE._04911_ ),
    .X(\u_cpu.REG_FILE._04920_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10031_  (.A(\u_cpu.REG_FILE._04920_ ),
    .X(\u_cpu.REG_FILE._00380_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10032_  (.A0(\u_cpu.REG_FILE.rf[10][29] ),
    .A1(\u_cpu.REG_FILE._04705_ ),
    .S(\u_cpu.REG_FILE._04911_ ),
    .X(\u_cpu.REG_FILE._04921_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10033_  (.A(\u_cpu.REG_FILE._04921_ ),
    .X(\u_cpu.REG_FILE._00381_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10034_  (.A0(\u_cpu.REG_FILE.rf[10][30] ),
    .A1(\u_cpu.REG_FILE._04707_ ),
    .S(\u_cpu.REG_FILE._04888_ ),
    .X(\u_cpu.REG_FILE._04922_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10035_  (.A(\u_cpu.REG_FILE._04922_ ),
    .X(\u_cpu.REG_FILE._00382_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10036_  (.A0(\u_cpu.REG_FILE.rf[10][31] ),
    .A1(\u_cpu.REG_FILE._04709_ ),
    .S(\u_cpu.REG_FILE._04888_ ),
    .X(\u_cpu.REG_FILE._04923_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10037_  (.A(\u_cpu.REG_FILE._04923_ ),
    .X(\u_cpu.REG_FILE._00383_ ));
 sky130_fd_sc_hd__or4bb_2 \u_cpu.REG_FILE._10038_  (.A(\u_cpu.REG_FILE._04424_ ),
    .B(\u_cpu.REG_FILE._04494_ ),
    .C_N(\u_cpu.REG_FILE._04495_ ),
    .D_N(\u_cpu.REG_FILE._04422_ ),
    .X(\u_cpu.REG_FILE._04924_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10039_  (.A(\u_cpu.REG_FILE._04924_ ),
    .X(\u_cpu.REG_FILE._04925_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10040_  (.A0(\u_cpu.REG_FILE._04420_ ),
    .A1(\u_cpu.REG_FILE.rf[11][0] ),
    .S(\u_cpu.REG_FILE._04925_ ),
    .X(\u_cpu.REG_FILE._04926_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10041_  (.A(\u_cpu.REG_FILE._04926_ ),
    .X(\u_cpu.REG_FILE._00384_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10042_  (.A0(\u_cpu.REG_FILE._04430_ ),
    .A1(\u_cpu.REG_FILE.rf[11][1] ),
    .S(\u_cpu.REG_FILE._04925_ ),
    .X(\u_cpu.REG_FILE._04927_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10043_  (.A(\u_cpu.REG_FILE._04927_ ),
    .X(\u_cpu.REG_FILE._00385_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10044_  (.A0(\u_cpu.REG_FILE._04432_ ),
    .A1(\u_cpu.REG_FILE.rf[11][2] ),
    .S(\u_cpu.REG_FILE._04925_ ),
    .X(\u_cpu.REG_FILE._04928_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10045_  (.A(\u_cpu.REG_FILE._04928_ ),
    .X(\u_cpu.REG_FILE._00386_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10046_  (.A0(\u_cpu.REG_FILE._04434_ ),
    .A1(\u_cpu.REG_FILE.rf[11][3] ),
    .S(\u_cpu.REG_FILE._04925_ ),
    .X(\u_cpu.REG_FILE._04929_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10047_  (.A(\u_cpu.REG_FILE._04929_ ),
    .X(\u_cpu.REG_FILE._00387_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10048_  (.A0(\u_cpu.REG_FILE._04436_ ),
    .A1(\u_cpu.REG_FILE.rf[11][4] ),
    .S(\u_cpu.REG_FILE._04925_ ),
    .X(\u_cpu.REG_FILE._04930_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10049_  (.A(\u_cpu.REG_FILE._04930_ ),
    .X(\u_cpu.REG_FILE._00388_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10050_  (.A0(\u_cpu.REG_FILE._04438_ ),
    .A1(\u_cpu.REG_FILE.rf[11][5] ),
    .S(\u_cpu.REG_FILE._04925_ ),
    .X(\u_cpu.REG_FILE._04931_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10051_  (.A(\u_cpu.REG_FILE._04931_ ),
    .X(\u_cpu.REG_FILE._00389_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10052_  (.A0(\u_cpu.REG_FILE._04440_ ),
    .A1(\u_cpu.REG_FILE.rf[11][6] ),
    .S(\u_cpu.REG_FILE._04925_ ),
    .X(\u_cpu.REG_FILE._04932_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10053_  (.A(\u_cpu.REG_FILE._04932_ ),
    .X(\u_cpu.REG_FILE._00390_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10054_  (.A0(\u_cpu.REG_FILE._04442_ ),
    .A1(\u_cpu.REG_FILE.rf[11][7] ),
    .S(\u_cpu.REG_FILE._04925_ ),
    .X(\u_cpu.REG_FILE._04933_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10055_  (.A(\u_cpu.REG_FILE._04933_ ),
    .X(\u_cpu.REG_FILE._00391_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10056_  (.A0(\u_cpu.REG_FILE._04444_ ),
    .A1(\u_cpu.REG_FILE.rf[11][8] ),
    .S(\u_cpu.REG_FILE._04925_ ),
    .X(\u_cpu.REG_FILE._04934_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10057_  (.A(\u_cpu.REG_FILE._04934_ ),
    .X(\u_cpu.REG_FILE._00392_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10058_  (.A0(\u_cpu.REG_FILE._04446_ ),
    .A1(\u_cpu.REG_FILE.rf[11][9] ),
    .S(\u_cpu.REG_FILE._04925_ ),
    .X(\u_cpu.REG_FILE._04935_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10059_  (.A(\u_cpu.REG_FILE._04935_ ),
    .X(\u_cpu.REG_FILE._00393_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10060_  (.A(\u_cpu.REG_FILE._04924_ ),
    .X(\u_cpu.REG_FILE._04936_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10061_  (.A0(\u_cpu.REG_FILE._04448_ ),
    .A1(\u_cpu.REG_FILE.rf[11][10] ),
    .S(\u_cpu.REG_FILE._04936_ ),
    .X(\u_cpu.REG_FILE._04937_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10062_  (.A(\u_cpu.REG_FILE._04937_ ),
    .X(\u_cpu.REG_FILE._00394_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10063_  (.A0(\u_cpu.REG_FILE._04451_ ),
    .A1(\u_cpu.REG_FILE.rf[11][11] ),
    .S(\u_cpu.REG_FILE._04936_ ),
    .X(\u_cpu.REG_FILE._04938_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10064_  (.A(\u_cpu.REG_FILE._04938_ ),
    .X(\u_cpu.REG_FILE._00395_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10065_  (.A0(\u_cpu.REG_FILE._04453_ ),
    .A1(\u_cpu.REG_FILE.rf[11][12] ),
    .S(\u_cpu.REG_FILE._04936_ ),
    .X(\u_cpu.REG_FILE._04939_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10066_  (.A(\u_cpu.REG_FILE._04939_ ),
    .X(\u_cpu.REG_FILE._00396_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10067_  (.A0(\u_cpu.REG_FILE._04455_ ),
    .A1(\u_cpu.REG_FILE.rf[11][13] ),
    .S(\u_cpu.REG_FILE._04936_ ),
    .X(\u_cpu.REG_FILE._04940_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10068_  (.A(\u_cpu.REG_FILE._04940_ ),
    .X(\u_cpu.REG_FILE._00397_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10069_  (.A0(\u_cpu.REG_FILE._04457_ ),
    .A1(\u_cpu.REG_FILE.rf[11][14] ),
    .S(\u_cpu.REG_FILE._04936_ ),
    .X(\u_cpu.REG_FILE._04941_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10070_  (.A(\u_cpu.REG_FILE._04941_ ),
    .X(\u_cpu.REG_FILE._00398_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10071_  (.A0(\u_cpu.REG_FILE._04459_ ),
    .A1(\u_cpu.REG_FILE.rf[11][15] ),
    .S(\u_cpu.REG_FILE._04936_ ),
    .X(\u_cpu.REG_FILE._04942_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10072_  (.A(\u_cpu.REG_FILE._04942_ ),
    .X(\u_cpu.REG_FILE._00399_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10073_  (.A0(\u_cpu.REG_FILE._04461_ ),
    .A1(\u_cpu.REG_FILE.rf[11][16] ),
    .S(\u_cpu.REG_FILE._04936_ ),
    .X(\u_cpu.REG_FILE._04943_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10074_  (.A(\u_cpu.REG_FILE._04943_ ),
    .X(\u_cpu.REG_FILE._00400_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10075_  (.A0(\u_cpu.REG_FILE._04463_ ),
    .A1(\u_cpu.REG_FILE.rf[11][17] ),
    .S(\u_cpu.REG_FILE._04936_ ),
    .X(\u_cpu.REG_FILE._04944_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10076_  (.A(\u_cpu.REG_FILE._04944_ ),
    .X(\u_cpu.REG_FILE._00401_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10077_  (.A0(\u_cpu.REG_FILE._04465_ ),
    .A1(\u_cpu.REG_FILE.rf[11][18] ),
    .S(\u_cpu.REG_FILE._04936_ ),
    .X(\u_cpu.REG_FILE._04945_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10078_  (.A(\u_cpu.REG_FILE._04945_ ),
    .X(\u_cpu.REG_FILE._00402_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10079_  (.A0(\u_cpu.REG_FILE._04467_ ),
    .A1(\u_cpu.REG_FILE.rf[11][19] ),
    .S(\u_cpu.REG_FILE._04936_ ),
    .X(\u_cpu.REG_FILE._04946_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10080_  (.A(\u_cpu.REG_FILE._04946_ ),
    .X(\u_cpu.REG_FILE._00403_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10081_  (.A(\u_cpu.REG_FILE._04924_ ),
    .X(\u_cpu.REG_FILE._04947_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10082_  (.A0(\u_cpu.REG_FILE._04469_ ),
    .A1(\u_cpu.REG_FILE.rf[11][20] ),
    .S(\u_cpu.REG_FILE._04947_ ),
    .X(\u_cpu.REG_FILE._04948_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10083_  (.A(\u_cpu.REG_FILE._04948_ ),
    .X(\u_cpu.REG_FILE._00404_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10084_  (.A0(\u_cpu.REG_FILE._04472_ ),
    .A1(\u_cpu.REG_FILE.rf[11][21] ),
    .S(\u_cpu.REG_FILE._04947_ ),
    .X(\u_cpu.REG_FILE._04949_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10085_  (.A(\u_cpu.REG_FILE._04949_ ),
    .X(\u_cpu.REG_FILE._00405_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10086_  (.A0(\u_cpu.REG_FILE._04474_ ),
    .A1(\u_cpu.REG_FILE.rf[11][22] ),
    .S(\u_cpu.REG_FILE._04947_ ),
    .X(\u_cpu.REG_FILE._04950_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10087_  (.A(\u_cpu.REG_FILE._04950_ ),
    .X(\u_cpu.REG_FILE._00406_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10088_  (.A0(\u_cpu.REG_FILE._04476_ ),
    .A1(\u_cpu.REG_FILE.rf[11][23] ),
    .S(\u_cpu.REG_FILE._04947_ ),
    .X(\u_cpu.REG_FILE._04951_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10089_  (.A(\u_cpu.REG_FILE._04951_ ),
    .X(\u_cpu.REG_FILE._00407_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10090_  (.A0(\u_cpu.REG_FILE._04478_ ),
    .A1(\u_cpu.REG_FILE.rf[11][24] ),
    .S(\u_cpu.REG_FILE._04947_ ),
    .X(\u_cpu.REG_FILE._04952_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10091_  (.A(\u_cpu.REG_FILE._04952_ ),
    .X(\u_cpu.REG_FILE._00408_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10092_  (.A0(\u_cpu.REG_FILE._04480_ ),
    .A1(\u_cpu.REG_FILE.rf[11][25] ),
    .S(\u_cpu.REG_FILE._04947_ ),
    .X(\u_cpu.REG_FILE._04953_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10093_  (.A(\u_cpu.REG_FILE._04953_ ),
    .X(\u_cpu.REG_FILE._00409_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10094_  (.A0(\u_cpu.REG_FILE._04482_ ),
    .A1(\u_cpu.REG_FILE.rf[11][26] ),
    .S(\u_cpu.REG_FILE._04947_ ),
    .X(\u_cpu.REG_FILE._04954_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10095_  (.A(\u_cpu.REG_FILE._04954_ ),
    .X(\u_cpu.REG_FILE._00410_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10096_  (.A0(\u_cpu.REG_FILE._04484_ ),
    .A1(\u_cpu.REG_FILE.rf[11][27] ),
    .S(\u_cpu.REG_FILE._04947_ ),
    .X(\u_cpu.REG_FILE._04955_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10097_  (.A(\u_cpu.REG_FILE._04955_ ),
    .X(\u_cpu.REG_FILE._00411_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10098_  (.A0(\u_cpu.REG_FILE._04486_ ),
    .A1(\u_cpu.REG_FILE.rf[11][28] ),
    .S(\u_cpu.REG_FILE._04947_ ),
    .X(\u_cpu.REG_FILE._04956_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10099_  (.A(\u_cpu.REG_FILE._04956_ ),
    .X(\u_cpu.REG_FILE._00412_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10100_  (.A0(\u_cpu.REG_FILE._04488_ ),
    .A1(\u_cpu.REG_FILE.rf[11][29] ),
    .S(\u_cpu.REG_FILE._04947_ ),
    .X(\u_cpu.REG_FILE._04957_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10101_  (.A(\u_cpu.REG_FILE._04957_ ),
    .X(\u_cpu.REG_FILE._00413_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10102_  (.A0(\u_cpu.REG_FILE._04490_ ),
    .A1(\u_cpu.REG_FILE.rf[11][30] ),
    .S(\u_cpu.REG_FILE._04924_ ),
    .X(\u_cpu.REG_FILE._04958_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10103_  (.A(\u_cpu.REG_FILE._04958_ ),
    .X(\u_cpu.REG_FILE._00414_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10104_  (.A0(\u_cpu.REG_FILE._04492_ ),
    .A1(\u_cpu.REG_FILE.rf[11][31] ),
    .S(\u_cpu.REG_FILE._04924_ ),
    .X(\u_cpu.REG_FILE._04959_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10105_  (.A(\u_cpu.REG_FILE._04959_ ),
    .X(\u_cpu.REG_FILE._00415_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu.REG_FILE._10106_  (.A_N(\u_cpu.REG_FILE._04496_ ),
    .B(\u_cpu.REG_FILE._04422_ ),
    .C(\u_cpu.REG_FILE._04494_ ),
    .D(\u_cpu.REG_FILE._04643_ ),
    .Y(\u_cpu.REG_FILE._04960_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10107_  (.A(\u_cpu.REG_FILE._04960_ ),
    .X(\u_cpu.REG_FILE._04961_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10108_  (.A0(\u_cpu.REG_FILE._04420_ ),
    .A1(\u_cpu.REG_FILE.rf[12][0] ),
    .S(\u_cpu.REG_FILE._04961_ ),
    .X(\u_cpu.REG_FILE._04962_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10109_  (.A(\u_cpu.REG_FILE._04962_ ),
    .X(\u_cpu.REG_FILE._00416_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10110_  (.A0(\u_cpu.REG_FILE._04430_ ),
    .A1(\u_cpu.REG_FILE.rf[12][1] ),
    .S(\u_cpu.REG_FILE._04961_ ),
    .X(\u_cpu.REG_FILE._04963_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10111_  (.A(\u_cpu.REG_FILE._04963_ ),
    .X(\u_cpu.REG_FILE._00417_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10112_  (.A0(\u_cpu.REG_FILE._04432_ ),
    .A1(\u_cpu.REG_FILE.rf[12][2] ),
    .S(\u_cpu.REG_FILE._04961_ ),
    .X(\u_cpu.REG_FILE._04964_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10113_  (.A(\u_cpu.REG_FILE._04964_ ),
    .X(\u_cpu.REG_FILE._00418_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10114_  (.A0(\u_cpu.REG_FILE._04434_ ),
    .A1(\u_cpu.REG_FILE.rf[12][3] ),
    .S(\u_cpu.REG_FILE._04961_ ),
    .X(\u_cpu.REG_FILE._04965_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10115_  (.A(\u_cpu.REG_FILE._04965_ ),
    .X(\u_cpu.REG_FILE._00419_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10116_  (.A0(\u_cpu.REG_FILE._04436_ ),
    .A1(\u_cpu.REG_FILE.rf[12][4] ),
    .S(\u_cpu.REG_FILE._04961_ ),
    .X(\u_cpu.REG_FILE._04966_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10117_  (.A(\u_cpu.REG_FILE._04966_ ),
    .X(\u_cpu.REG_FILE._00420_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10118_  (.A0(\u_cpu.REG_FILE._04438_ ),
    .A1(\u_cpu.REG_FILE.rf[12][5] ),
    .S(\u_cpu.REG_FILE._04961_ ),
    .X(\u_cpu.REG_FILE._04967_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10119_  (.A(\u_cpu.REG_FILE._04967_ ),
    .X(\u_cpu.REG_FILE._00421_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10120_  (.A0(\u_cpu.REG_FILE._04440_ ),
    .A1(\u_cpu.REG_FILE.rf[12][6] ),
    .S(\u_cpu.REG_FILE._04961_ ),
    .X(\u_cpu.REG_FILE._04968_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10121_  (.A(\u_cpu.REG_FILE._04968_ ),
    .X(\u_cpu.REG_FILE._00422_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10122_  (.A0(\u_cpu.REG_FILE._04442_ ),
    .A1(\u_cpu.REG_FILE.rf[12][7] ),
    .S(\u_cpu.REG_FILE._04961_ ),
    .X(\u_cpu.REG_FILE._04969_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10123_  (.A(\u_cpu.REG_FILE._04969_ ),
    .X(\u_cpu.REG_FILE._00423_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10124_  (.A0(\u_cpu.REG_FILE._04444_ ),
    .A1(\u_cpu.REG_FILE.rf[12][8] ),
    .S(\u_cpu.REG_FILE._04961_ ),
    .X(\u_cpu.REG_FILE._04970_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10125_  (.A(\u_cpu.REG_FILE._04970_ ),
    .X(\u_cpu.REG_FILE._00424_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10126_  (.A0(\u_cpu.REG_FILE._04446_ ),
    .A1(\u_cpu.REG_FILE.rf[12][9] ),
    .S(\u_cpu.REG_FILE._04961_ ),
    .X(\u_cpu.REG_FILE._04971_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10127_  (.A(\u_cpu.REG_FILE._04971_ ),
    .X(\u_cpu.REG_FILE._00425_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10128_  (.A(\u_cpu.REG_FILE._04960_ ),
    .X(\u_cpu.REG_FILE._04972_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10129_  (.A0(\u_cpu.REG_FILE._04448_ ),
    .A1(\u_cpu.REG_FILE.rf[12][10] ),
    .S(\u_cpu.REG_FILE._04972_ ),
    .X(\u_cpu.REG_FILE._04973_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10130_  (.A(\u_cpu.REG_FILE._04973_ ),
    .X(\u_cpu.REG_FILE._00426_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10131_  (.A0(\u_cpu.REG_FILE._04451_ ),
    .A1(\u_cpu.REG_FILE.rf[12][11] ),
    .S(\u_cpu.REG_FILE._04972_ ),
    .X(\u_cpu.REG_FILE._04974_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10132_  (.A(\u_cpu.REG_FILE._04974_ ),
    .X(\u_cpu.REG_FILE._00427_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10133_  (.A0(\u_cpu.REG_FILE._04453_ ),
    .A1(\u_cpu.REG_FILE.rf[12][12] ),
    .S(\u_cpu.REG_FILE._04972_ ),
    .X(\u_cpu.REG_FILE._04975_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10134_  (.A(\u_cpu.REG_FILE._04975_ ),
    .X(\u_cpu.REG_FILE._00428_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10135_  (.A0(\u_cpu.REG_FILE._04455_ ),
    .A1(\u_cpu.REG_FILE.rf[12][13] ),
    .S(\u_cpu.REG_FILE._04972_ ),
    .X(\u_cpu.REG_FILE._04976_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10136_  (.A(\u_cpu.REG_FILE._04976_ ),
    .X(\u_cpu.REG_FILE._00429_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10137_  (.A0(\u_cpu.REG_FILE._04457_ ),
    .A1(\u_cpu.REG_FILE.rf[12][14] ),
    .S(\u_cpu.REG_FILE._04972_ ),
    .X(\u_cpu.REG_FILE._04977_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10138_  (.A(\u_cpu.REG_FILE._04977_ ),
    .X(\u_cpu.REG_FILE._00430_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10139_  (.A0(\u_cpu.REG_FILE._04459_ ),
    .A1(\u_cpu.REG_FILE.rf[12][15] ),
    .S(\u_cpu.REG_FILE._04972_ ),
    .X(\u_cpu.REG_FILE._04978_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10140_  (.A(\u_cpu.REG_FILE._04978_ ),
    .X(\u_cpu.REG_FILE._00431_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10141_  (.A0(\u_cpu.REG_FILE._04461_ ),
    .A1(\u_cpu.REG_FILE.rf[12][16] ),
    .S(\u_cpu.REG_FILE._04972_ ),
    .X(\u_cpu.REG_FILE._04979_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10142_  (.A(\u_cpu.REG_FILE._04979_ ),
    .X(\u_cpu.REG_FILE._00432_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10143_  (.A0(\u_cpu.REG_FILE._04463_ ),
    .A1(\u_cpu.REG_FILE.rf[12][17] ),
    .S(\u_cpu.REG_FILE._04972_ ),
    .X(\u_cpu.REG_FILE._04980_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10144_  (.A(\u_cpu.REG_FILE._04980_ ),
    .X(\u_cpu.REG_FILE._00433_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10145_  (.A0(\u_cpu.REG_FILE._04465_ ),
    .A1(\u_cpu.REG_FILE.rf[12][18] ),
    .S(\u_cpu.REG_FILE._04972_ ),
    .X(\u_cpu.REG_FILE._04981_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10146_  (.A(\u_cpu.REG_FILE._04981_ ),
    .X(\u_cpu.REG_FILE._00434_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10147_  (.A0(\u_cpu.REG_FILE._04467_ ),
    .A1(\u_cpu.REG_FILE.rf[12][19] ),
    .S(\u_cpu.REG_FILE._04972_ ),
    .X(\u_cpu.REG_FILE._04982_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10148_  (.A(\u_cpu.REG_FILE._04982_ ),
    .X(\u_cpu.REG_FILE._00435_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10149_  (.A(\u_cpu.REG_FILE._04960_ ),
    .X(\u_cpu.REG_FILE._04983_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10150_  (.A0(\u_cpu.REG_FILE._04469_ ),
    .A1(\u_cpu.REG_FILE.rf[12][20] ),
    .S(\u_cpu.REG_FILE._04983_ ),
    .X(\u_cpu.REG_FILE._04984_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10151_  (.A(\u_cpu.REG_FILE._04984_ ),
    .X(\u_cpu.REG_FILE._00436_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10152_  (.A0(\u_cpu.REG_FILE._04472_ ),
    .A1(\u_cpu.REG_FILE.rf[12][21] ),
    .S(\u_cpu.REG_FILE._04983_ ),
    .X(\u_cpu.REG_FILE._04985_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10153_  (.A(\u_cpu.REG_FILE._04985_ ),
    .X(\u_cpu.REG_FILE._00437_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10154_  (.A0(\u_cpu.REG_FILE._04474_ ),
    .A1(\u_cpu.REG_FILE.rf[12][22] ),
    .S(\u_cpu.REG_FILE._04983_ ),
    .X(\u_cpu.REG_FILE._04986_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10155_  (.A(\u_cpu.REG_FILE._04986_ ),
    .X(\u_cpu.REG_FILE._00438_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10156_  (.A0(\u_cpu.REG_FILE._04476_ ),
    .A1(\u_cpu.REG_FILE.rf[12][23] ),
    .S(\u_cpu.REG_FILE._04983_ ),
    .X(\u_cpu.REG_FILE._04987_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10157_  (.A(\u_cpu.REG_FILE._04987_ ),
    .X(\u_cpu.REG_FILE._00439_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10158_  (.A0(\u_cpu.REG_FILE._04478_ ),
    .A1(\u_cpu.REG_FILE.rf[12][24] ),
    .S(\u_cpu.REG_FILE._04983_ ),
    .X(\u_cpu.REG_FILE._04988_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10159_  (.A(\u_cpu.REG_FILE._04988_ ),
    .X(\u_cpu.REG_FILE._00440_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10160_  (.A0(\u_cpu.REG_FILE._04480_ ),
    .A1(\u_cpu.REG_FILE.rf[12][25] ),
    .S(\u_cpu.REG_FILE._04983_ ),
    .X(\u_cpu.REG_FILE._04989_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10161_  (.A(\u_cpu.REG_FILE._04989_ ),
    .X(\u_cpu.REG_FILE._00441_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10162_  (.A0(\u_cpu.REG_FILE._04482_ ),
    .A1(\u_cpu.REG_FILE.rf[12][26] ),
    .S(\u_cpu.REG_FILE._04983_ ),
    .X(\u_cpu.REG_FILE._04990_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10163_  (.A(\u_cpu.REG_FILE._04990_ ),
    .X(\u_cpu.REG_FILE._00442_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10164_  (.A0(\u_cpu.REG_FILE._04484_ ),
    .A1(\u_cpu.REG_FILE.rf[12][27] ),
    .S(\u_cpu.REG_FILE._04983_ ),
    .X(\u_cpu.REG_FILE._04991_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10165_  (.A(\u_cpu.REG_FILE._04991_ ),
    .X(\u_cpu.REG_FILE._00443_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10166_  (.A0(\u_cpu.REG_FILE._04486_ ),
    .A1(\u_cpu.REG_FILE.rf[12][28] ),
    .S(\u_cpu.REG_FILE._04983_ ),
    .X(\u_cpu.REG_FILE._04992_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10167_  (.A(\u_cpu.REG_FILE._04992_ ),
    .X(\u_cpu.REG_FILE._00444_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10168_  (.A0(\u_cpu.REG_FILE._04488_ ),
    .A1(\u_cpu.REG_FILE.rf[12][29] ),
    .S(\u_cpu.REG_FILE._04983_ ),
    .X(\u_cpu.REG_FILE._04993_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10169_  (.A(\u_cpu.REG_FILE._04993_ ),
    .X(\u_cpu.REG_FILE._00445_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10170_  (.A0(\u_cpu.REG_FILE._04490_ ),
    .A1(\u_cpu.REG_FILE.rf[12][30] ),
    .S(\u_cpu.REG_FILE._04960_ ),
    .X(\u_cpu.REG_FILE._04994_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10171_  (.A(\u_cpu.REG_FILE._04994_ ),
    .X(\u_cpu.REG_FILE._00446_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10172_  (.A0(\u_cpu.REG_FILE._04492_ ),
    .A1(\u_cpu.REG_FILE.rf[12][31] ),
    .S(\u_cpu.REG_FILE._04960_ ),
    .X(\u_cpu.REG_FILE._04995_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10173_  (.A(\u_cpu.REG_FILE._04995_ ),
    .X(\u_cpu.REG_FILE._00447_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.REG_FILE._10174_  (.A_N(\u_cpu.REG_FILE._04424_ ),
    .B(\u_cpu.REG_FILE.a3[3] ),
    .C(\u_cpu.REG_FILE.a3[2] ),
    .D(\u_cpu.REG_FILE._04423_ ),
    .X(\u_cpu.REG_FILE._04996_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10175_  (.A(\u_cpu.REG_FILE._04996_ ),
    .X(\u_cpu.REG_FILE._04997_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10176_  (.A(\u_cpu.REG_FILE._04997_ ),
    .X(\u_cpu.REG_FILE._04998_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10177_  (.A0(\u_cpu.REG_FILE.rf[13][0] ),
    .A1(\u_cpu.REG_FILE._04642_ ),
    .S(\u_cpu.REG_FILE._04998_ ),
    .X(\u_cpu.REG_FILE._04999_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10178_  (.A(\u_cpu.REG_FILE._04999_ ),
    .X(\u_cpu.REG_FILE._00448_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10179_  (.A0(\u_cpu.REG_FILE.rf[13][1] ),
    .A1(\u_cpu.REG_FILE._04647_ ),
    .S(\u_cpu.REG_FILE._04998_ ),
    .X(\u_cpu.REG_FILE._05000_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10180_  (.A(\u_cpu.REG_FILE._05000_ ),
    .X(\u_cpu.REG_FILE._00449_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10181_  (.A0(\u_cpu.REG_FILE.rf[13][2] ),
    .A1(\u_cpu.REG_FILE._04649_ ),
    .S(\u_cpu.REG_FILE._04998_ ),
    .X(\u_cpu.REG_FILE._05001_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10182_  (.A(\u_cpu.REG_FILE._05001_ ),
    .X(\u_cpu.REG_FILE._00450_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10183_  (.A0(\u_cpu.REG_FILE.rf[13][3] ),
    .A1(\u_cpu.REG_FILE._04651_ ),
    .S(\u_cpu.REG_FILE._04998_ ),
    .X(\u_cpu.REG_FILE._05002_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10184_  (.A(\u_cpu.REG_FILE._05002_ ),
    .X(\u_cpu.REG_FILE._00451_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10185_  (.A0(\u_cpu.REG_FILE.rf[13][4] ),
    .A1(\u_cpu.REG_FILE._04653_ ),
    .S(\u_cpu.REG_FILE._04998_ ),
    .X(\u_cpu.REG_FILE._05003_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10186_  (.A(\u_cpu.REG_FILE._05003_ ),
    .X(\u_cpu.REG_FILE._00452_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10187_  (.A0(\u_cpu.REG_FILE.rf[13][5] ),
    .A1(\u_cpu.REG_FILE._04655_ ),
    .S(\u_cpu.REG_FILE._04998_ ),
    .X(\u_cpu.REG_FILE._05004_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10188_  (.A(\u_cpu.REG_FILE._05004_ ),
    .X(\u_cpu.REG_FILE._00453_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10189_  (.A0(\u_cpu.REG_FILE.rf[13][6] ),
    .A1(\u_cpu.REG_FILE._04657_ ),
    .S(\u_cpu.REG_FILE._04998_ ),
    .X(\u_cpu.REG_FILE._05005_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10190_  (.A(\u_cpu.REG_FILE._05005_ ),
    .X(\u_cpu.REG_FILE._00454_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10191_  (.A0(\u_cpu.REG_FILE.rf[13][7] ),
    .A1(\u_cpu.REG_FILE._04659_ ),
    .S(\u_cpu.REG_FILE._04998_ ),
    .X(\u_cpu.REG_FILE._05006_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10192_  (.A(\u_cpu.REG_FILE._05006_ ),
    .X(\u_cpu.REG_FILE._00455_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10193_  (.A0(\u_cpu.REG_FILE.rf[13][8] ),
    .A1(\u_cpu.REG_FILE._04661_ ),
    .S(\u_cpu.REG_FILE._04998_ ),
    .X(\u_cpu.REG_FILE._05007_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10194_  (.A(\u_cpu.REG_FILE._05007_ ),
    .X(\u_cpu.REG_FILE._00456_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10195_  (.A0(\u_cpu.REG_FILE.rf[13][9] ),
    .A1(\u_cpu.REG_FILE._04663_ ),
    .S(\u_cpu.REG_FILE._04998_ ),
    .X(\u_cpu.REG_FILE._05008_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10196_  (.A(\u_cpu.REG_FILE._05008_ ),
    .X(\u_cpu.REG_FILE._00457_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10197_  (.A(\u_cpu.REG_FILE._04997_ ),
    .X(\u_cpu.REG_FILE._05009_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10198_  (.A0(\u_cpu.REG_FILE.rf[13][10] ),
    .A1(\u_cpu.REG_FILE._04665_ ),
    .S(\u_cpu.REG_FILE._05009_ ),
    .X(\u_cpu.REG_FILE._05010_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10199_  (.A(\u_cpu.REG_FILE._05010_ ),
    .X(\u_cpu.REG_FILE._00458_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10200_  (.A0(\u_cpu.REG_FILE.rf[13][11] ),
    .A1(\u_cpu.REG_FILE._04668_ ),
    .S(\u_cpu.REG_FILE._05009_ ),
    .X(\u_cpu.REG_FILE._05011_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10201_  (.A(\u_cpu.REG_FILE._05011_ ),
    .X(\u_cpu.REG_FILE._00459_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10202_  (.A0(\u_cpu.REG_FILE.rf[13][12] ),
    .A1(\u_cpu.REG_FILE._04670_ ),
    .S(\u_cpu.REG_FILE._05009_ ),
    .X(\u_cpu.REG_FILE._05012_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10203_  (.A(\u_cpu.REG_FILE._05012_ ),
    .X(\u_cpu.REG_FILE._00460_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10204_  (.A0(\u_cpu.REG_FILE.rf[13][13] ),
    .A1(\u_cpu.REG_FILE._04672_ ),
    .S(\u_cpu.REG_FILE._05009_ ),
    .X(\u_cpu.REG_FILE._05013_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10205_  (.A(\u_cpu.REG_FILE._05013_ ),
    .X(\u_cpu.REG_FILE._00461_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10206_  (.A0(\u_cpu.REG_FILE.rf[13][14] ),
    .A1(\u_cpu.REG_FILE._04674_ ),
    .S(\u_cpu.REG_FILE._05009_ ),
    .X(\u_cpu.REG_FILE._05014_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10207_  (.A(\u_cpu.REG_FILE._05014_ ),
    .X(\u_cpu.REG_FILE._00462_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10208_  (.A0(\u_cpu.REG_FILE.rf[13][15] ),
    .A1(\u_cpu.REG_FILE._04676_ ),
    .S(\u_cpu.REG_FILE._05009_ ),
    .X(\u_cpu.REG_FILE._05015_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10209_  (.A(\u_cpu.REG_FILE._05015_ ),
    .X(\u_cpu.REG_FILE._00463_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10210_  (.A0(\u_cpu.REG_FILE.rf[13][16] ),
    .A1(\u_cpu.REG_FILE._04678_ ),
    .S(\u_cpu.REG_FILE._05009_ ),
    .X(\u_cpu.REG_FILE._05016_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10211_  (.A(\u_cpu.REG_FILE._05016_ ),
    .X(\u_cpu.REG_FILE._00464_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10212_  (.A0(\u_cpu.REG_FILE.rf[13][17] ),
    .A1(\u_cpu.REG_FILE._04680_ ),
    .S(\u_cpu.REG_FILE._05009_ ),
    .X(\u_cpu.REG_FILE._05017_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10213_  (.A(\u_cpu.REG_FILE._05017_ ),
    .X(\u_cpu.REG_FILE._00465_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10214_  (.A0(\u_cpu.REG_FILE.rf[13][18] ),
    .A1(\u_cpu.REG_FILE._04682_ ),
    .S(\u_cpu.REG_FILE._05009_ ),
    .X(\u_cpu.REG_FILE._05018_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10215_  (.A(\u_cpu.REG_FILE._05018_ ),
    .X(\u_cpu.REG_FILE._00466_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10216_  (.A0(\u_cpu.REG_FILE.rf[13][19] ),
    .A1(\u_cpu.REG_FILE._04684_ ),
    .S(\u_cpu.REG_FILE._05009_ ),
    .X(\u_cpu.REG_FILE._05019_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10217_  (.A(\u_cpu.REG_FILE._05019_ ),
    .X(\u_cpu.REG_FILE._00467_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10218_  (.A(\u_cpu.REG_FILE._04997_ ),
    .X(\u_cpu.REG_FILE._05020_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10219_  (.A0(\u_cpu.REG_FILE.rf[13][20] ),
    .A1(\u_cpu.REG_FILE._04686_ ),
    .S(\u_cpu.REG_FILE._05020_ ),
    .X(\u_cpu.REG_FILE._05021_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10220_  (.A(\u_cpu.REG_FILE._05021_ ),
    .X(\u_cpu.REG_FILE._00468_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10221_  (.A0(\u_cpu.REG_FILE.rf[13][21] ),
    .A1(\u_cpu.REG_FILE._04689_ ),
    .S(\u_cpu.REG_FILE._05020_ ),
    .X(\u_cpu.REG_FILE._05022_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10222_  (.A(\u_cpu.REG_FILE._05022_ ),
    .X(\u_cpu.REG_FILE._00469_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10223_  (.A0(\u_cpu.REG_FILE.rf[13][22] ),
    .A1(\u_cpu.REG_FILE._04691_ ),
    .S(\u_cpu.REG_FILE._05020_ ),
    .X(\u_cpu.REG_FILE._05023_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10224_  (.A(\u_cpu.REG_FILE._05023_ ),
    .X(\u_cpu.REG_FILE._00470_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10225_  (.A0(\u_cpu.REG_FILE.rf[13][23] ),
    .A1(\u_cpu.REG_FILE._04693_ ),
    .S(\u_cpu.REG_FILE._05020_ ),
    .X(\u_cpu.REG_FILE._05024_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10226_  (.A(\u_cpu.REG_FILE._05024_ ),
    .X(\u_cpu.REG_FILE._00471_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10227_  (.A0(\u_cpu.REG_FILE.rf[13][24] ),
    .A1(\u_cpu.REG_FILE._04695_ ),
    .S(\u_cpu.REG_FILE._05020_ ),
    .X(\u_cpu.REG_FILE._05025_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10228_  (.A(\u_cpu.REG_FILE._05025_ ),
    .X(\u_cpu.REG_FILE._00472_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10229_  (.A0(\u_cpu.REG_FILE.rf[13][25] ),
    .A1(\u_cpu.REG_FILE._04697_ ),
    .S(\u_cpu.REG_FILE._05020_ ),
    .X(\u_cpu.REG_FILE._05026_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10230_  (.A(\u_cpu.REG_FILE._05026_ ),
    .X(\u_cpu.REG_FILE._00473_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10231_  (.A0(\u_cpu.REG_FILE.rf[13][26] ),
    .A1(\u_cpu.REG_FILE._04699_ ),
    .S(\u_cpu.REG_FILE._05020_ ),
    .X(\u_cpu.REG_FILE._05027_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10232_  (.A(\u_cpu.REG_FILE._05027_ ),
    .X(\u_cpu.REG_FILE._00474_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10233_  (.A0(\u_cpu.REG_FILE.rf[13][27] ),
    .A1(\u_cpu.REG_FILE._04701_ ),
    .S(\u_cpu.REG_FILE._05020_ ),
    .X(\u_cpu.REG_FILE._05028_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10234_  (.A(\u_cpu.REG_FILE._05028_ ),
    .X(\u_cpu.REG_FILE._00475_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10235_  (.A0(\u_cpu.REG_FILE.rf[13][28] ),
    .A1(\u_cpu.REG_FILE._04703_ ),
    .S(\u_cpu.REG_FILE._05020_ ),
    .X(\u_cpu.REG_FILE._05029_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10236_  (.A(\u_cpu.REG_FILE._05029_ ),
    .X(\u_cpu.REG_FILE._00476_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10237_  (.A0(\u_cpu.REG_FILE.rf[13][29] ),
    .A1(\u_cpu.REG_FILE._04705_ ),
    .S(\u_cpu.REG_FILE._05020_ ),
    .X(\u_cpu.REG_FILE._05030_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10238_  (.A(\u_cpu.REG_FILE._05030_ ),
    .X(\u_cpu.REG_FILE._00477_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10239_  (.A0(\u_cpu.REG_FILE.rf[13][30] ),
    .A1(\u_cpu.REG_FILE._04707_ ),
    .S(\u_cpu.REG_FILE._04997_ ),
    .X(\u_cpu.REG_FILE._05031_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10240_  (.A(\u_cpu.REG_FILE._05031_ ),
    .X(\u_cpu.REG_FILE._00478_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10241_  (.A0(\u_cpu.REG_FILE.rf[13][31] ),
    .A1(\u_cpu.REG_FILE._04709_ ),
    .S(\u_cpu.REG_FILE._04997_ ),
    .X(\u_cpu.REG_FILE._05032_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10242_  (.A(\u_cpu.REG_FILE._05032_ ),
    .X(\u_cpu.REG_FILE._00479_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.REG_FILE._10243_  (.A_N(\u_cpu.REG_FILE._04424_ ),
    .B(\u_cpu.REG_FILE.a3[3] ),
    .C(\u_cpu.REG_FILE.a3[2] ),
    .D(\u_cpu.REG_FILE._04747_ ),
    .X(\u_cpu.REG_FILE._05033_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10244_  (.A(\u_cpu.REG_FILE._05033_ ),
    .X(\u_cpu.REG_FILE._05034_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10245_  (.A(\u_cpu.REG_FILE._05034_ ),
    .X(\u_cpu.REG_FILE._05035_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10246_  (.A0(\u_cpu.REG_FILE.rf[14][0] ),
    .A1(\u_cpu.REG_FILE._04642_ ),
    .S(\u_cpu.REG_FILE._05035_ ),
    .X(\u_cpu.REG_FILE._05036_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10247_  (.A(\u_cpu.REG_FILE._05036_ ),
    .X(\u_cpu.REG_FILE._00480_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10248_  (.A0(\u_cpu.REG_FILE.rf[14][1] ),
    .A1(\u_cpu.REG_FILE._04647_ ),
    .S(\u_cpu.REG_FILE._05035_ ),
    .X(\u_cpu.REG_FILE._05037_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10249_  (.A(\u_cpu.REG_FILE._05037_ ),
    .X(\u_cpu.REG_FILE._00481_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10250_  (.A0(\u_cpu.REG_FILE.rf[14][2] ),
    .A1(\u_cpu.REG_FILE._04649_ ),
    .S(\u_cpu.REG_FILE._05035_ ),
    .X(\u_cpu.REG_FILE._05038_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10251_  (.A(\u_cpu.REG_FILE._05038_ ),
    .X(\u_cpu.REG_FILE._00482_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10252_  (.A0(\u_cpu.REG_FILE.rf[14][3] ),
    .A1(\u_cpu.REG_FILE._04651_ ),
    .S(\u_cpu.REG_FILE._05035_ ),
    .X(\u_cpu.REG_FILE._05039_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10253_  (.A(\u_cpu.REG_FILE._05039_ ),
    .X(\u_cpu.REG_FILE._00483_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10254_  (.A0(\u_cpu.REG_FILE.rf[14][4] ),
    .A1(\u_cpu.REG_FILE._04653_ ),
    .S(\u_cpu.REG_FILE._05035_ ),
    .X(\u_cpu.REG_FILE._05040_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10255_  (.A(\u_cpu.REG_FILE._05040_ ),
    .X(\u_cpu.REG_FILE._00484_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10256_  (.A0(\u_cpu.REG_FILE.rf[14][5] ),
    .A1(\u_cpu.REG_FILE._04655_ ),
    .S(\u_cpu.REG_FILE._05035_ ),
    .X(\u_cpu.REG_FILE._05041_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10257_  (.A(\u_cpu.REG_FILE._05041_ ),
    .X(\u_cpu.REG_FILE._00485_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10258_  (.A0(\u_cpu.REG_FILE.rf[14][6] ),
    .A1(\u_cpu.REG_FILE._04657_ ),
    .S(\u_cpu.REG_FILE._05035_ ),
    .X(\u_cpu.REG_FILE._05042_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10259_  (.A(\u_cpu.REG_FILE._05042_ ),
    .X(\u_cpu.REG_FILE._00486_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10260_  (.A0(\u_cpu.REG_FILE.rf[14][7] ),
    .A1(\u_cpu.REG_FILE._04659_ ),
    .S(\u_cpu.REG_FILE._05035_ ),
    .X(\u_cpu.REG_FILE._05043_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10261_  (.A(\u_cpu.REG_FILE._05043_ ),
    .X(\u_cpu.REG_FILE._00487_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10262_  (.A0(\u_cpu.REG_FILE.rf[14][8] ),
    .A1(\u_cpu.REG_FILE._04661_ ),
    .S(\u_cpu.REG_FILE._05035_ ),
    .X(\u_cpu.REG_FILE._05044_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10263_  (.A(\u_cpu.REG_FILE._05044_ ),
    .X(\u_cpu.REG_FILE._00488_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10264_  (.A0(\u_cpu.REG_FILE.rf[14][9] ),
    .A1(\u_cpu.REG_FILE._04663_ ),
    .S(\u_cpu.REG_FILE._05035_ ),
    .X(\u_cpu.REG_FILE._05045_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10265_  (.A(\u_cpu.REG_FILE._05045_ ),
    .X(\u_cpu.REG_FILE._00489_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10266_  (.A(\u_cpu.REG_FILE._05034_ ),
    .X(\u_cpu.REG_FILE._05046_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10267_  (.A0(\u_cpu.REG_FILE.rf[14][10] ),
    .A1(\u_cpu.REG_FILE._04665_ ),
    .S(\u_cpu.REG_FILE._05046_ ),
    .X(\u_cpu.REG_FILE._05047_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10268_  (.A(\u_cpu.REG_FILE._05047_ ),
    .X(\u_cpu.REG_FILE._00490_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10269_  (.A0(\u_cpu.REG_FILE.rf[14][11] ),
    .A1(\u_cpu.REG_FILE._04668_ ),
    .S(\u_cpu.REG_FILE._05046_ ),
    .X(\u_cpu.REG_FILE._05048_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10270_  (.A(\u_cpu.REG_FILE._05048_ ),
    .X(\u_cpu.REG_FILE._00491_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10271_  (.A0(\u_cpu.REG_FILE.rf[14][12] ),
    .A1(\u_cpu.REG_FILE._04670_ ),
    .S(\u_cpu.REG_FILE._05046_ ),
    .X(\u_cpu.REG_FILE._05049_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10272_  (.A(\u_cpu.REG_FILE._05049_ ),
    .X(\u_cpu.REG_FILE._00492_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10273_  (.A0(\u_cpu.REG_FILE.rf[14][13] ),
    .A1(\u_cpu.REG_FILE._04672_ ),
    .S(\u_cpu.REG_FILE._05046_ ),
    .X(\u_cpu.REG_FILE._05050_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10274_  (.A(\u_cpu.REG_FILE._05050_ ),
    .X(\u_cpu.REG_FILE._00493_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10275_  (.A0(\u_cpu.REG_FILE.rf[14][14] ),
    .A1(\u_cpu.REG_FILE._04674_ ),
    .S(\u_cpu.REG_FILE._05046_ ),
    .X(\u_cpu.REG_FILE._05051_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10276_  (.A(\u_cpu.REG_FILE._05051_ ),
    .X(\u_cpu.REG_FILE._00494_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10277_  (.A0(\u_cpu.REG_FILE.rf[14][15] ),
    .A1(\u_cpu.REG_FILE._04676_ ),
    .S(\u_cpu.REG_FILE._05046_ ),
    .X(\u_cpu.REG_FILE._05052_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10278_  (.A(\u_cpu.REG_FILE._05052_ ),
    .X(\u_cpu.REG_FILE._00495_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10279_  (.A0(\u_cpu.REG_FILE.rf[14][16] ),
    .A1(\u_cpu.REG_FILE._04678_ ),
    .S(\u_cpu.REG_FILE._05046_ ),
    .X(\u_cpu.REG_FILE._05053_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10280_  (.A(\u_cpu.REG_FILE._05053_ ),
    .X(\u_cpu.REG_FILE._00496_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10281_  (.A0(\u_cpu.REG_FILE.rf[14][17] ),
    .A1(\u_cpu.REG_FILE._04680_ ),
    .S(\u_cpu.REG_FILE._05046_ ),
    .X(\u_cpu.REG_FILE._05054_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10282_  (.A(\u_cpu.REG_FILE._05054_ ),
    .X(\u_cpu.REG_FILE._00497_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10283_  (.A0(\u_cpu.REG_FILE.rf[14][18] ),
    .A1(\u_cpu.REG_FILE._04682_ ),
    .S(\u_cpu.REG_FILE._05046_ ),
    .X(\u_cpu.REG_FILE._05055_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10284_  (.A(\u_cpu.REG_FILE._05055_ ),
    .X(\u_cpu.REG_FILE._00498_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10285_  (.A0(\u_cpu.REG_FILE.rf[14][19] ),
    .A1(\u_cpu.REG_FILE._04684_ ),
    .S(\u_cpu.REG_FILE._05046_ ),
    .X(\u_cpu.REG_FILE._05056_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10286_  (.A(\u_cpu.REG_FILE._05056_ ),
    .X(\u_cpu.REG_FILE._00499_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10287_  (.A(\u_cpu.REG_FILE._05034_ ),
    .X(\u_cpu.REG_FILE._05057_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10288_  (.A0(\u_cpu.REG_FILE.rf[14][20] ),
    .A1(\u_cpu.REG_FILE._04686_ ),
    .S(\u_cpu.REG_FILE._05057_ ),
    .X(\u_cpu.REG_FILE._05058_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10289_  (.A(\u_cpu.REG_FILE._05058_ ),
    .X(\u_cpu.REG_FILE._00500_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10290_  (.A0(\u_cpu.REG_FILE.rf[14][21] ),
    .A1(\u_cpu.REG_FILE._04689_ ),
    .S(\u_cpu.REG_FILE._05057_ ),
    .X(\u_cpu.REG_FILE._05059_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10291_  (.A(\u_cpu.REG_FILE._05059_ ),
    .X(\u_cpu.REG_FILE._00501_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10292_  (.A0(\u_cpu.REG_FILE.rf[14][22] ),
    .A1(\u_cpu.REG_FILE._04691_ ),
    .S(\u_cpu.REG_FILE._05057_ ),
    .X(\u_cpu.REG_FILE._05060_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10293_  (.A(\u_cpu.REG_FILE._05060_ ),
    .X(\u_cpu.REG_FILE._00502_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10294_  (.A0(\u_cpu.REG_FILE.rf[14][23] ),
    .A1(\u_cpu.REG_FILE._04693_ ),
    .S(\u_cpu.REG_FILE._05057_ ),
    .X(\u_cpu.REG_FILE._05061_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10295_  (.A(\u_cpu.REG_FILE._05061_ ),
    .X(\u_cpu.REG_FILE._00503_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10296_  (.A0(\u_cpu.REG_FILE.rf[14][24] ),
    .A1(\u_cpu.REG_FILE._04695_ ),
    .S(\u_cpu.REG_FILE._05057_ ),
    .X(\u_cpu.REG_FILE._05062_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10297_  (.A(\u_cpu.REG_FILE._05062_ ),
    .X(\u_cpu.REG_FILE._00504_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10298_  (.A0(\u_cpu.REG_FILE.rf[14][25] ),
    .A1(\u_cpu.REG_FILE._04697_ ),
    .S(\u_cpu.REG_FILE._05057_ ),
    .X(\u_cpu.REG_FILE._05063_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10299_  (.A(\u_cpu.REG_FILE._05063_ ),
    .X(\u_cpu.REG_FILE._00505_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10300_  (.A0(\u_cpu.REG_FILE.rf[14][26] ),
    .A1(\u_cpu.REG_FILE._04699_ ),
    .S(\u_cpu.REG_FILE._05057_ ),
    .X(\u_cpu.REG_FILE._05064_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10301_  (.A(\u_cpu.REG_FILE._05064_ ),
    .X(\u_cpu.REG_FILE._00506_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10302_  (.A0(\u_cpu.REG_FILE.rf[14][27] ),
    .A1(\u_cpu.REG_FILE._04701_ ),
    .S(\u_cpu.REG_FILE._05057_ ),
    .X(\u_cpu.REG_FILE._05065_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10303_  (.A(\u_cpu.REG_FILE._05065_ ),
    .X(\u_cpu.REG_FILE._00507_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10304_  (.A0(\u_cpu.REG_FILE.rf[14][28] ),
    .A1(\u_cpu.REG_FILE._04703_ ),
    .S(\u_cpu.REG_FILE._05057_ ),
    .X(\u_cpu.REG_FILE._05066_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10305_  (.A(\u_cpu.REG_FILE._05066_ ),
    .X(\u_cpu.REG_FILE._00508_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10306_  (.A0(\u_cpu.REG_FILE.rf[14][29] ),
    .A1(\u_cpu.REG_FILE._04705_ ),
    .S(\u_cpu.REG_FILE._05057_ ),
    .X(\u_cpu.REG_FILE._05067_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10307_  (.A(\u_cpu.REG_FILE._05067_ ),
    .X(\u_cpu.REG_FILE._00509_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10308_  (.A0(\u_cpu.REG_FILE.rf[14][30] ),
    .A1(\u_cpu.REG_FILE._04707_ ),
    .S(\u_cpu.REG_FILE._05034_ ),
    .X(\u_cpu.REG_FILE._05068_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10309_  (.A(\u_cpu.REG_FILE._05068_ ),
    .X(\u_cpu.REG_FILE._00510_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10310_  (.A0(\u_cpu.REG_FILE.rf[14][31] ),
    .A1(\u_cpu.REG_FILE._04709_ ),
    .S(\u_cpu.REG_FILE._05034_ ),
    .X(\u_cpu.REG_FILE._05069_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10311_  (.A(\u_cpu.REG_FILE._05069_ ),
    .X(\u_cpu.REG_FILE._00511_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.REG_FILE._10312_  (.A_N(\u_cpu.REG_FILE._04424_ ),
    .B(\u_cpu.REG_FILE.a3[3] ),
    .C(\u_cpu.REG_FILE.a3[2] ),
    .D(\u_cpu.REG_FILE._04495_ ),
    .X(\u_cpu.REG_FILE._05070_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10313_  (.A(\u_cpu.REG_FILE._05070_ ),
    .X(\u_cpu.REG_FILE._05071_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10314_  (.A(\u_cpu.REG_FILE._05071_ ),
    .X(\u_cpu.REG_FILE._05072_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10315_  (.A0(\u_cpu.REG_FILE.rf[15][0] ),
    .A1(\u_cpu.REG_FILE._04642_ ),
    .S(\u_cpu.REG_FILE._05072_ ),
    .X(\u_cpu.REG_FILE._05073_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10316_  (.A(\u_cpu.REG_FILE._05073_ ),
    .X(\u_cpu.REG_FILE._00512_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10317_  (.A0(\u_cpu.REG_FILE.rf[15][1] ),
    .A1(\u_cpu.REG_FILE._04647_ ),
    .S(\u_cpu.REG_FILE._05072_ ),
    .X(\u_cpu.REG_FILE._05074_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10318_  (.A(\u_cpu.REG_FILE._05074_ ),
    .X(\u_cpu.REG_FILE._00513_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10319_  (.A0(\u_cpu.REG_FILE.rf[15][2] ),
    .A1(\u_cpu.REG_FILE._04649_ ),
    .S(\u_cpu.REG_FILE._05072_ ),
    .X(\u_cpu.REG_FILE._05075_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10320_  (.A(\u_cpu.REG_FILE._05075_ ),
    .X(\u_cpu.REG_FILE._00514_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10321_  (.A0(\u_cpu.REG_FILE.rf[15][3] ),
    .A1(\u_cpu.REG_FILE._04651_ ),
    .S(\u_cpu.REG_FILE._05072_ ),
    .X(\u_cpu.REG_FILE._05076_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10322_  (.A(\u_cpu.REG_FILE._05076_ ),
    .X(\u_cpu.REG_FILE._00515_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10323_  (.A0(\u_cpu.REG_FILE.rf[15][4] ),
    .A1(\u_cpu.REG_FILE._04653_ ),
    .S(\u_cpu.REG_FILE._05072_ ),
    .X(\u_cpu.REG_FILE._05077_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10324_  (.A(\u_cpu.REG_FILE._05077_ ),
    .X(\u_cpu.REG_FILE._00516_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10325_  (.A0(\u_cpu.REG_FILE.rf[15][5] ),
    .A1(\u_cpu.REG_FILE._04655_ ),
    .S(\u_cpu.REG_FILE._05072_ ),
    .X(\u_cpu.REG_FILE._05078_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10326_  (.A(\u_cpu.REG_FILE._05078_ ),
    .X(\u_cpu.REG_FILE._00517_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10327_  (.A0(\u_cpu.REG_FILE.rf[15][6] ),
    .A1(\u_cpu.REG_FILE._04657_ ),
    .S(\u_cpu.REG_FILE._05072_ ),
    .X(\u_cpu.REG_FILE._05079_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10328_  (.A(\u_cpu.REG_FILE._05079_ ),
    .X(\u_cpu.REG_FILE._00518_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10329_  (.A0(\u_cpu.REG_FILE.rf[15][7] ),
    .A1(\u_cpu.REG_FILE._04659_ ),
    .S(\u_cpu.REG_FILE._05072_ ),
    .X(\u_cpu.REG_FILE._05080_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10330_  (.A(\u_cpu.REG_FILE._05080_ ),
    .X(\u_cpu.REG_FILE._00519_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10331_  (.A0(\u_cpu.REG_FILE.rf[15][8] ),
    .A1(\u_cpu.REG_FILE._04661_ ),
    .S(\u_cpu.REG_FILE._05072_ ),
    .X(\u_cpu.REG_FILE._05081_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10332_  (.A(\u_cpu.REG_FILE._05081_ ),
    .X(\u_cpu.REG_FILE._00520_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10333_  (.A0(\u_cpu.REG_FILE.rf[15][9] ),
    .A1(\u_cpu.REG_FILE._04663_ ),
    .S(\u_cpu.REG_FILE._05072_ ),
    .X(\u_cpu.REG_FILE._05082_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10334_  (.A(\u_cpu.REG_FILE._05082_ ),
    .X(\u_cpu.REG_FILE._00521_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10335_  (.A(\u_cpu.REG_FILE._05071_ ),
    .X(\u_cpu.REG_FILE._05083_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10336_  (.A0(\u_cpu.REG_FILE.rf[15][10] ),
    .A1(\u_cpu.REG_FILE._04665_ ),
    .S(\u_cpu.REG_FILE._05083_ ),
    .X(\u_cpu.REG_FILE._05084_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10337_  (.A(\u_cpu.REG_FILE._05084_ ),
    .X(\u_cpu.REG_FILE._00522_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10338_  (.A0(\u_cpu.REG_FILE.rf[15][11] ),
    .A1(\u_cpu.REG_FILE._04668_ ),
    .S(\u_cpu.REG_FILE._05083_ ),
    .X(\u_cpu.REG_FILE._05085_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10339_  (.A(\u_cpu.REG_FILE._05085_ ),
    .X(\u_cpu.REG_FILE._00523_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10340_  (.A0(\u_cpu.REG_FILE.rf[15][12] ),
    .A1(\u_cpu.REG_FILE._04670_ ),
    .S(\u_cpu.REG_FILE._05083_ ),
    .X(\u_cpu.REG_FILE._05086_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10341_  (.A(\u_cpu.REG_FILE._05086_ ),
    .X(\u_cpu.REG_FILE._00524_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10342_  (.A0(\u_cpu.REG_FILE.rf[15][13] ),
    .A1(\u_cpu.REG_FILE._04672_ ),
    .S(\u_cpu.REG_FILE._05083_ ),
    .X(\u_cpu.REG_FILE._05087_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10343_  (.A(\u_cpu.REG_FILE._05087_ ),
    .X(\u_cpu.REG_FILE._00525_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10344_  (.A0(\u_cpu.REG_FILE.rf[15][14] ),
    .A1(\u_cpu.REG_FILE._04674_ ),
    .S(\u_cpu.REG_FILE._05083_ ),
    .X(\u_cpu.REG_FILE._05088_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10345_  (.A(\u_cpu.REG_FILE._05088_ ),
    .X(\u_cpu.REG_FILE._00526_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10346_  (.A0(\u_cpu.REG_FILE.rf[15][15] ),
    .A1(\u_cpu.REG_FILE._04676_ ),
    .S(\u_cpu.REG_FILE._05083_ ),
    .X(\u_cpu.REG_FILE._05089_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10347_  (.A(\u_cpu.REG_FILE._05089_ ),
    .X(\u_cpu.REG_FILE._00527_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10348_  (.A0(\u_cpu.REG_FILE.rf[15][16] ),
    .A1(\u_cpu.REG_FILE._04678_ ),
    .S(\u_cpu.REG_FILE._05083_ ),
    .X(\u_cpu.REG_FILE._05090_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10349_  (.A(\u_cpu.REG_FILE._05090_ ),
    .X(\u_cpu.REG_FILE._00528_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10350_  (.A0(\u_cpu.REG_FILE.rf[15][17] ),
    .A1(\u_cpu.REG_FILE._04680_ ),
    .S(\u_cpu.REG_FILE._05083_ ),
    .X(\u_cpu.REG_FILE._05091_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10351_  (.A(\u_cpu.REG_FILE._05091_ ),
    .X(\u_cpu.REG_FILE._00529_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10352_  (.A0(\u_cpu.REG_FILE.rf[15][18] ),
    .A1(\u_cpu.REG_FILE._04682_ ),
    .S(\u_cpu.REG_FILE._05083_ ),
    .X(\u_cpu.REG_FILE._05092_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10353_  (.A(\u_cpu.REG_FILE._05092_ ),
    .X(\u_cpu.REG_FILE._00530_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10354_  (.A0(\u_cpu.REG_FILE.rf[15][19] ),
    .A1(\u_cpu.REG_FILE._04684_ ),
    .S(\u_cpu.REG_FILE._05083_ ),
    .X(\u_cpu.REG_FILE._05093_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10355_  (.A(\u_cpu.REG_FILE._05093_ ),
    .X(\u_cpu.REG_FILE._00531_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10356_  (.A(\u_cpu.REG_FILE._05071_ ),
    .X(\u_cpu.REG_FILE._05094_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10357_  (.A0(\u_cpu.REG_FILE.rf[15][20] ),
    .A1(\u_cpu.REG_FILE._04686_ ),
    .S(\u_cpu.REG_FILE._05094_ ),
    .X(\u_cpu.REG_FILE._05095_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10358_  (.A(\u_cpu.REG_FILE._05095_ ),
    .X(\u_cpu.REG_FILE._00532_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10359_  (.A0(\u_cpu.REG_FILE.rf[15][21] ),
    .A1(\u_cpu.REG_FILE._04689_ ),
    .S(\u_cpu.REG_FILE._05094_ ),
    .X(\u_cpu.REG_FILE._05096_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10360_  (.A(\u_cpu.REG_FILE._05096_ ),
    .X(\u_cpu.REG_FILE._00533_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10361_  (.A0(\u_cpu.REG_FILE.rf[15][22] ),
    .A1(\u_cpu.REG_FILE._04691_ ),
    .S(\u_cpu.REG_FILE._05094_ ),
    .X(\u_cpu.REG_FILE._05097_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10362_  (.A(\u_cpu.REG_FILE._05097_ ),
    .X(\u_cpu.REG_FILE._00534_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10363_  (.A0(\u_cpu.REG_FILE.rf[15][23] ),
    .A1(\u_cpu.REG_FILE._04693_ ),
    .S(\u_cpu.REG_FILE._05094_ ),
    .X(\u_cpu.REG_FILE._05098_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10364_  (.A(\u_cpu.REG_FILE._05098_ ),
    .X(\u_cpu.REG_FILE._00535_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10365_  (.A0(\u_cpu.REG_FILE.rf[15][24] ),
    .A1(\u_cpu.REG_FILE._04695_ ),
    .S(\u_cpu.REG_FILE._05094_ ),
    .X(\u_cpu.REG_FILE._05099_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10366_  (.A(\u_cpu.REG_FILE._05099_ ),
    .X(\u_cpu.REG_FILE._00536_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10367_  (.A0(\u_cpu.REG_FILE.rf[15][25] ),
    .A1(\u_cpu.REG_FILE._04697_ ),
    .S(\u_cpu.REG_FILE._05094_ ),
    .X(\u_cpu.REG_FILE._05100_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10368_  (.A(\u_cpu.REG_FILE._05100_ ),
    .X(\u_cpu.REG_FILE._00537_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10369_  (.A0(\u_cpu.REG_FILE.rf[15][26] ),
    .A1(\u_cpu.REG_FILE._04699_ ),
    .S(\u_cpu.REG_FILE._05094_ ),
    .X(\u_cpu.REG_FILE._05101_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10370_  (.A(\u_cpu.REG_FILE._05101_ ),
    .X(\u_cpu.REG_FILE._00538_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10371_  (.A0(\u_cpu.REG_FILE.rf[15][27] ),
    .A1(\u_cpu.REG_FILE._04701_ ),
    .S(\u_cpu.REG_FILE._05094_ ),
    .X(\u_cpu.REG_FILE._05102_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10372_  (.A(\u_cpu.REG_FILE._05102_ ),
    .X(\u_cpu.REG_FILE._00539_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10373_  (.A0(\u_cpu.REG_FILE.rf[15][28] ),
    .A1(\u_cpu.REG_FILE._04703_ ),
    .S(\u_cpu.REG_FILE._05094_ ),
    .X(\u_cpu.REG_FILE._05103_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10374_  (.A(\u_cpu.REG_FILE._05103_ ),
    .X(\u_cpu.REG_FILE._00540_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10375_  (.A0(\u_cpu.REG_FILE.rf[15][29] ),
    .A1(\u_cpu.REG_FILE._04705_ ),
    .S(\u_cpu.REG_FILE._05094_ ),
    .X(\u_cpu.REG_FILE._05104_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10376_  (.A(\u_cpu.REG_FILE._05104_ ),
    .X(\u_cpu.REG_FILE._00541_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10377_  (.A0(\u_cpu.REG_FILE.rf[15][30] ),
    .A1(\u_cpu.REG_FILE._04707_ ),
    .S(\u_cpu.REG_FILE._05071_ ),
    .X(\u_cpu.REG_FILE._05105_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10378_  (.A(\u_cpu.REG_FILE._05105_ ),
    .X(\u_cpu.REG_FILE._00542_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10379_  (.A0(\u_cpu.REG_FILE.rf[15][31] ),
    .A1(\u_cpu.REG_FILE._04709_ ),
    .S(\u_cpu.REG_FILE._05071_ ),
    .X(\u_cpu.REG_FILE._05106_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10380_  (.A(\u_cpu.REG_FILE._05106_ ),
    .X(\u_cpu.REG_FILE._00543_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu.REG_FILE._10381_  (.A(\u_cpu.REG_FILE._04421_ ),
    .B(\u_cpu.REG_FILE._04425_ ),
    .Y(\u_cpu.REG_FILE._05107_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.REG_FILE._10382_  (.A(\u_cpu.REG_FILE._04496_ ),
    .B(\u_cpu.REG_FILE._05107_ ),
    .C(\u_cpu.REG_FILE._04643_ ),
    .X(\u_cpu.REG_FILE._05108_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10383_  (.A(\u_cpu.REG_FILE._05108_ ),
    .X(\u_cpu.REG_FILE._05109_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10384_  (.A0(\u_cpu.REG_FILE.rf[16][0] ),
    .A1(\u_cpu.REG_FILE._04642_ ),
    .S(\u_cpu.REG_FILE._05109_ ),
    .X(\u_cpu.REG_FILE._05110_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10385_  (.A(\u_cpu.REG_FILE._05110_ ),
    .X(\u_cpu.REG_FILE._00544_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10386_  (.A0(\u_cpu.REG_FILE.rf[16][1] ),
    .A1(\u_cpu.REG_FILE._04647_ ),
    .S(\u_cpu.REG_FILE._05109_ ),
    .X(\u_cpu.REG_FILE._05111_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10387_  (.A(\u_cpu.REG_FILE._05111_ ),
    .X(\u_cpu.REG_FILE._00545_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10388_  (.A0(\u_cpu.REG_FILE.rf[16][2] ),
    .A1(\u_cpu.REG_FILE._04649_ ),
    .S(\u_cpu.REG_FILE._05109_ ),
    .X(\u_cpu.REG_FILE._05112_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10389_  (.A(\u_cpu.REG_FILE._05112_ ),
    .X(\u_cpu.REG_FILE._00546_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10390_  (.A0(\u_cpu.REG_FILE.rf[16][3] ),
    .A1(\u_cpu.REG_FILE._04651_ ),
    .S(\u_cpu.REG_FILE._05109_ ),
    .X(\u_cpu.REG_FILE._05113_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10391_  (.A(\u_cpu.REG_FILE._05113_ ),
    .X(\u_cpu.REG_FILE._00547_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10392_  (.A0(\u_cpu.REG_FILE.rf[16][4] ),
    .A1(\u_cpu.REG_FILE._04653_ ),
    .S(\u_cpu.REG_FILE._05109_ ),
    .X(\u_cpu.REG_FILE._05114_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10393_  (.A(\u_cpu.REG_FILE._05114_ ),
    .X(\u_cpu.REG_FILE._00548_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10394_  (.A0(\u_cpu.REG_FILE.rf[16][5] ),
    .A1(\u_cpu.REG_FILE._04655_ ),
    .S(\u_cpu.REG_FILE._05109_ ),
    .X(\u_cpu.REG_FILE._05115_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10395_  (.A(\u_cpu.REG_FILE._05115_ ),
    .X(\u_cpu.REG_FILE._00549_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10396_  (.A0(\u_cpu.REG_FILE.rf[16][6] ),
    .A1(\u_cpu.REG_FILE._04657_ ),
    .S(\u_cpu.REG_FILE._05109_ ),
    .X(\u_cpu.REG_FILE._05116_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10397_  (.A(\u_cpu.REG_FILE._05116_ ),
    .X(\u_cpu.REG_FILE._00550_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10398_  (.A0(\u_cpu.REG_FILE.rf[16][7] ),
    .A1(\u_cpu.REG_FILE._04659_ ),
    .S(\u_cpu.REG_FILE._05109_ ),
    .X(\u_cpu.REG_FILE._05117_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10399_  (.A(\u_cpu.REG_FILE._05117_ ),
    .X(\u_cpu.REG_FILE._00551_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10400_  (.A0(\u_cpu.REG_FILE.rf[16][8] ),
    .A1(\u_cpu.REG_FILE._04661_ ),
    .S(\u_cpu.REG_FILE._05109_ ),
    .X(\u_cpu.REG_FILE._05118_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10401_  (.A(\u_cpu.REG_FILE._05118_ ),
    .X(\u_cpu.REG_FILE._00552_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10402_  (.A0(\u_cpu.REG_FILE.rf[16][9] ),
    .A1(\u_cpu.REG_FILE._04663_ ),
    .S(\u_cpu.REG_FILE._05109_ ),
    .X(\u_cpu.REG_FILE._05119_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10403_  (.A(\u_cpu.REG_FILE._05119_ ),
    .X(\u_cpu.REG_FILE._00553_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10404_  (.A(\u_cpu.REG_FILE._05108_ ),
    .X(\u_cpu.REG_FILE._05120_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10405_  (.A0(\u_cpu.REG_FILE.rf[16][10] ),
    .A1(\u_cpu.REG_FILE._04665_ ),
    .S(\u_cpu.REG_FILE._05120_ ),
    .X(\u_cpu.REG_FILE._05121_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10406_  (.A(\u_cpu.REG_FILE._05121_ ),
    .X(\u_cpu.REG_FILE._00554_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10407_  (.A0(\u_cpu.REG_FILE.rf[16][11] ),
    .A1(\u_cpu.REG_FILE._04668_ ),
    .S(\u_cpu.REG_FILE._05120_ ),
    .X(\u_cpu.REG_FILE._05122_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10408_  (.A(\u_cpu.REG_FILE._05122_ ),
    .X(\u_cpu.REG_FILE._00555_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10409_  (.A0(\u_cpu.REG_FILE.rf[16][12] ),
    .A1(\u_cpu.REG_FILE._04670_ ),
    .S(\u_cpu.REG_FILE._05120_ ),
    .X(\u_cpu.REG_FILE._05123_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10410_  (.A(\u_cpu.REG_FILE._05123_ ),
    .X(\u_cpu.REG_FILE._00556_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10411_  (.A0(\u_cpu.REG_FILE.rf[16][13] ),
    .A1(\u_cpu.REG_FILE._04672_ ),
    .S(\u_cpu.REG_FILE._05120_ ),
    .X(\u_cpu.REG_FILE._05124_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10412_  (.A(\u_cpu.REG_FILE._05124_ ),
    .X(\u_cpu.REG_FILE._00557_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10413_  (.A0(\u_cpu.REG_FILE.rf[16][14] ),
    .A1(\u_cpu.REG_FILE._04674_ ),
    .S(\u_cpu.REG_FILE._05120_ ),
    .X(\u_cpu.REG_FILE._05125_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10414_  (.A(\u_cpu.REG_FILE._05125_ ),
    .X(\u_cpu.REG_FILE._00558_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10415_  (.A0(\u_cpu.REG_FILE.rf[16][15] ),
    .A1(\u_cpu.REG_FILE._04676_ ),
    .S(\u_cpu.REG_FILE._05120_ ),
    .X(\u_cpu.REG_FILE._05126_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10416_  (.A(\u_cpu.REG_FILE._05126_ ),
    .X(\u_cpu.REG_FILE._00559_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10417_  (.A0(\u_cpu.REG_FILE.rf[16][16] ),
    .A1(\u_cpu.REG_FILE._04678_ ),
    .S(\u_cpu.REG_FILE._05120_ ),
    .X(\u_cpu.REG_FILE._05127_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10418_  (.A(\u_cpu.REG_FILE._05127_ ),
    .X(\u_cpu.REG_FILE._00560_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10419_  (.A0(\u_cpu.REG_FILE.rf[16][17] ),
    .A1(\u_cpu.REG_FILE._04680_ ),
    .S(\u_cpu.REG_FILE._05120_ ),
    .X(\u_cpu.REG_FILE._05128_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10420_  (.A(\u_cpu.REG_FILE._05128_ ),
    .X(\u_cpu.REG_FILE._00561_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10421_  (.A0(\u_cpu.REG_FILE.rf[16][18] ),
    .A1(\u_cpu.REG_FILE._04682_ ),
    .S(\u_cpu.REG_FILE._05120_ ),
    .X(\u_cpu.REG_FILE._05129_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10422_  (.A(\u_cpu.REG_FILE._05129_ ),
    .X(\u_cpu.REG_FILE._00562_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10423_  (.A0(\u_cpu.REG_FILE.rf[16][19] ),
    .A1(\u_cpu.REG_FILE._04684_ ),
    .S(\u_cpu.REG_FILE._05120_ ),
    .X(\u_cpu.REG_FILE._05130_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10424_  (.A(\u_cpu.REG_FILE._05130_ ),
    .X(\u_cpu.REG_FILE._00563_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10425_  (.A(\u_cpu.REG_FILE._05108_ ),
    .X(\u_cpu.REG_FILE._05131_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10426_  (.A0(\u_cpu.REG_FILE.rf[16][20] ),
    .A1(\u_cpu.REG_FILE._04686_ ),
    .S(\u_cpu.REG_FILE._05131_ ),
    .X(\u_cpu.REG_FILE._05132_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10427_  (.A(\u_cpu.REG_FILE._05132_ ),
    .X(\u_cpu.REG_FILE._00564_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10428_  (.A0(\u_cpu.REG_FILE.rf[16][21] ),
    .A1(\u_cpu.REG_FILE._04689_ ),
    .S(\u_cpu.REG_FILE._05131_ ),
    .X(\u_cpu.REG_FILE._05133_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10429_  (.A(\u_cpu.REG_FILE._05133_ ),
    .X(\u_cpu.REG_FILE._00565_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10430_  (.A0(\u_cpu.REG_FILE.rf[16][22] ),
    .A1(\u_cpu.REG_FILE._04691_ ),
    .S(\u_cpu.REG_FILE._05131_ ),
    .X(\u_cpu.REG_FILE._05134_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10431_  (.A(\u_cpu.REG_FILE._05134_ ),
    .X(\u_cpu.REG_FILE._00566_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10432_  (.A0(\u_cpu.REG_FILE.rf[16][23] ),
    .A1(\u_cpu.REG_FILE._04693_ ),
    .S(\u_cpu.REG_FILE._05131_ ),
    .X(\u_cpu.REG_FILE._05135_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10433_  (.A(\u_cpu.REG_FILE._05135_ ),
    .X(\u_cpu.REG_FILE._00567_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10434_  (.A0(\u_cpu.REG_FILE.rf[16][24] ),
    .A1(\u_cpu.REG_FILE._04695_ ),
    .S(\u_cpu.REG_FILE._05131_ ),
    .X(\u_cpu.REG_FILE._05136_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10435_  (.A(\u_cpu.REG_FILE._05136_ ),
    .X(\u_cpu.REG_FILE._00568_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10436_  (.A0(\u_cpu.REG_FILE.rf[16][25] ),
    .A1(\u_cpu.REG_FILE._04697_ ),
    .S(\u_cpu.REG_FILE._05131_ ),
    .X(\u_cpu.REG_FILE._05137_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10437_  (.A(\u_cpu.REG_FILE._05137_ ),
    .X(\u_cpu.REG_FILE._00569_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10438_  (.A0(\u_cpu.REG_FILE.rf[16][26] ),
    .A1(\u_cpu.REG_FILE._04699_ ),
    .S(\u_cpu.REG_FILE._05131_ ),
    .X(\u_cpu.REG_FILE._05138_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10439_  (.A(\u_cpu.REG_FILE._05138_ ),
    .X(\u_cpu.REG_FILE._00570_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10440_  (.A0(\u_cpu.REG_FILE.rf[16][27] ),
    .A1(\u_cpu.REG_FILE._04701_ ),
    .S(\u_cpu.REG_FILE._05131_ ),
    .X(\u_cpu.REG_FILE._05139_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10441_  (.A(\u_cpu.REG_FILE._05139_ ),
    .X(\u_cpu.REG_FILE._00571_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10442_  (.A0(\u_cpu.REG_FILE.rf[16][28] ),
    .A1(\u_cpu.REG_FILE._04703_ ),
    .S(\u_cpu.REG_FILE._05131_ ),
    .X(\u_cpu.REG_FILE._05140_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10443_  (.A(\u_cpu.REG_FILE._05140_ ),
    .X(\u_cpu.REG_FILE._00572_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10444_  (.A0(\u_cpu.REG_FILE.rf[16][29] ),
    .A1(\u_cpu.REG_FILE._04705_ ),
    .S(\u_cpu.REG_FILE._05131_ ),
    .X(\u_cpu.REG_FILE._05141_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10445_  (.A(\u_cpu.REG_FILE._05141_ ),
    .X(\u_cpu.REG_FILE._00573_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10446_  (.A0(\u_cpu.REG_FILE.rf[16][30] ),
    .A1(\u_cpu.REG_FILE._04707_ ),
    .S(\u_cpu.REG_FILE._05108_ ),
    .X(\u_cpu.REG_FILE._05142_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10447_  (.A(\u_cpu.REG_FILE._05142_ ),
    .X(\u_cpu.REG_FILE._00574_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10448_  (.A0(\u_cpu.REG_FILE.rf[16][31] ),
    .A1(\u_cpu.REG_FILE._04709_ ),
    .S(\u_cpu.REG_FILE._05108_ ),
    .X(\u_cpu.REG_FILE._05143_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10449_  (.A(\u_cpu.REG_FILE._05143_ ),
    .X(\u_cpu.REG_FILE._00575_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu.REG_FILE._10450_  (.A(\u_cpu.REG_FILE._04496_ ),
    .B(\u_cpu.REG_FILE._04423_ ),
    .C(\u_cpu.REG_FILE._05107_ ),
    .Y(\u_cpu.REG_FILE._05144_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10451_  (.A(\u_cpu.REG_FILE._05144_ ),
    .X(\u_cpu.REG_FILE._05145_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10452_  (.A0(\u_cpu.REG_FILE._04420_ ),
    .A1(\u_cpu.REG_FILE.rf[17][0] ),
    .S(\u_cpu.REG_FILE._05145_ ),
    .X(\u_cpu.REG_FILE._05146_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10453_  (.A(\u_cpu.REG_FILE._05146_ ),
    .X(\u_cpu.REG_FILE._00576_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10454_  (.A0(\u_cpu.REG_FILE._04430_ ),
    .A1(\u_cpu.REG_FILE.rf[17][1] ),
    .S(\u_cpu.REG_FILE._05145_ ),
    .X(\u_cpu.REG_FILE._05147_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10455_  (.A(\u_cpu.REG_FILE._05147_ ),
    .X(\u_cpu.REG_FILE._00577_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10456_  (.A0(\u_cpu.REG_FILE._04432_ ),
    .A1(\u_cpu.REG_FILE.rf[17][2] ),
    .S(\u_cpu.REG_FILE._05145_ ),
    .X(\u_cpu.REG_FILE._05148_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10457_  (.A(\u_cpu.REG_FILE._05148_ ),
    .X(\u_cpu.REG_FILE._00578_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10458_  (.A0(\u_cpu.REG_FILE._04434_ ),
    .A1(\u_cpu.REG_FILE.rf[17][3] ),
    .S(\u_cpu.REG_FILE._05145_ ),
    .X(\u_cpu.REG_FILE._05149_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10459_  (.A(\u_cpu.REG_FILE._05149_ ),
    .X(\u_cpu.REG_FILE._00579_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10460_  (.A0(\u_cpu.REG_FILE._04436_ ),
    .A1(\u_cpu.REG_FILE.rf[17][4] ),
    .S(\u_cpu.REG_FILE._05145_ ),
    .X(\u_cpu.REG_FILE._05150_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10461_  (.A(\u_cpu.REG_FILE._05150_ ),
    .X(\u_cpu.REG_FILE._00580_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10462_  (.A0(\u_cpu.REG_FILE._04438_ ),
    .A1(\u_cpu.REG_FILE.rf[17][5] ),
    .S(\u_cpu.REG_FILE._05145_ ),
    .X(\u_cpu.REG_FILE._05151_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10463_  (.A(\u_cpu.REG_FILE._05151_ ),
    .X(\u_cpu.REG_FILE._00581_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10464_  (.A0(\u_cpu.REG_FILE._04440_ ),
    .A1(\u_cpu.REG_FILE.rf[17][6] ),
    .S(\u_cpu.REG_FILE._05145_ ),
    .X(\u_cpu.REG_FILE._05152_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10465_  (.A(\u_cpu.REG_FILE._05152_ ),
    .X(\u_cpu.REG_FILE._00582_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10466_  (.A0(\u_cpu.REG_FILE._04442_ ),
    .A1(\u_cpu.REG_FILE.rf[17][7] ),
    .S(\u_cpu.REG_FILE._05145_ ),
    .X(\u_cpu.REG_FILE._05153_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10467_  (.A(\u_cpu.REG_FILE._05153_ ),
    .X(\u_cpu.REG_FILE._00583_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10468_  (.A0(\u_cpu.REG_FILE._04444_ ),
    .A1(\u_cpu.REG_FILE.rf[17][8] ),
    .S(\u_cpu.REG_FILE._05145_ ),
    .X(\u_cpu.REG_FILE._05154_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10469_  (.A(\u_cpu.REG_FILE._05154_ ),
    .X(\u_cpu.REG_FILE._00584_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10470_  (.A0(\u_cpu.REG_FILE._04446_ ),
    .A1(\u_cpu.REG_FILE.rf[17][9] ),
    .S(\u_cpu.REG_FILE._05145_ ),
    .X(\u_cpu.REG_FILE._05155_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10471_  (.A(\u_cpu.REG_FILE._05155_ ),
    .X(\u_cpu.REG_FILE._00585_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10472_  (.A(\u_cpu.REG_FILE._05144_ ),
    .X(\u_cpu.REG_FILE._05156_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10473_  (.A0(\u_cpu.REG_FILE._04448_ ),
    .A1(\u_cpu.REG_FILE.rf[17][10] ),
    .S(\u_cpu.REG_FILE._05156_ ),
    .X(\u_cpu.REG_FILE._05157_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10474_  (.A(\u_cpu.REG_FILE._05157_ ),
    .X(\u_cpu.REG_FILE._00586_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10475_  (.A0(\u_cpu.REG_FILE._04451_ ),
    .A1(\u_cpu.REG_FILE.rf[17][11] ),
    .S(\u_cpu.REG_FILE._05156_ ),
    .X(\u_cpu.REG_FILE._05158_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10476_  (.A(\u_cpu.REG_FILE._05158_ ),
    .X(\u_cpu.REG_FILE._00587_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10477_  (.A0(\u_cpu.REG_FILE._04453_ ),
    .A1(\u_cpu.REG_FILE.rf[17][12] ),
    .S(\u_cpu.REG_FILE._05156_ ),
    .X(\u_cpu.REG_FILE._05159_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10478_  (.A(\u_cpu.REG_FILE._05159_ ),
    .X(\u_cpu.REG_FILE._00588_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10479_  (.A0(\u_cpu.REG_FILE._04455_ ),
    .A1(\u_cpu.REG_FILE.rf[17][13] ),
    .S(\u_cpu.REG_FILE._05156_ ),
    .X(\u_cpu.REG_FILE._05160_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10480_  (.A(\u_cpu.REG_FILE._05160_ ),
    .X(\u_cpu.REG_FILE._00589_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10481_  (.A0(\u_cpu.REG_FILE._04457_ ),
    .A1(\u_cpu.REG_FILE.rf[17][14] ),
    .S(\u_cpu.REG_FILE._05156_ ),
    .X(\u_cpu.REG_FILE._05161_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10482_  (.A(\u_cpu.REG_FILE._05161_ ),
    .X(\u_cpu.REG_FILE._00590_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10483_  (.A0(\u_cpu.REG_FILE._04459_ ),
    .A1(\u_cpu.REG_FILE.rf[17][15] ),
    .S(\u_cpu.REG_FILE._05156_ ),
    .X(\u_cpu.REG_FILE._05162_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10484_  (.A(\u_cpu.REG_FILE._05162_ ),
    .X(\u_cpu.REG_FILE._00591_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10485_  (.A0(\u_cpu.REG_FILE._04461_ ),
    .A1(\u_cpu.REG_FILE.rf[17][16] ),
    .S(\u_cpu.REG_FILE._05156_ ),
    .X(\u_cpu.REG_FILE._05163_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10486_  (.A(\u_cpu.REG_FILE._05163_ ),
    .X(\u_cpu.REG_FILE._00592_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10487_  (.A0(\u_cpu.REG_FILE._04463_ ),
    .A1(\u_cpu.REG_FILE.rf[17][17] ),
    .S(\u_cpu.REG_FILE._05156_ ),
    .X(\u_cpu.REG_FILE._05164_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10488_  (.A(\u_cpu.REG_FILE._05164_ ),
    .X(\u_cpu.REG_FILE._00593_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10489_  (.A0(\u_cpu.REG_FILE._04465_ ),
    .A1(\u_cpu.REG_FILE.rf[17][18] ),
    .S(\u_cpu.REG_FILE._05156_ ),
    .X(\u_cpu.REG_FILE._05165_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10490_  (.A(\u_cpu.REG_FILE._05165_ ),
    .X(\u_cpu.REG_FILE._00594_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10491_  (.A0(\u_cpu.REG_FILE._04467_ ),
    .A1(\u_cpu.REG_FILE.rf[17][19] ),
    .S(\u_cpu.REG_FILE._05156_ ),
    .X(\u_cpu.REG_FILE._05166_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10492_  (.A(\u_cpu.REG_FILE._05166_ ),
    .X(\u_cpu.REG_FILE._00595_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10493_  (.A(\u_cpu.REG_FILE._05144_ ),
    .X(\u_cpu.REG_FILE._05167_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10494_  (.A0(\u_cpu.REG_FILE._04469_ ),
    .A1(\u_cpu.REG_FILE.rf[17][20] ),
    .S(\u_cpu.REG_FILE._05167_ ),
    .X(\u_cpu.REG_FILE._05168_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10495_  (.A(\u_cpu.REG_FILE._05168_ ),
    .X(\u_cpu.REG_FILE._00596_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10496_  (.A0(\u_cpu.REG_FILE._04472_ ),
    .A1(\u_cpu.REG_FILE.rf[17][21] ),
    .S(\u_cpu.REG_FILE._05167_ ),
    .X(\u_cpu.REG_FILE._05169_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10497_  (.A(\u_cpu.REG_FILE._05169_ ),
    .X(\u_cpu.REG_FILE._00597_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10498_  (.A0(\u_cpu.REG_FILE._04474_ ),
    .A1(\u_cpu.REG_FILE.rf[17][22] ),
    .S(\u_cpu.REG_FILE._05167_ ),
    .X(\u_cpu.REG_FILE._05170_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10499_  (.A(\u_cpu.REG_FILE._05170_ ),
    .X(\u_cpu.REG_FILE._00598_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10500_  (.A0(\u_cpu.REG_FILE._04476_ ),
    .A1(\u_cpu.REG_FILE.rf[17][23] ),
    .S(\u_cpu.REG_FILE._05167_ ),
    .X(\u_cpu.REG_FILE._05171_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10501_  (.A(\u_cpu.REG_FILE._05171_ ),
    .X(\u_cpu.REG_FILE._00599_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10502_  (.A0(\u_cpu.REG_FILE._04478_ ),
    .A1(\u_cpu.REG_FILE.rf[17][24] ),
    .S(\u_cpu.REG_FILE._05167_ ),
    .X(\u_cpu.REG_FILE._05172_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10503_  (.A(\u_cpu.REG_FILE._05172_ ),
    .X(\u_cpu.REG_FILE._00600_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10504_  (.A0(\u_cpu.REG_FILE._04480_ ),
    .A1(\u_cpu.REG_FILE.rf[17][25] ),
    .S(\u_cpu.REG_FILE._05167_ ),
    .X(\u_cpu.REG_FILE._05173_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10505_  (.A(\u_cpu.REG_FILE._05173_ ),
    .X(\u_cpu.REG_FILE._00601_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10506_  (.A0(\u_cpu.REG_FILE._04482_ ),
    .A1(\u_cpu.REG_FILE.rf[17][26] ),
    .S(\u_cpu.REG_FILE._05167_ ),
    .X(\u_cpu.REG_FILE._05174_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10507_  (.A(\u_cpu.REG_FILE._05174_ ),
    .X(\u_cpu.REG_FILE._00602_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10508_  (.A0(\u_cpu.REG_FILE._04484_ ),
    .A1(\u_cpu.REG_FILE.rf[17][27] ),
    .S(\u_cpu.REG_FILE._05167_ ),
    .X(\u_cpu.REG_FILE._05175_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10509_  (.A(\u_cpu.REG_FILE._05175_ ),
    .X(\u_cpu.REG_FILE._00603_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10510_  (.A0(\u_cpu.REG_FILE._04486_ ),
    .A1(\u_cpu.REG_FILE.rf[17][28] ),
    .S(\u_cpu.REG_FILE._05167_ ),
    .X(\u_cpu.REG_FILE._05176_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10511_  (.A(\u_cpu.REG_FILE._05176_ ),
    .X(\u_cpu.REG_FILE._00604_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10512_  (.A0(\u_cpu.REG_FILE._04488_ ),
    .A1(\u_cpu.REG_FILE.rf[17][29] ),
    .S(\u_cpu.REG_FILE._05167_ ),
    .X(\u_cpu.REG_FILE._05177_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10513_  (.A(\u_cpu.REG_FILE._05177_ ),
    .X(\u_cpu.REG_FILE._00605_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10514_  (.A0(\u_cpu.REG_FILE._04490_ ),
    .A1(\u_cpu.REG_FILE.rf[17][30] ),
    .S(\u_cpu.REG_FILE._05144_ ),
    .X(\u_cpu.REG_FILE._05178_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10515_  (.A(\u_cpu.REG_FILE._05178_ ),
    .X(\u_cpu.REG_FILE._00606_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10516_  (.A0(\u_cpu.REG_FILE._04492_ ),
    .A1(\u_cpu.REG_FILE.rf[17][31] ),
    .S(\u_cpu.REG_FILE._05144_ ),
    .X(\u_cpu.REG_FILE._05179_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10517_  (.A(\u_cpu.REG_FILE._05179_ ),
    .X(\u_cpu.REG_FILE._00607_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu.REG_FILE._10518_  (.A(\u_cpu.REG_FILE._04496_ ),
    .B(\u_cpu.REG_FILE._05107_ ),
    .C(\u_cpu.REG_FILE._04747_ ),
    .X(\u_cpu.REG_FILE._05180_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10519_  (.A(\u_cpu.REG_FILE._05180_ ),
    .X(\u_cpu.REG_FILE._05181_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10520_  (.A0(\u_cpu.REG_FILE.rf[18][0] ),
    .A1(\u_cpu.REG_FILE._04642_ ),
    .S(\u_cpu.REG_FILE._05181_ ),
    .X(\u_cpu.REG_FILE._05182_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10521_  (.A(\u_cpu.REG_FILE._05182_ ),
    .X(\u_cpu.REG_FILE._00608_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10522_  (.A0(\u_cpu.REG_FILE.rf[18][1] ),
    .A1(\u_cpu.REG_FILE._04647_ ),
    .S(\u_cpu.REG_FILE._05181_ ),
    .X(\u_cpu.REG_FILE._05183_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10523_  (.A(\u_cpu.REG_FILE._05183_ ),
    .X(\u_cpu.REG_FILE._00609_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10524_  (.A0(\u_cpu.REG_FILE.rf[18][2] ),
    .A1(\u_cpu.REG_FILE._04649_ ),
    .S(\u_cpu.REG_FILE._05181_ ),
    .X(\u_cpu.REG_FILE._05184_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10525_  (.A(\u_cpu.REG_FILE._05184_ ),
    .X(\u_cpu.REG_FILE._00610_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10526_  (.A0(\u_cpu.REG_FILE.rf[18][3] ),
    .A1(\u_cpu.REG_FILE._04651_ ),
    .S(\u_cpu.REG_FILE._05181_ ),
    .X(\u_cpu.REG_FILE._05185_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10527_  (.A(\u_cpu.REG_FILE._05185_ ),
    .X(\u_cpu.REG_FILE._00611_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10528_  (.A0(\u_cpu.REG_FILE.rf[18][4] ),
    .A1(\u_cpu.REG_FILE._04653_ ),
    .S(\u_cpu.REG_FILE._05181_ ),
    .X(\u_cpu.REG_FILE._05186_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10529_  (.A(\u_cpu.REG_FILE._05186_ ),
    .X(\u_cpu.REG_FILE._00612_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10530_  (.A0(\u_cpu.REG_FILE.rf[18][5] ),
    .A1(\u_cpu.REG_FILE._04655_ ),
    .S(\u_cpu.REG_FILE._05181_ ),
    .X(\u_cpu.REG_FILE._05187_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10531_  (.A(\u_cpu.REG_FILE._05187_ ),
    .X(\u_cpu.REG_FILE._00613_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10532_  (.A0(\u_cpu.REG_FILE.rf[18][6] ),
    .A1(\u_cpu.REG_FILE._04657_ ),
    .S(\u_cpu.REG_FILE._05181_ ),
    .X(\u_cpu.REG_FILE._05188_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10533_  (.A(\u_cpu.REG_FILE._05188_ ),
    .X(\u_cpu.REG_FILE._00614_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10534_  (.A0(\u_cpu.REG_FILE.rf[18][7] ),
    .A1(\u_cpu.REG_FILE._04659_ ),
    .S(\u_cpu.REG_FILE._05181_ ),
    .X(\u_cpu.REG_FILE._05189_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10535_  (.A(\u_cpu.REG_FILE._05189_ ),
    .X(\u_cpu.REG_FILE._00615_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10536_  (.A0(\u_cpu.REG_FILE.rf[18][8] ),
    .A1(\u_cpu.REG_FILE._04661_ ),
    .S(\u_cpu.REG_FILE._05181_ ),
    .X(\u_cpu.REG_FILE._05190_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10537_  (.A(\u_cpu.REG_FILE._05190_ ),
    .X(\u_cpu.REG_FILE._00616_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10538_  (.A0(\u_cpu.REG_FILE.rf[18][9] ),
    .A1(\u_cpu.REG_FILE._04663_ ),
    .S(\u_cpu.REG_FILE._05181_ ),
    .X(\u_cpu.REG_FILE._05191_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10539_  (.A(\u_cpu.REG_FILE._05191_ ),
    .X(\u_cpu.REG_FILE._00617_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10540_  (.A(\u_cpu.REG_FILE._05180_ ),
    .X(\u_cpu.REG_FILE._05192_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10541_  (.A0(\u_cpu.REG_FILE.rf[18][10] ),
    .A1(\u_cpu.REG_FILE._04665_ ),
    .S(\u_cpu.REG_FILE._05192_ ),
    .X(\u_cpu.REG_FILE._05193_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10542_  (.A(\u_cpu.REG_FILE._05193_ ),
    .X(\u_cpu.REG_FILE._00618_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10543_  (.A0(\u_cpu.REG_FILE.rf[18][11] ),
    .A1(\u_cpu.REG_FILE._04668_ ),
    .S(\u_cpu.REG_FILE._05192_ ),
    .X(\u_cpu.REG_FILE._05194_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10544_  (.A(\u_cpu.REG_FILE._05194_ ),
    .X(\u_cpu.REG_FILE._00619_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10545_  (.A0(\u_cpu.REG_FILE.rf[18][12] ),
    .A1(\u_cpu.REG_FILE._04670_ ),
    .S(\u_cpu.REG_FILE._05192_ ),
    .X(\u_cpu.REG_FILE._05195_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10546_  (.A(\u_cpu.REG_FILE._05195_ ),
    .X(\u_cpu.REG_FILE._00620_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10547_  (.A0(\u_cpu.REG_FILE.rf[18][13] ),
    .A1(\u_cpu.REG_FILE._04672_ ),
    .S(\u_cpu.REG_FILE._05192_ ),
    .X(\u_cpu.REG_FILE._05196_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10548_  (.A(\u_cpu.REG_FILE._05196_ ),
    .X(\u_cpu.REG_FILE._00621_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10549_  (.A0(\u_cpu.REG_FILE.rf[18][14] ),
    .A1(\u_cpu.REG_FILE._04674_ ),
    .S(\u_cpu.REG_FILE._05192_ ),
    .X(\u_cpu.REG_FILE._05197_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10550_  (.A(\u_cpu.REG_FILE._05197_ ),
    .X(\u_cpu.REG_FILE._00622_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10551_  (.A0(\u_cpu.REG_FILE.rf[18][15] ),
    .A1(\u_cpu.REG_FILE._04676_ ),
    .S(\u_cpu.REG_FILE._05192_ ),
    .X(\u_cpu.REG_FILE._05198_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10552_  (.A(\u_cpu.REG_FILE._05198_ ),
    .X(\u_cpu.REG_FILE._00623_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10553_  (.A0(\u_cpu.REG_FILE.rf[18][16] ),
    .A1(\u_cpu.REG_FILE._04678_ ),
    .S(\u_cpu.REG_FILE._05192_ ),
    .X(\u_cpu.REG_FILE._05199_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10554_  (.A(\u_cpu.REG_FILE._05199_ ),
    .X(\u_cpu.REG_FILE._00624_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10555_  (.A0(\u_cpu.REG_FILE.rf[18][17] ),
    .A1(\u_cpu.REG_FILE._04680_ ),
    .S(\u_cpu.REG_FILE._05192_ ),
    .X(\u_cpu.REG_FILE._05200_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10556_  (.A(\u_cpu.REG_FILE._05200_ ),
    .X(\u_cpu.REG_FILE._00625_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10557_  (.A0(\u_cpu.REG_FILE.rf[18][18] ),
    .A1(\u_cpu.REG_FILE._04682_ ),
    .S(\u_cpu.REG_FILE._05192_ ),
    .X(\u_cpu.REG_FILE._05201_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10558_  (.A(\u_cpu.REG_FILE._05201_ ),
    .X(\u_cpu.REG_FILE._00626_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10559_  (.A0(\u_cpu.REG_FILE.rf[18][19] ),
    .A1(\u_cpu.REG_FILE._04684_ ),
    .S(\u_cpu.REG_FILE._05192_ ),
    .X(\u_cpu.REG_FILE._05202_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10560_  (.A(\u_cpu.REG_FILE._05202_ ),
    .X(\u_cpu.REG_FILE._00627_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10561_  (.A(\u_cpu.REG_FILE._05180_ ),
    .X(\u_cpu.REG_FILE._05203_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10562_  (.A0(\u_cpu.REG_FILE.rf[18][20] ),
    .A1(\u_cpu.REG_FILE._04686_ ),
    .S(\u_cpu.REG_FILE._05203_ ),
    .X(\u_cpu.REG_FILE._05204_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10563_  (.A(\u_cpu.REG_FILE._05204_ ),
    .X(\u_cpu.REG_FILE._00628_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10564_  (.A0(\u_cpu.REG_FILE.rf[18][21] ),
    .A1(\u_cpu.REG_FILE._04689_ ),
    .S(\u_cpu.REG_FILE._05203_ ),
    .X(\u_cpu.REG_FILE._05205_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10565_  (.A(\u_cpu.REG_FILE._05205_ ),
    .X(\u_cpu.REG_FILE._00629_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10566_  (.A0(\u_cpu.REG_FILE.rf[18][22] ),
    .A1(\u_cpu.REG_FILE._04691_ ),
    .S(\u_cpu.REG_FILE._05203_ ),
    .X(\u_cpu.REG_FILE._05206_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10567_  (.A(\u_cpu.REG_FILE._05206_ ),
    .X(\u_cpu.REG_FILE._00630_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10568_  (.A0(\u_cpu.REG_FILE.rf[18][23] ),
    .A1(\u_cpu.REG_FILE._04693_ ),
    .S(\u_cpu.REG_FILE._05203_ ),
    .X(\u_cpu.REG_FILE._05207_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10569_  (.A(\u_cpu.REG_FILE._05207_ ),
    .X(\u_cpu.REG_FILE._00631_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10570_  (.A0(\u_cpu.REG_FILE.rf[18][24] ),
    .A1(\u_cpu.REG_FILE._04695_ ),
    .S(\u_cpu.REG_FILE._05203_ ),
    .X(\u_cpu.REG_FILE._05208_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10571_  (.A(\u_cpu.REG_FILE._05208_ ),
    .X(\u_cpu.REG_FILE._00632_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10572_  (.A0(\u_cpu.REG_FILE.rf[18][25] ),
    .A1(\u_cpu.REG_FILE._04697_ ),
    .S(\u_cpu.REG_FILE._05203_ ),
    .X(\u_cpu.REG_FILE._05209_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10573_  (.A(\u_cpu.REG_FILE._05209_ ),
    .X(\u_cpu.REG_FILE._00633_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10574_  (.A0(\u_cpu.REG_FILE.rf[18][26] ),
    .A1(\u_cpu.REG_FILE._04699_ ),
    .S(\u_cpu.REG_FILE._05203_ ),
    .X(\u_cpu.REG_FILE._05210_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10575_  (.A(\u_cpu.REG_FILE._05210_ ),
    .X(\u_cpu.REG_FILE._00634_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10576_  (.A0(\u_cpu.REG_FILE.rf[18][27] ),
    .A1(\u_cpu.REG_FILE._04701_ ),
    .S(\u_cpu.REG_FILE._05203_ ),
    .X(\u_cpu.REG_FILE._05211_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10577_  (.A(\u_cpu.REG_FILE._05211_ ),
    .X(\u_cpu.REG_FILE._00635_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10578_  (.A0(\u_cpu.REG_FILE.rf[18][28] ),
    .A1(\u_cpu.REG_FILE._04703_ ),
    .S(\u_cpu.REG_FILE._05203_ ),
    .X(\u_cpu.REG_FILE._05212_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10579_  (.A(\u_cpu.REG_FILE._05212_ ),
    .X(\u_cpu.REG_FILE._00636_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10580_  (.A0(\u_cpu.REG_FILE.rf[18][29] ),
    .A1(\u_cpu.REG_FILE._04705_ ),
    .S(\u_cpu.REG_FILE._05203_ ),
    .X(\u_cpu.REG_FILE._05213_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10581_  (.A(\u_cpu.REG_FILE._05213_ ),
    .X(\u_cpu.REG_FILE._00637_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10582_  (.A0(\u_cpu.REG_FILE.rf[18][30] ),
    .A1(\u_cpu.REG_FILE._04707_ ),
    .S(\u_cpu.REG_FILE._05180_ ),
    .X(\u_cpu.REG_FILE._05214_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10583_  (.A(\u_cpu.REG_FILE._05214_ ),
    .X(\u_cpu.REG_FILE._00638_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10584_  (.A0(\u_cpu.REG_FILE.rf[18][31] ),
    .A1(\u_cpu.REG_FILE._04709_ ),
    .S(\u_cpu.REG_FILE._05180_ ),
    .X(\u_cpu.REG_FILE._05215_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10585_  (.A(\u_cpu.REG_FILE._05215_ ),
    .X(\u_cpu.REG_FILE._00639_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10586_  (.A(\u_cpu.REG_FILE.wd3[0] ),
    .X(\u_cpu.REG_FILE._05216_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.REG_FILE._10587_  (.A_N(\u_cpu.REG_FILE.a3[1] ),
    .B(\u_cpu.REG_FILE.a3[0] ),
    .C(\u_cpu.REG_FILE.we3 ),
    .D(\u_cpu.REG_FILE._04605_ ),
    .X(\u_cpu.REG_FILE._05217_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10588_  (.A(\u_cpu.REG_FILE._05217_ ),
    .X(\u_cpu.REG_FILE._05218_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10589_  (.A(\u_cpu.REG_FILE._05218_ ),
    .X(\u_cpu.REG_FILE._05219_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10590_  (.A0(\u_cpu.REG_FILE.rf[1][0] ),
    .A1(\u_cpu.REG_FILE._05216_ ),
    .S(\u_cpu.REG_FILE._05219_ ),
    .X(\u_cpu.REG_FILE._05220_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10591_  (.A(\u_cpu.REG_FILE._05220_ ),
    .X(\u_cpu.REG_FILE._00640_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10592_  (.A(\u_cpu.REG_FILE.wd3[1] ),
    .X(\u_cpu.REG_FILE._05221_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10593_  (.A0(\u_cpu.REG_FILE.rf[1][1] ),
    .A1(\u_cpu.REG_FILE._05221_ ),
    .S(\u_cpu.REG_FILE._05219_ ),
    .X(\u_cpu.REG_FILE._05222_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10594_  (.A(\u_cpu.REG_FILE._05222_ ),
    .X(\u_cpu.REG_FILE._00641_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10595_  (.A(\u_cpu.REG_FILE.wd3[2] ),
    .X(\u_cpu.REG_FILE._05223_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10596_  (.A0(\u_cpu.REG_FILE.rf[1][2] ),
    .A1(\u_cpu.REG_FILE._05223_ ),
    .S(\u_cpu.REG_FILE._05219_ ),
    .X(\u_cpu.REG_FILE._05224_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10597_  (.A(\u_cpu.REG_FILE._05224_ ),
    .X(\u_cpu.REG_FILE._00642_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10598_  (.A(\u_cpu.REG_FILE.wd3[3] ),
    .X(\u_cpu.REG_FILE._05225_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10599_  (.A0(\u_cpu.REG_FILE.rf[1][3] ),
    .A1(\u_cpu.REG_FILE._05225_ ),
    .S(\u_cpu.REG_FILE._05219_ ),
    .X(\u_cpu.REG_FILE._05226_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10600_  (.A(\u_cpu.REG_FILE._05226_ ),
    .X(\u_cpu.REG_FILE._00643_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10601_  (.A(\u_cpu.REG_FILE.wd3[4] ),
    .X(\u_cpu.REG_FILE._05227_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10602_  (.A0(\u_cpu.REG_FILE.rf[1][4] ),
    .A1(\u_cpu.REG_FILE._05227_ ),
    .S(\u_cpu.REG_FILE._05219_ ),
    .X(\u_cpu.REG_FILE._05228_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10603_  (.A(\u_cpu.REG_FILE._05228_ ),
    .X(\u_cpu.REG_FILE._00644_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10604_  (.A(\u_cpu.REG_FILE.wd3[5] ),
    .X(\u_cpu.REG_FILE._05229_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10605_  (.A0(\u_cpu.REG_FILE.rf[1][5] ),
    .A1(\u_cpu.REG_FILE._05229_ ),
    .S(\u_cpu.REG_FILE._05219_ ),
    .X(\u_cpu.REG_FILE._05230_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10606_  (.A(\u_cpu.REG_FILE._05230_ ),
    .X(\u_cpu.REG_FILE._00645_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10607_  (.A(\u_cpu.REG_FILE.wd3[6] ),
    .X(\u_cpu.REG_FILE._05231_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10608_  (.A0(\u_cpu.REG_FILE.rf[1][6] ),
    .A1(\u_cpu.REG_FILE._05231_ ),
    .S(\u_cpu.REG_FILE._05219_ ),
    .X(\u_cpu.REG_FILE._05232_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10609_  (.A(\u_cpu.REG_FILE._05232_ ),
    .X(\u_cpu.REG_FILE._00646_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10610_  (.A(\u_cpu.REG_FILE.wd3[7] ),
    .X(\u_cpu.REG_FILE._05233_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10611_  (.A0(\u_cpu.REG_FILE.rf[1][7] ),
    .A1(\u_cpu.REG_FILE._05233_ ),
    .S(\u_cpu.REG_FILE._05219_ ),
    .X(\u_cpu.REG_FILE._05234_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10612_  (.A(\u_cpu.REG_FILE._05234_ ),
    .X(\u_cpu.REG_FILE._00647_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10613_  (.A(\u_cpu.REG_FILE.wd3[8] ),
    .X(\u_cpu.REG_FILE._05235_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10614_  (.A0(\u_cpu.REG_FILE.rf[1][8] ),
    .A1(\u_cpu.REG_FILE._05235_ ),
    .S(\u_cpu.REG_FILE._05219_ ),
    .X(\u_cpu.REG_FILE._05236_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10615_  (.A(\u_cpu.REG_FILE._05236_ ),
    .X(\u_cpu.REG_FILE._00648_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10616_  (.A(\u_cpu.REG_FILE.wd3[9] ),
    .X(\u_cpu.REG_FILE._05237_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10617_  (.A0(\u_cpu.REG_FILE.rf[1][9] ),
    .A1(\u_cpu.REG_FILE._05237_ ),
    .S(\u_cpu.REG_FILE._05219_ ),
    .X(\u_cpu.REG_FILE._05238_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10618_  (.A(\u_cpu.REG_FILE._05238_ ),
    .X(\u_cpu.REG_FILE._00649_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10619_  (.A(\u_cpu.REG_FILE.wd3[10] ),
    .X(\u_cpu.REG_FILE._05239_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10620_  (.A(\u_cpu.REG_FILE._05218_ ),
    .X(\u_cpu.REG_FILE._05240_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10621_  (.A0(\u_cpu.REG_FILE.rf[1][10] ),
    .A1(\u_cpu.REG_FILE._05239_ ),
    .S(\u_cpu.REG_FILE._05240_ ),
    .X(\u_cpu.REG_FILE._05241_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10622_  (.A(\u_cpu.REG_FILE._05241_ ),
    .X(\u_cpu.REG_FILE._00650_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10623_  (.A(\u_cpu.REG_FILE.wd3[11] ),
    .X(\u_cpu.REG_FILE._05242_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10624_  (.A0(\u_cpu.REG_FILE.rf[1][11] ),
    .A1(\u_cpu.REG_FILE._05242_ ),
    .S(\u_cpu.REG_FILE._05240_ ),
    .X(\u_cpu.REG_FILE._05243_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10625_  (.A(\u_cpu.REG_FILE._05243_ ),
    .X(\u_cpu.REG_FILE._00651_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10626_  (.A(\u_cpu.REG_FILE.wd3[12] ),
    .X(\u_cpu.REG_FILE._05244_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10627_  (.A0(\u_cpu.REG_FILE.rf[1][12] ),
    .A1(\u_cpu.REG_FILE._05244_ ),
    .S(\u_cpu.REG_FILE._05240_ ),
    .X(\u_cpu.REG_FILE._05245_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10628_  (.A(\u_cpu.REG_FILE._05245_ ),
    .X(\u_cpu.REG_FILE._00652_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10629_  (.A(\u_cpu.REG_FILE.wd3[13] ),
    .X(\u_cpu.REG_FILE._05246_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10630_  (.A0(\u_cpu.REG_FILE.rf[1][13] ),
    .A1(\u_cpu.REG_FILE._05246_ ),
    .S(\u_cpu.REG_FILE._05240_ ),
    .X(\u_cpu.REG_FILE._05247_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10631_  (.A(\u_cpu.REG_FILE._05247_ ),
    .X(\u_cpu.REG_FILE._00653_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10632_  (.A(\u_cpu.REG_FILE.wd3[14] ),
    .X(\u_cpu.REG_FILE._05248_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10633_  (.A0(\u_cpu.REG_FILE.rf[1][14] ),
    .A1(\u_cpu.REG_FILE._05248_ ),
    .S(\u_cpu.REG_FILE._05240_ ),
    .X(\u_cpu.REG_FILE._05249_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10634_  (.A(\u_cpu.REG_FILE._05249_ ),
    .X(\u_cpu.REG_FILE._00654_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10635_  (.A(\u_cpu.REG_FILE.wd3[15] ),
    .X(\u_cpu.REG_FILE._05250_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10636_  (.A0(\u_cpu.REG_FILE.rf[1][15] ),
    .A1(\u_cpu.REG_FILE._05250_ ),
    .S(\u_cpu.REG_FILE._05240_ ),
    .X(\u_cpu.REG_FILE._05251_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10637_  (.A(\u_cpu.REG_FILE._05251_ ),
    .X(\u_cpu.REG_FILE._00655_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10638_  (.A(\u_cpu.REG_FILE.wd3[16] ),
    .X(\u_cpu.REG_FILE._05252_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10639_  (.A0(\u_cpu.REG_FILE.rf[1][16] ),
    .A1(\u_cpu.REG_FILE._05252_ ),
    .S(\u_cpu.REG_FILE._05240_ ),
    .X(\u_cpu.REG_FILE._05253_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10640_  (.A(\u_cpu.REG_FILE._05253_ ),
    .X(\u_cpu.REG_FILE._00656_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10641_  (.A(\u_cpu.REG_FILE.wd3[17] ),
    .X(\u_cpu.REG_FILE._05254_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10642_  (.A0(\u_cpu.REG_FILE.rf[1][17] ),
    .A1(\u_cpu.REG_FILE._05254_ ),
    .S(\u_cpu.REG_FILE._05240_ ),
    .X(\u_cpu.REG_FILE._05255_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10643_  (.A(\u_cpu.REG_FILE._05255_ ),
    .X(\u_cpu.REG_FILE._00657_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10644_  (.A(\u_cpu.REG_FILE.wd3[18] ),
    .X(\u_cpu.REG_FILE._05256_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10645_  (.A0(\u_cpu.REG_FILE.rf[1][18] ),
    .A1(\u_cpu.REG_FILE._05256_ ),
    .S(\u_cpu.REG_FILE._05240_ ),
    .X(\u_cpu.REG_FILE._05257_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10646_  (.A(\u_cpu.REG_FILE._05257_ ),
    .X(\u_cpu.REG_FILE._00658_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10647_  (.A(\u_cpu.REG_FILE.wd3[19] ),
    .X(\u_cpu.REG_FILE._05258_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10648_  (.A0(\u_cpu.REG_FILE.rf[1][19] ),
    .A1(\u_cpu.REG_FILE._05258_ ),
    .S(\u_cpu.REG_FILE._05240_ ),
    .X(\u_cpu.REG_FILE._05259_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10649_  (.A(\u_cpu.REG_FILE._05259_ ),
    .X(\u_cpu.REG_FILE._00659_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10650_  (.A(\u_cpu.REG_FILE.wd3[20] ),
    .X(\u_cpu.REG_FILE._05260_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10651_  (.A(\u_cpu.REG_FILE._05218_ ),
    .X(\u_cpu.REG_FILE._05261_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10652_  (.A0(\u_cpu.REG_FILE.rf[1][20] ),
    .A1(\u_cpu.REG_FILE._05260_ ),
    .S(\u_cpu.REG_FILE._05261_ ),
    .X(\u_cpu.REG_FILE._05262_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10653_  (.A(\u_cpu.REG_FILE._05262_ ),
    .X(\u_cpu.REG_FILE._00660_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10654_  (.A(\u_cpu.REG_FILE.wd3[21] ),
    .X(\u_cpu.REG_FILE._05263_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10655_  (.A0(\u_cpu.REG_FILE.rf[1][21] ),
    .A1(\u_cpu.REG_FILE._05263_ ),
    .S(\u_cpu.REG_FILE._05261_ ),
    .X(\u_cpu.REG_FILE._05264_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10656_  (.A(\u_cpu.REG_FILE._05264_ ),
    .X(\u_cpu.REG_FILE._00661_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10657_  (.A(\u_cpu.REG_FILE.wd3[22] ),
    .X(\u_cpu.REG_FILE._05265_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10658_  (.A0(\u_cpu.REG_FILE.rf[1][22] ),
    .A1(\u_cpu.REG_FILE._05265_ ),
    .S(\u_cpu.REG_FILE._05261_ ),
    .X(\u_cpu.REG_FILE._05266_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10659_  (.A(\u_cpu.REG_FILE._05266_ ),
    .X(\u_cpu.REG_FILE._00662_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10660_  (.A(\u_cpu.REG_FILE.wd3[23] ),
    .X(\u_cpu.REG_FILE._05267_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10661_  (.A0(\u_cpu.REG_FILE.rf[1][23] ),
    .A1(\u_cpu.REG_FILE._05267_ ),
    .S(\u_cpu.REG_FILE._05261_ ),
    .X(\u_cpu.REG_FILE._05268_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10662_  (.A(\u_cpu.REG_FILE._05268_ ),
    .X(\u_cpu.REG_FILE._00663_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10663_  (.A(\u_cpu.REG_FILE.wd3[24] ),
    .X(\u_cpu.REG_FILE._05269_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10664_  (.A0(\u_cpu.REG_FILE.rf[1][24] ),
    .A1(\u_cpu.REG_FILE._05269_ ),
    .S(\u_cpu.REG_FILE._05261_ ),
    .X(\u_cpu.REG_FILE._05270_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10665_  (.A(\u_cpu.REG_FILE._05270_ ),
    .X(\u_cpu.REG_FILE._00664_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10666_  (.A(\u_cpu.REG_FILE.wd3[25] ),
    .X(\u_cpu.REG_FILE._05271_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10667_  (.A0(\u_cpu.REG_FILE.rf[1][25] ),
    .A1(\u_cpu.REG_FILE._05271_ ),
    .S(\u_cpu.REG_FILE._05261_ ),
    .X(\u_cpu.REG_FILE._05272_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10668_  (.A(\u_cpu.REG_FILE._05272_ ),
    .X(\u_cpu.REG_FILE._00665_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10669_  (.A(\u_cpu.REG_FILE.wd3[26] ),
    .X(\u_cpu.REG_FILE._05273_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10670_  (.A0(\u_cpu.REG_FILE.rf[1][26] ),
    .A1(\u_cpu.REG_FILE._05273_ ),
    .S(\u_cpu.REG_FILE._05261_ ),
    .X(\u_cpu.REG_FILE._05274_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10671_  (.A(\u_cpu.REG_FILE._05274_ ),
    .X(\u_cpu.REG_FILE._00666_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10672_  (.A(\u_cpu.REG_FILE.wd3[27] ),
    .X(\u_cpu.REG_FILE._05275_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10673_  (.A0(\u_cpu.REG_FILE.rf[1][27] ),
    .A1(\u_cpu.REG_FILE._05275_ ),
    .S(\u_cpu.REG_FILE._05261_ ),
    .X(\u_cpu.REG_FILE._05276_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10674_  (.A(\u_cpu.REG_FILE._05276_ ),
    .X(\u_cpu.REG_FILE._00667_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10675_  (.A(\u_cpu.REG_FILE.wd3[28] ),
    .X(\u_cpu.REG_FILE._05277_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10676_  (.A0(\u_cpu.REG_FILE.rf[1][28] ),
    .A1(\u_cpu.REG_FILE._05277_ ),
    .S(\u_cpu.REG_FILE._05261_ ),
    .X(\u_cpu.REG_FILE._05278_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10677_  (.A(\u_cpu.REG_FILE._05278_ ),
    .X(\u_cpu.REG_FILE._00668_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10678_  (.A(\u_cpu.REG_FILE.wd3[29] ),
    .X(\u_cpu.REG_FILE._05279_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10679_  (.A0(\u_cpu.REG_FILE.rf[1][29] ),
    .A1(\u_cpu.REG_FILE._05279_ ),
    .S(\u_cpu.REG_FILE._05261_ ),
    .X(\u_cpu.REG_FILE._05280_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10680_  (.A(\u_cpu.REG_FILE._05280_ ),
    .X(\u_cpu.REG_FILE._00669_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10681_  (.A(\u_cpu.REG_FILE.wd3[30] ),
    .X(\u_cpu.REG_FILE._05281_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10682_  (.A0(\u_cpu.REG_FILE.rf[1][30] ),
    .A1(\u_cpu.REG_FILE._05281_ ),
    .S(\u_cpu.REG_FILE._05218_ ),
    .X(\u_cpu.REG_FILE._05282_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10683_  (.A(\u_cpu.REG_FILE._05282_ ),
    .X(\u_cpu.REG_FILE._00670_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10684_  (.A(\u_cpu.REG_FILE.wd3[31] ),
    .X(\u_cpu.REG_FILE._05283_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10685_  (.A0(\u_cpu.REG_FILE.rf[1][31] ),
    .A1(\u_cpu.REG_FILE._05283_ ),
    .S(\u_cpu.REG_FILE._05218_ ),
    .X(\u_cpu.REG_FILE._05284_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10686_  (.A(\u_cpu.REG_FILE._05284_ ),
    .X(\u_cpu.REG_FILE._00671_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.REG_FILE._10687_  (.A_N(\u_cpu.REG_FILE._04421_ ),
    .B(\u_cpu.REG_FILE._04425_ ),
    .C(\u_cpu.REG_FILE._04643_ ),
    .D(\u_cpu.REG_FILE.a3[4] ),
    .X(\u_cpu.REG_FILE._05285_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10688_  (.A(\u_cpu.REG_FILE._05285_ ),
    .X(\u_cpu.REG_FILE._05286_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10689_  (.A(\u_cpu.REG_FILE._05286_ ),
    .X(\u_cpu.REG_FILE._05287_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10690_  (.A0(\u_cpu.REG_FILE.rf[20][0] ),
    .A1(\u_cpu.REG_FILE._05216_ ),
    .S(\u_cpu.REG_FILE._05287_ ),
    .X(\u_cpu.REG_FILE._05288_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10691_  (.A(\u_cpu.REG_FILE._05288_ ),
    .X(\u_cpu.REG_FILE._00672_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10692_  (.A0(\u_cpu.REG_FILE.rf[20][1] ),
    .A1(\u_cpu.REG_FILE._05221_ ),
    .S(\u_cpu.REG_FILE._05287_ ),
    .X(\u_cpu.REG_FILE._05289_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10693_  (.A(\u_cpu.REG_FILE._05289_ ),
    .X(\u_cpu.REG_FILE._00673_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10694_  (.A0(\u_cpu.REG_FILE.rf[20][2] ),
    .A1(\u_cpu.REG_FILE._05223_ ),
    .S(\u_cpu.REG_FILE._05287_ ),
    .X(\u_cpu.REG_FILE._05290_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10695_  (.A(\u_cpu.REG_FILE._05290_ ),
    .X(\u_cpu.REG_FILE._00674_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10696_  (.A0(\u_cpu.REG_FILE.rf[20][3] ),
    .A1(\u_cpu.REG_FILE._05225_ ),
    .S(\u_cpu.REG_FILE._05287_ ),
    .X(\u_cpu.REG_FILE._05291_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10697_  (.A(\u_cpu.REG_FILE._05291_ ),
    .X(\u_cpu.REG_FILE._00675_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10698_  (.A0(\u_cpu.REG_FILE.rf[20][4] ),
    .A1(\u_cpu.REG_FILE._05227_ ),
    .S(\u_cpu.REG_FILE._05287_ ),
    .X(\u_cpu.REG_FILE._05292_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10699_  (.A(\u_cpu.REG_FILE._05292_ ),
    .X(\u_cpu.REG_FILE._00676_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10700_  (.A0(\u_cpu.REG_FILE.rf[20][5] ),
    .A1(\u_cpu.REG_FILE._05229_ ),
    .S(\u_cpu.REG_FILE._05287_ ),
    .X(\u_cpu.REG_FILE._05293_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10701_  (.A(\u_cpu.REG_FILE._05293_ ),
    .X(\u_cpu.REG_FILE._00677_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10702_  (.A0(\u_cpu.REG_FILE.rf[20][6] ),
    .A1(\u_cpu.REG_FILE._05231_ ),
    .S(\u_cpu.REG_FILE._05287_ ),
    .X(\u_cpu.REG_FILE._05294_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10703_  (.A(\u_cpu.REG_FILE._05294_ ),
    .X(\u_cpu.REG_FILE._00678_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10704_  (.A0(\u_cpu.REG_FILE.rf[20][7] ),
    .A1(\u_cpu.REG_FILE._05233_ ),
    .S(\u_cpu.REG_FILE._05287_ ),
    .X(\u_cpu.REG_FILE._05295_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10705_  (.A(\u_cpu.REG_FILE._05295_ ),
    .X(\u_cpu.REG_FILE._00679_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10706_  (.A0(\u_cpu.REG_FILE.rf[20][8] ),
    .A1(\u_cpu.REG_FILE._05235_ ),
    .S(\u_cpu.REG_FILE._05287_ ),
    .X(\u_cpu.REG_FILE._05296_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10707_  (.A(\u_cpu.REG_FILE._05296_ ),
    .X(\u_cpu.REG_FILE._00680_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10708_  (.A0(\u_cpu.REG_FILE.rf[20][9] ),
    .A1(\u_cpu.REG_FILE._05237_ ),
    .S(\u_cpu.REG_FILE._05287_ ),
    .X(\u_cpu.REG_FILE._05297_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10709_  (.A(\u_cpu.REG_FILE._05297_ ),
    .X(\u_cpu.REG_FILE._00681_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10710_  (.A(\u_cpu.REG_FILE._05286_ ),
    .X(\u_cpu.REG_FILE._05298_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10711_  (.A0(\u_cpu.REG_FILE.rf[20][10] ),
    .A1(\u_cpu.REG_FILE._05239_ ),
    .S(\u_cpu.REG_FILE._05298_ ),
    .X(\u_cpu.REG_FILE._05299_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10712_  (.A(\u_cpu.REG_FILE._05299_ ),
    .X(\u_cpu.REG_FILE._00682_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10713_  (.A0(\u_cpu.REG_FILE.rf[20][11] ),
    .A1(\u_cpu.REG_FILE._05242_ ),
    .S(\u_cpu.REG_FILE._05298_ ),
    .X(\u_cpu.REG_FILE._05300_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10714_  (.A(\u_cpu.REG_FILE._05300_ ),
    .X(\u_cpu.REG_FILE._00683_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10715_  (.A0(\u_cpu.REG_FILE.rf[20][12] ),
    .A1(\u_cpu.REG_FILE._05244_ ),
    .S(\u_cpu.REG_FILE._05298_ ),
    .X(\u_cpu.REG_FILE._05301_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10716_  (.A(\u_cpu.REG_FILE._05301_ ),
    .X(\u_cpu.REG_FILE._00684_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10717_  (.A0(\u_cpu.REG_FILE.rf[20][13] ),
    .A1(\u_cpu.REG_FILE._05246_ ),
    .S(\u_cpu.REG_FILE._05298_ ),
    .X(\u_cpu.REG_FILE._05302_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10718_  (.A(\u_cpu.REG_FILE._05302_ ),
    .X(\u_cpu.REG_FILE._00685_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10719_  (.A0(\u_cpu.REG_FILE.rf[20][14] ),
    .A1(\u_cpu.REG_FILE._05248_ ),
    .S(\u_cpu.REG_FILE._05298_ ),
    .X(\u_cpu.REG_FILE._05303_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10720_  (.A(\u_cpu.REG_FILE._05303_ ),
    .X(\u_cpu.REG_FILE._00686_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10721_  (.A0(\u_cpu.REG_FILE.rf[20][15] ),
    .A1(\u_cpu.REG_FILE._05250_ ),
    .S(\u_cpu.REG_FILE._05298_ ),
    .X(\u_cpu.REG_FILE._05304_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10722_  (.A(\u_cpu.REG_FILE._05304_ ),
    .X(\u_cpu.REG_FILE._00687_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10723_  (.A0(\u_cpu.REG_FILE.rf[20][16] ),
    .A1(\u_cpu.REG_FILE._05252_ ),
    .S(\u_cpu.REG_FILE._05298_ ),
    .X(\u_cpu.REG_FILE._05305_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10724_  (.A(\u_cpu.REG_FILE._05305_ ),
    .X(\u_cpu.REG_FILE._00688_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10725_  (.A0(\u_cpu.REG_FILE.rf[20][17] ),
    .A1(\u_cpu.REG_FILE._05254_ ),
    .S(\u_cpu.REG_FILE._05298_ ),
    .X(\u_cpu.REG_FILE._05306_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10726_  (.A(\u_cpu.REG_FILE._05306_ ),
    .X(\u_cpu.REG_FILE._00689_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10727_  (.A0(\u_cpu.REG_FILE.rf[20][18] ),
    .A1(\u_cpu.REG_FILE._05256_ ),
    .S(\u_cpu.REG_FILE._05298_ ),
    .X(\u_cpu.REG_FILE._05307_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10728_  (.A(\u_cpu.REG_FILE._05307_ ),
    .X(\u_cpu.REG_FILE._00690_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10729_  (.A0(\u_cpu.REG_FILE.rf[20][19] ),
    .A1(\u_cpu.REG_FILE._05258_ ),
    .S(\u_cpu.REG_FILE._05298_ ),
    .X(\u_cpu.REG_FILE._05308_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10730_  (.A(\u_cpu.REG_FILE._05308_ ),
    .X(\u_cpu.REG_FILE._00691_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10731_  (.A(\u_cpu.REG_FILE._05286_ ),
    .X(\u_cpu.REG_FILE._05309_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10732_  (.A0(\u_cpu.REG_FILE.rf[20][20] ),
    .A1(\u_cpu.REG_FILE._05260_ ),
    .S(\u_cpu.REG_FILE._05309_ ),
    .X(\u_cpu.REG_FILE._05310_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10733_  (.A(\u_cpu.REG_FILE._05310_ ),
    .X(\u_cpu.REG_FILE._00692_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10734_  (.A0(\u_cpu.REG_FILE.rf[20][21] ),
    .A1(\u_cpu.REG_FILE._05263_ ),
    .S(\u_cpu.REG_FILE._05309_ ),
    .X(\u_cpu.REG_FILE._05311_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10735_  (.A(\u_cpu.REG_FILE._05311_ ),
    .X(\u_cpu.REG_FILE._00693_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10736_  (.A0(\u_cpu.REG_FILE.rf[20][22] ),
    .A1(\u_cpu.REG_FILE._05265_ ),
    .S(\u_cpu.REG_FILE._05309_ ),
    .X(\u_cpu.REG_FILE._05312_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10737_  (.A(\u_cpu.REG_FILE._05312_ ),
    .X(\u_cpu.REG_FILE._00694_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10738_  (.A0(\u_cpu.REG_FILE.rf[20][23] ),
    .A1(\u_cpu.REG_FILE._05267_ ),
    .S(\u_cpu.REG_FILE._05309_ ),
    .X(\u_cpu.REG_FILE._05313_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10739_  (.A(\u_cpu.REG_FILE._05313_ ),
    .X(\u_cpu.REG_FILE._00695_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10740_  (.A0(\u_cpu.REG_FILE.rf[20][24] ),
    .A1(\u_cpu.REG_FILE._05269_ ),
    .S(\u_cpu.REG_FILE._05309_ ),
    .X(\u_cpu.REG_FILE._05314_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10741_  (.A(\u_cpu.REG_FILE._05314_ ),
    .X(\u_cpu.REG_FILE._00696_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10742_  (.A0(\u_cpu.REG_FILE.rf[20][25] ),
    .A1(\u_cpu.REG_FILE._05271_ ),
    .S(\u_cpu.REG_FILE._05309_ ),
    .X(\u_cpu.REG_FILE._05315_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10743_  (.A(\u_cpu.REG_FILE._05315_ ),
    .X(\u_cpu.REG_FILE._00697_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10744_  (.A0(\u_cpu.REG_FILE.rf[20][26] ),
    .A1(\u_cpu.REG_FILE._05273_ ),
    .S(\u_cpu.REG_FILE._05309_ ),
    .X(\u_cpu.REG_FILE._05316_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10745_  (.A(\u_cpu.REG_FILE._05316_ ),
    .X(\u_cpu.REG_FILE._00698_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10746_  (.A0(\u_cpu.REG_FILE.rf[20][27] ),
    .A1(\u_cpu.REG_FILE._05275_ ),
    .S(\u_cpu.REG_FILE._05309_ ),
    .X(\u_cpu.REG_FILE._05317_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10747_  (.A(\u_cpu.REG_FILE._05317_ ),
    .X(\u_cpu.REG_FILE._00699_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10748_  (.A0(\u_cpu.REG_FILE.rf[20][28] ),
    .A1(\u_cpu.REG_FILE._05277_ ),
    .S(\u_cpu.REG_FILE._05309_ ),
    .X(\u_cpu.REG_FILE._05318_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10749_  (.A(\u_cpu.REG_FILE._05318_ ),
    .X(\u_cpu.REG_FILE._00700_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10750_  (.A0(\u_cpu.REG_FILE.rf[20][29] ),
    .A1(\u_cpu.REG_FILE._05279_ ),
    .S(\u_cpu.REG_FILE._05309_ ),
    .X(\u_cpu.REG_FILE._05319_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10751_  (.A(\u_cpu.REG_FILE._05319_ ),
    .X(\u_cpu.REG_FILE._00701_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10752_  (.A0(\u_cpu.REG_FILE.rf[20][30] ),
    .A1(\u_cpu.REG_FILE._05281_ ),
    .S(\u_cpu.REG_FILE._05286_ ),
    .X(\u_cpu.REG_FILE._05320_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10753_  (.A(\u_cpu.REG_FILE._05320_ ),
    .X(\u_cpu.REG_FILE._00702_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10754_  (.A0(\u_cpu.REG_FILE.rf[20][31] ),
    .A1(\u_cpu.REG_FILE._05283_ ),
    .S(\u_cpu.REG_FILE._05286_ ),
    .X(\u_cpu.REG_FILE._05321_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10755_  (.A(\u_cpu.REG_FILE._05321_ ),
    .X(\u_cpu.REG_FILE._00703_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.REG_FILE._10756_  (.A_N(\u_cpu.REG_FILE._04421_ ),
    .B(\u_cpu.REG_FILE._04425_ ),
    .C(\u_cpu.REG_FILE._04423_ ),
    .D(\u_cpu.REG_FILE.a3[4] ),
    .X(\u_cpu.REG_FILE._05322_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10757_  (.A(\u_cpu.REG_FILE._05322_ ),
    .X(\u_cpu.REG_FILE._05323_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10758_  (.A(\u_cpu.REG_FILE._05323_ ),
    .X(\u_cpu.REG_FILE._05324_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10759_  (.A0(\u_cpu.REG_FILE.rf[21][0] ),
    .A1(\u_cpu.REG_FILE._05216_ ),
    .S(\u_cpu.REG_FILE._05324_ ),
    .X(\u_cpu.REG_FILE._05325_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10760_  (.A(\u_cpu.REG_FILE._05325_ ),
    .X(\u_cpu.REG_FILE._00704_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10761_  (.A0(\u_cpu.REG_FILE.rf[21][1] ),
    .A1(\u_cpu.REG_FILE._05221_ ),
    .S(\u_cpu.REG_FILE._05324_ ),
    .X(\u_cpu.REG_FILE._05326_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10762_  (.A(\u_cpu.REG_FILE._05326_ ),
    .X(\u_cpu.REG_FILE._00705_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10763_  (.A0(\u_cpu.REG_FILE.rf[21][2] ),
    .A1(\u_cpu.REG_FILE._05223_ ),
    .S(\u_cpu.REG_FILE._05324_ ),
    .X(\u_cpu.REG_FILE._05327_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10764_  (.A(\u_cpu.REG_FILE._05327_ ),
    .X(\u_cpu.REG_FILE._00706_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10765_  (.A0(\u_cpu.REG_FILE.rf[21][3] ),
    .A1(\u_cpu.REG_FILE._05225_ ),
    .S(\u_cpu.REG_FILE._05324_ ),
    .X(\u_cpu.REG_FILE._05328_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10766_  (.A(\u_cpu.REG_FILE._05328_ ),
    .X(\u_cpu.REG_FILE._00707_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10767_  (.A0(\u_cpu.REG_FILE.rf[21][4] ),
    .A1(\u_cpu.REG_FILE._05227_ ),
    .S(\u_cpu.REG_FILE._05324_ ),
    .X(\u_cpu.REG_FILE._05329_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10768_  (.A(\u_cpu.REG_FILE._05329_ ),
    .X(\u_cpu.REG_FILE._00708_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10769_  (.A0(\u_cpu.REG_FILE.rf[21][5] ),
    .A1(\u_cpu.REG_FILE._05229_ ),
    .S(\u_cpu.REG_FILE._05324_ ),
    .X(\u_cpu.REG_FILE._05330_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10770_  (.A(\u_cpu.REG_FILE._05330_ ),
    .X(\u_cpu.REG_FILE._00709_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10771_  (.A0(\u_cpu.REG_FILE.rf[21][6] ),
    .A1(\u_cpu.REG_FILE._05231_ ),
    .S(\u_cpu.REG_FILE._05324_ ),
    .X(\u_cpu.REG_FILE._05331_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10772_  (.A(\u_cpu.REG_FILE._05331_ ),
    .X(\u_cpu.REG_FILE._00710_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10773_  (.A0(\u_cpu.REG_FILE.rf[21][7] ),
    .A1(\u_cpu.REG_FILE._05233_ ),
    .S(\u_cpu.REG_FILE._05324_ ),
    .X(\u_cpu.REG_FILE._05332_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10774_  (.A(\u_cpu.REG_FILE._05332_ ),
    .X(\u_cpu.REG_FILE._00711_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10775_  (.A0(\u_cpu.REG_FILE.rf[21][8] ),
    .A1(\u_cpu.REG_FILE._05235_ ),
    .S(\u_cpu.REG_FILE._05324_ ),
    .X(\u_cpu.REG_FILE._05333_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10776_  (.A(\u_cpu.REG_FILE._05333_ ),
    .X(\u_cpu.REG_FILE._00712_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10777_  (.A0(\u_cpu.REG_FILE.rf[21][9] ),
    .A1(\u_cpu.REG_FILE._05237_ ),
    .S(\u_cpu.REG_FILE._05324_ ),
    .X(\u_cpu.REG_FILE._05334_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10778_  (.A(\u_cpu.REG_FILE._05334_ ),
    .X(\u_cpu.REG_FILE._00713_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10779_  (.A(\u_cpu.REG_FILE._05323_ ),
    .X(\u_cpu.REG_FILE._05335_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10780_  (.A0(\u_cpu.REG_FILE.rf[21][10] ),
    .A1(\u_cpu.REG_FILE._05239_ ),
    .S(\u_cpu.REG_FILE._05335_ ),
    .X(\u_cpu.REG_FILE._05336_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10781_  (.A(\u_cpu.REG_FILE._05336_ ),
    .X(\u_cpu.REG_FILE._00714_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10782_  (.A0(\u_cpu.REG_FILE.rf[21][11] ),
    .A1(\u_cpu.REG_FILE._05242_ ),
    .S(\u_cpu.REG_FILE._05335_ ),
    .X(\u_cpu.REG_FILE._05337_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10783_  (.A(\u_cpu.REG_FILE._05337_ ),
    .X(\u_cpu.REG_FILE._00715_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10784_  (.A0(\u_cpu.REG_FILE.rf[21][12] ),
    .A1(\u_cpu.REG_FILE._05244_ ),
    .S(\u_cpu.REG_FILE._05335_ ),
    .X(\u_cpu.REG_FILE._05338_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10785_  (.A(\u_cpu.REG_FILE._05338_ ),
    .X(\u_cpu.REG_FILE._00716_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10786_  (.A0(\u_cpu.REG_FILE.rf[21][13] ),
    .A1(\u_cpu.REG_FILE._05246_ ),
    .S(\u_cpu.REG_FILE._05335_ ),
    .X(\u_cpu.REG_FILE._05339_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10787_  (.A(\u_cpu.REG_FILE._05339_ ),
    .X(\u_cpu.REG_FILE._00717_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10788_  (.A0(\u_cpu.REG_FILE.rf[21][14] ),
    .A1(\u_cpu.REG_FILE._05248_ ),
    .S(\u_cpu.REG_FILE._05335_ ),
    .X(\u_cpu.REG_FILE._05340_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10789_  (.A(\u_cpu.REG_FILE._05340_ ),
    .X(\u_cpu.REG_FILE._00718_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10790_  (.A0(\u_cpu.REG_FILE.rf[21][15] ),
    .A1(\u_cpu.REG_FILE._05250_ ),
    .S(\u_cpu.REG_FILE._05335_ ),
    .X(\u_cpu.REG_FILE._05341_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10791_  (.A(\u_cpu.REG_FILE._05341_ ),
    .X(\u_cpu.REG_FILE._00719_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10792_  (.A0(\u_cpu.REG_FILE.rf[21][16] ),
    .A1(\u_cpu.REG_FILE._05252_ ),
    .S(\u_cpu.REG_FILE._05335_ ),
    .X(\u_cpu.REG_FILE._05342_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10793_  (.A(\u_cpu.REG_FILE._05342_ ),
    .X(\u_cpu.REG_FILE._00720_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10794_  (.A0(\u_cpu.REG_FILE.rf[21][17] ),
    .A1(\u_cpu.REG_FILE._05254_ ),
    .S(\u_cpu.REG_FILE._05335_ ),
    .X(\u_cpu.REG_FILE._05343_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10795_  (.A(\u_cpu.REG_FILE._05343_ ),
    .X(\u_cpu.REG_FILE._00721_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10796_  (.A0(\u_cpu.REG_FILE.rf[21][18] ),
    .A1(\u_cpu.REG_FILE._05256_ ),
    .S(\u_cpu.REG_FILE._05335_ ),
    .X(\u_cpu.REG_FILE._05344_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10797_  (.A(\u_cpu.REG_FILE._05344_ ),
    .X(\u_cpu.REG_FILE._00722_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10798_  (.A0(\u_cpu.REG_FILE.rf[21][19] ),
    .A1(\u_cpu.REG_FILE._05258_ ),
    .S(\u_cpu.REG_FILE._05335_ ),
    .X(\u_cpu.REG_FILE._05345_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10799_  (.A(\u_cpu.REG_FILE._05345_ ),
    .X(\u_cpu.REG_FILE._00723_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10800_  (.A(\u_cpu.REG_FILE._05323_ ),
    .X(\u_cpu.REG_FILE._05346_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10801_  (.A0(\u_cpu.REG_FILE.rf[21][20] ),
    .A1(\u_cpu.REG_FILE._05260_ ),
    .S(\u_cpu.REG_FILE._05346_ ),
    .X(\u_cpu.REG_FILE._05347_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10802_  (.A(\u_cpu.REG_FILE._05347_ ),
    .X(\u_cpu.REG_FILE._00724_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10803_  (.A0(\u_cpu.REG_FILE.rf[21][21] ),
    .A1(\u_cpu.REG_FILE._05263_ ),
    .S(\u_cpu.REG_FILE._05346_ ),
    .X(\u_cpu.REG_FILE._05348_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10804_  (.A(\u_cpu.REG_FILE._05348_ ),
    .X(\u_cpu.REG_FILE._00725_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10805_  (.A0(\u_cpu.REG_FILE.rf[21][22] ),
    .A1(\u_cpu.REG_FILE._05265_ ),
    .S(\u_cpu.REG_FILE._05346_ ),
    .X(\u_cpu.REG_FILE._05349_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10806_  (.A(\u_cpu.REG_FILE._05349_ ),
    .X(\u_cpu.REG_FILE._00726_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10807_  (.A0(\u_cpu.REG_FILE.rf[21][23] ),
    .A1(\u_cpu.REG_FILE._05267_ ),
    .S(\u_cpu.REG_FILE._05346_ ),
    .X(\u_cpu.REG_FILE._05350_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10808_  (.A(\u_cpu.REG_FILE._05350_ ),
    .X(\u_cpu.REG_FILE._00727_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10809_  (.A0(\u_cpu.REG_FILE.rf[21][24] ),
    .A1(\u_cpu.REG_FILE._05269_ ),
    .S(\u_cpu.REG_FILE._05346_ ),
    .X(\u_cpu.REG_FILE._05351_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10810_  (.A(\u_cpu.REG_FILE._05351_ ),
    .X(\u_cpu.REG_FILE._00728_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10811_  (.A0(\u_cpu.REG_FILE.rf[21][25] ),
    .A1(\u_cpu.REG_FILE._05271_ ),
    .S(\u_cpu.REG_FILE._05346_ ),
    .X(\u_cpu.REG_FILE._05352_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10812_  (.A(\u_cpu.REG_FILE._05352_ ),
    .X(\u_cpu.REG_FILE._00729_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10813_  (.A0(\u_cpu.REG_FILE.rf[21][26] ),
    .A1(\u_cpu.REG_FILE._05273_ ),
    .S(\u_cpu.REG_FILE._05346_ ),
    .X(\u_cpu.REG_FILE._05353_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10814_  (.A(\u_cpu.REG_FILE._05353_ ),
    .X(\u_cpu.REG_FILE._00730_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10815_  (.A0(\u_cpu.REG_FILE.rf[21][27] ),
    .A1(\u_cpu.REG_FILE._05275_ ),
    .S(\u_cpu.REG_FILE._05346_ ),
    .X(\u_cpu.REG_FILE._05354_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10816_  (.A(\u_cpu.REG_FILE._05354_ ),
    .X(\u_cpu.REG_FILE._00731_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10817_  (.A0(\u_cpu.REG_FILE.rf[21][28] ),
    .A1(\u_cpu.REG_FILE._05277_ ),
    .S(\u_cpu.REG_FILE._05346_ ),
    .X(\u_cpu.REG_FILE._05355_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10818_  (.A(\u_cpu.REG_FILE._05355_ ),
    .X(\u_cpu.REG_FILE._00732_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10819_  (.A0(\u_cpu.REG_FILE.rf[21][29] ),
    .A1(\u_cpu.REG_FILE._05279_ ),
    .S(\u_cpu.REG_FILE._05346_ ),
    .X(\u_cpu.REG_FILE._05356_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10820_  (.A(\u_cpu.REG_FILE._05356_ ),
    .X(\u_cpu.REG_FILE._00733_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10821_  (.A0(\u_cpu.REG_FILE.rf[21][30] ),
    .A1(\u_cpu.REG_FILE._05281_ ),
    .S(\u_cpu.REG_FILE._05323_ ),
    .X(\u_cpu.REG_FILE._05357_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10822_  (.A(\u_cpu.REG_FILE._05357_ ),
    .X(\u_cpu.REG_FILE._00734_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10823_  (.A0(\u_cpu.REG_FILE.rf[21][31] ),
    .A1(\u_cpu.REG_FILE._05283_ ),
    .S(\u_cpu.REG_FILE._05323_ ),
    .X(\u_cpu.REG_FILE._05358_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10824_  (.A(\u_cpu.REG_FILE._05358_ ),
    .X(\u_cpu.REG_FILE._00735_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.REG_FILE._10825_  (.A_N(\u_cpu.REG_FILE._04421_ ),
    .B(\u_cpu.REG_FILE._04425_ ),
    .C(\u_cpu.REG_FILE._04747_ ),
    .D(\u_cpu.REG_FILE.a3[4] ),
    .X(\u_cpu.REG_FILE._05359_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10826_  (.A(\u_cpu.REG_FILE._05359_ ),
    .X(\u_cpu.REG_FILE._05360_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10827_  (.A(\u_cpu.REG_FILE._05360_ ),
    .X(\u_cpu.REG_FILE._05361_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10828_  (.A0(\u_cpu.REG_FILE.rf[22][0] ),
    .A1(\u_cpu.REG_FILE._05216_ ),
    .S(\u_cpu.REG_FILE._05361_ ),
    .X(\u_cpu.REG_FILE._05362_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10829_  (.A(\u_cpu.REG_FILE._05362_ ),
    .X(\u_cpu.REG_FILE._00736_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10830_  (.A0(\u_cpu.REG_FILE.rf[22][1] ),
    .A1(\u_cpu.REG_FILE._05221_ ),
    .S(\u_cpu.REG_FILE._05361_ ),
    .X(\u_cpu.REG_FILE._05363_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10831_  (.A(\u_cpu.REG_FILE._05363_ ),
    .X(\u_cpu.REG_FILE._00737_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10832_  (.A0(\u_cpu.REG_FILE.rf[22][2] ),
    .A1(\u_cpu.REG_FILE._05223_ ),
    .S(\u_cpu.REG_FILE._05361_ ),
    .X(\u_cpu.REG_FILE._05364_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10833_  (.A(\u_cpu.REG_FILE._05364_ ),
    .X(\u_cpu.REG_FILE._00738_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10834_  (.A0(\u_cpu.REG_FILE.rf[22][3] ),
    .A1(\u_cpu.REG_FILE._05225_ ),
    .S(\u_cpu.REG_FILE._05361_ ),
    .X(\u_cpu.REG_FILE._05365_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10835_  (.A(\u_cpu.REG_FILE._05365_ ),
    .X(\u_cpu.REG_FILE._00739_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10836_  (.A0(\u_cpu.REG_FILE.rf[22][4] ),
    .A1(\u_cpu.REG_FILE._05227_ ),
    .S(\u_cpu.REG_FILE._05361_ ),
    .X(\u_cpu.REG_FILE._05366_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10837_  (.A(\u_cpu.REG_FILE._05366_ ),
    .X(\u_cpu.REG_FILE._00740_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10838_  (.A0(\u_cpu.REG_FILE.rf[22][5] ),
    .A1(\u_cpu.REG_FILE._05229_ ),
    .S(\u_cpu.REG_FILE._05361_ ),
    .X(\u_cpu.REG_FILE._05367_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10839_  (.A(\u_cpu.REG_FILE._05367_ ),
    .X(\u_cpu.REG_FILE._00741_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10840_  (.A0(\u_cpu.REG_FILE.rf[22][6] ),
    .A1(\u_cpu.REG_FILE._05231_ ),
    .S(\u_cpu.REG_FILE._05361_ ),
    .X(\u_cpu.REG_FILE._05368_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10841_  (.A(\u_cpu.REG_FILE._05368_ ),
    .X(\u_cpu.REG_FILE._00742_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10842_  (.A0(\u_cpu.REG_FILE.rf[22][7] ),
    .A1(\u_cpu.REG_FILE._05233_ ),
    .S(\u_cpu.REG_FILE._05361_ ),
    .X(\u_cpu.REG_FILE._05369_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10843_  (.A(\u_cpu.REG_FILE._05369_ ),
    .X(\u_cpu.REG_FILE._00743_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10844_  (.A0(\u_cpu.REG_FILE.rf[22][8] ),
    .A1(\u_cpu.REG_FILE._05235_ ),
    .S(\u_cpu.REG_FILE._05361_ ),
    .X(\u_cpu.REG_FILE._05370_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10845_  (.A(\u_cpu.REG_FILE._05370_ ),
    .X(\u_cpu.REG_FILE._00744_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10846_  (.A0(\u_cpu.REG_FILE.rf[22][9] ),
    .A1(\u_cpu.REG_FILE._05237_ ),
    .S(\u_cpu.REG_FILE._05361_ ),
    .X(\u_cpu.REG_FILE._05371_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10847_  (.A(\u_cpu.REG_FILE._05371_ ),
    .X(\u_cpu.REG_FILE._00745_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10848_  (.A(\u_cpu.REG_FILE._05360_ ),
    .X(\u_cpu.REG_FILE._05372_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10849_  (.A0(\u_cpu.REG_FILE.rf[22][10] ),
    .A1(\u_cpu.REG_FILE._05239_ ),
    .S(\u_cpu.REG_FILE._05372_ ),
    .X(\u_cpu.REG_FILE._05373_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10850_  (.A(\u_cpu.REG_FILE._05373_ ),
    .X(\u_cpu.REG_FILE._00746_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10851_  (.A0(\u_cpu.REG_FILE.rf[22][11] ),
    .A1(\u_cpu.REG_FILE._05242_ ),
    .S(\u_cpu.REG_FILE._05372_ ),
    .X(\u_cpu.REG_FILE._05374_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10852_  (.A(\u_cpu.REG_FILE._05374_ ),
    .X(\u_cpu.REG_FILE._00747_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10853_  (.A0(\u_cpu.REG_FILE.rf[22][12] ),
    .A1(\u_cpu.REG_FILE._05244_ ),
    .S(\u_cpu.REG_FILE._05372_ ),
    .X(\u_cpu.REG_FILE._05375_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10854_  (.A(\u_cpu.REG_FILE._05375_ ),
    .X(\u_cpu.REG_FILE._00748_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10855_  (.A0(\u_cpu.REG_FILE.rf[22][13] ),
    .A1(\u_cpu.REG_FILE._05246_ ),
    .S(\u_cpu.REG_FILE._05372_ ),
    .X(\u_cpu.REG_FILE._05376_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10856_  (.A(\u_cpu.REG_FILE._05376_ ),
    .X(\u_cpu.REG_FILE._00749_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10857_  (.A0(\u_cpu.REG_FILE.rf[22][14] ),
    .A1(\u_cpu.REG_FILE._05248_ ),
    .S(\u_cpu.REG_FILE._05372_ ),
    .X(\u_cpu.REG_FILE._05377_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10858_  (.A(\u_cpu.REG_FILE._05377_ ),
    .X(\u_cpu.REG_FILE._00750_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10859_  (.A0(\u_cpu.REG_FILE.rf[22][15] ),
    .A1(\u_cpu.REG_FILE._05250_ ),
    .S(\u_cpu.REG_FILE._05372_ ),
    .X(\u_cpu.REG_FILE._05378_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10860_  (.A(\u_cpu.REG_FILE._05378_ ),
    .X(\u_cpu.REG_FILE._00751_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10861_  (.A0(\u_cpu.REG_FILE.rf[22][16] ),
    .A1(\u_cpu.REG_FILE._05252_ ),
    .S(\u_cpu.REG_FILE._05372_ ),
    .X(\u_cpu.REG_FILE._05379_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10862_  (.A(\u_cpu.REG_FILE._05379_ ),
    .X(\u_cpu.REG_FILE._00752_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10863_  (.A0(\u_cpu.REG_FILE.rf[22][17] ),
    .A1(\u_cpu.REG_FILE._05254_ ),
    .S(\u_cpu.REG_FILE._05372_ ),
    .X(\u_cpu.REG_FILE._05380_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10864_  (.A(\u_cpu.REG_FILE._05380_ ),
    .X(\u_cpu.REG_FILE._00753_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10865_  (.A0(\u_cpu.REG_FILE.rf[22][18] ),
    .A1(\u_cpu.REG_FILE._05256_ ),
    .S(\u_cpu.REG_FILE._05372_ ),
    .X(\u_cpu.REG_FILE._05381_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10866_  (.A(\u_cpu.REG_FILE._05381_ ),
    .X(\u_cpu.REG_FILE._00754_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10867_  (.A0(\u_cpu.REG_FILE.rf[22][19] ),
    .A1(\u_cpu.REG_FILE._05258_ ),
    .S(\u_cpu.REG_FILE._05372_ ),
    .X(\u_cpu.REG_FILE._05382_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10868_  (.A(\u_cpu.REG_FILE._05382_ ),
    .X(\u_cpu.REG_FILE._00755_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10869_  (.A(\u_cpu.REG_FILE._05360_ ),
    .X(\u_cpu.REG_FILE._05383_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10870_  (.A0(\u_cpu.REG_FILE.rf[22][20] ),
    .A1(\u_cpu.REG_FILE._05260_ ),
    .S(\u_cpu.REG_FILE._05383_ ),
    .X(\u_cpu.REG_FILE._05384_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10871_  (.A(\u_cpu.REG_FILE._05384_ ),
    .X(\u_cpu.REG_FILE._00756_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10872_  (.A0(\u_cpu.REG_FILE.rf[22][21] ),
    .A1(\u_cpu.REG_FILE._05263_ ),
    .S(\u_cpu.REG_FILE._05383_ ),
    .X(\u_cpu.REG_FILE._05385_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10873_  (.A(\u_cpu.REG_FILE._05385_ ),
    .X(\u_cpu.REG_FILE._00757_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10874_  (.A0(\u_cpu.REG_FILE.rf[22][22] ),
    .A1(\u_cpu.REG_FILE._05265_ ),
    .S(\u_cpu.REG_FILE._05383_ ),
    .X(\u_cpu.REG_FILE._05386_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10875_  (.A(\u_cpu.REG_FILE._05386_ ),
    .X(\u_cpu.REG_FILE._00758_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10876_  (.A0(\u_cpu.REG_FILE.rf[22][23] ),
    .A1(\u_cpu.REG_FILE._05267_ ),
    .S(\u_cpu.REG_FILE._05383_ ),
    .X(\u_cpu.REG_FILE._05387_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10877_  (.A(\u_cpu.REG_FILE._05387_ ),
    .X(\u_cpu.REG_FILE._00759_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10878_  (.A0(\u_cpu.REG_FILE.rf[22][24] ),
    .A1(\u_cpu.REG_FILE._05269_ ),
    .S(\u_cpu.REG_FILE._05383_ ),
    .X(\u_cpu.REG_FILE._05388_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10879_  (.A(\u_cpu.REG_FILE._05388_ ),
    .X(\u_cpu.REG_FILE._00760_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10880_  (.A0(\u_cpu.REG_FILE.rf[22][25] ),
    .A1(\u_cpu.REG_FILE._05271_ ),
    .S(\u_cpu.REG_FILE._05383_ ),
    .X(\u_cpu.REG_FILE._05389_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10881_  (.A(\u_cpu.REG_FILE._05389_ ),
    .X(\u_cpu.REG_FILE._00761_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10882_  (.A0(\u_cpu.REG_FILE.rf[22][26] ),
    .A1(\u_cpu.REG_FILE._05273_ ),
    .S(\u_cpu.REG_FILE._05383_ ),
    .X(\u_cpu.REG_FILE._05390_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10883_  (.A(\u_cpu.REG_FILE._05390_ ),
    .X(\u_cpu.REG_FILE._00762_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10884_  (.A0(\u_cpu.REG_FILE.rf[22][27] ),
    .A1(\u_cpu.REG_FILE._05275_ ),
    .S(\u_cpu.REG_FILE._05383_ ),
    .X(\u_cpu.REG_FILE._05391_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10885_  (.A(\u_cpu.REG_FILE._05391_ ),
    .X(\u_cpu.REG_FILE._00763_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10886_  (.A0(\u_cpu.REG_FILE.rf[22][28] ),
    .A1(\u_cpu.REG_FILE._05277_ ),
    .S(\u_cpu.REG_FILE._05383_ ),
    .X(\u_cpu.REG_FILE._05392_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10887_  (.A(\u_cpu.REG_FILE._05392_ ),
    .X(\u_cpu.REG_FILE._00764_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10888_  (.A0(\u_cpu.REG_FILE.rf[22][29] ),
    .A1(\u_cpu.REG_FILE._05279_ ),
    .S(\u_cpu.REG_FILE._05383_ ),
    .X(\u_cpu.REG_FILE._05393_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10889_  (.A(\u_cpu.REG_FILE._05393_ ),
    .X(\u_cpu.REG_FILE._00765_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10890_  (.A0(\u_cpu.REG_FILE.rf[22][30] ),
    .A1(\u_cpu.REG_FILE._05281_ ),
    .S(\u_cpu.REG_FILE._05360_ ),
    .X(\u_cpu.REG_FILE._05394_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10891_  (.A(\u_cpu.REG_FILE._05394_ ),
    .X(\u_cpu.REG_FILE._00766_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10892_  (.A0(\u_cpu.REG_FILE.rf[22][31] ),
    .A1(\u_cpu.REG_FILE._05283_ ),
    .S(\u_cpu.REG_FILE._05360_ ),
    .X(\u_cpu.REG_FILE._05395_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10893_  (.A(\u_cpu.REG_FILE._05395_ ),
    .X(\u_cpu.REG_FILE._00767_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.REG_FILE._10894_  (.A_N(\u_cpu.REG_FILE._04421_ ),
    .B(\u_cpu.REG_FILE.a3[2] ),
    .C(\u_cpu.REG_FILE._04495_ ),
    .D(\u_cpu.REG_FILE.a3[4] ),
    .X(\u_cpu.REG_FILE._05396_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10895_  (.A(\u_cpu.REG_FILE._05396_ ),
    .X(\u_cpu.REG_FILE._05397_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10896_  (.A(\u_cpu.REG_FILE._05397_ ),
    .X(\u_cpu.REG_FILE._05398_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10897_  (.A0(\u_cpu.REG_FILE.rf[23][0] ),
    .A1(\u_cpu.REG_FILE._05216_ ),
    .S(\u_cpu.REG_FILE._05398_ ),
    .X(\u_cpu.REG_FILE._05399_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10898_  (.A(\u_cpu.REG_FILE._05399_ ),
    .X(\u_cpu.REG_FILE._00768_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10899_  (.A0(\u_cpu.REG_FILE.rf[23][1] ),
    .A1(\u_cpu.REG_FILE._05221_ ),
    .S(\u_cpu.REG_FILE._05398_ ),
    .X(\u_cpu.REG_FILE._05400_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10900_  (.A(\u_cpu.REG_FILE._05400_ ),
    .X(\u_cpu.REG_FILE._00769_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10901_  (.A0(\u_cpu.REG_FILE.rf[23][2] ),
    .A1(\u_cpu.REG_FILE._05223_ ),
    .S(\u_cpu.REG_FILE._05398_ ),
    .X(\u_cpu.REG_FILE._05401_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10902_  (.A(\u_cpu.REG_FILE._05401_ ),
    .X(\u_cpu.REG_FILE._00770_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10903_  (.A0(\u_cpu.REG_FILE.rf[23][3] ),
    .A1(\u_cpu.REG_FILE._05225_ ),
    .S(\u_cpu.REG_FILE._05398_ ),
    .X(\u_cpu.REG_FILE._05402_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10904_  (.A(\u_cpu.REG_FILE._05402_ ),
    .X(\u_cpu.REG_FILE._00771_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10905_  (.A0(\u_cpu.REG_FILE.rf[23][4] ),
    .A1(\u_cpu.REG_FILE._05227_ ),
    .S(\u_cpu.REG_FILE._05398_ ),
    .X(\u_cpu.REG_FILE._05403_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10906_  (.A(\u_cpu.REG_FILE._05403_ ),
    .X(\u_cpu.REG_FILE._00772_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10907_  (.A0(\u_cpu.REG_FILE.rf[23][5] ),
    .A1(\u_cpu.REG_FILE._05229_ ),
    .S(\u_cpu.REG_FILE._05398_ ),
    .X(\u_cpu.REG_FILE._05404_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10908_  (.A(\u_cpu.REG_FILE._05404_ ),
    .X(\u_cpu.REG_FILE._00773_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10909_  (.A0(\u_cpu.REG_FILE.rf[23][6] ),
    .A1(\u_cpu.REG_FILE._05231_ ),
    .S(\u_cpu.REG_FILE._05398_ ),
    .X(\u_cpu.REG_FILE._05405_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10910_  (.A(\u_cpu.REG_FILE._05405_ ),
    .X(\u_cpu.REG_FILE._00774_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10911_  (.A0(\u_cpu.REG_FILE.rf[23][7] ),
    .A1(\u_cpu.REG_FILE._05233_ ),
    .S(\u_cpu.REG_FILE._05398_ ),
    .X(\u_cpu.REG_FILE._05406_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10912_  (.A(\u_cpu.REG_FILE._05406_ ),
    .X(\u_cpu.REG_FILE._00775_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10913_  (.A0(\u_cpu.REG_FILE.rf[23][8] ),
    .A1(\u_cpu.REG_FILE._05235_ ),
    .S(\u_cpu.REG_FILE._05398_ ),
    .X(\u_cpu.REG_FILE._05407_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10914_  (.A(\u_cpu.REG_FILE._05407_ ),
    .X(\u_cpu.REG_FILE._00776_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10915_  (.A0(\u_cpu.REG_FILE.rf[23][9] ),
    .A1(\u_cpu.REG_FILE._05237_ ),
    .S(\u_cpu.REG_FILE._05398_ ),
    .X(\u_cpu.REG_FILE._05408_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10916_  (.A(\u_cpu.REG_FILE._05408_ ),
    .X(\u_cpu.REG_FILE._00777_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10917_  (.A(\u_cpu.REG_FILE._05397_ ),
    .X(\u_cpu.REG_FILE._05409_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10918_  (.A0(\u_cpu.REG_FILE.rf[23][10] ),
    .A1(\u_cpu.REG_FILE._05239_ ),
    .S(\u_cpu.REG_FILE._05409_ ),
    .X(\u_cpu.REG_FILE._05410_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10919_  (.A(\u_cpu.REG_FILE._05410_ ),
    .X(\u_cpu.REG_FILE._00778_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10920_  (.A0(\u_cpu.REG_FILE.rf[23][11] ),
    .A1(\u_cpu.REG_FILE._05242_ ),
    .S(\u_cpu.REG_FILE._05409_ ),
    .X(\u_cpu.REG_FILE._05411_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10921_  (.A(\u_cpu.REG_FILE._05411_ ),
    .X(\u_cpu.REG_FILE._00779_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10922_  (.A0(\u_cpu.REG_FILE.rf[23][12] ),
    .A1(\u_cpu.REG_FILE._05244_ ),
    .S(\u_cpu.REG_FILE._05409_ ),
    .X(\u_cpu.REG_FILE._05412_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10923_  (.A(\u_cpu.REG_FILE._05412_ ),
    .X(\u_cpu.REG_FILE._00780_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10924_  (.A0(\u_cpu.REG_FILE.rf[23][13] ),
    .A1(\u_cpu.REG_FILE._05246_ ),
    .S(\u_cpu.REG_FILE._05409_ ),
    .X(\u_cpu.REG_FILE._05413_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10925_  (.A(\u_cpu.REG_FILE._05413_ ),
    .X(\u_cpu.REG_FILE._00781_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10926_  (.A0(\u_cpu.REG_FILE.rf[23][14] ),
    .A1(\u_cpu.REG_FILE._05248_ ),
    .S(\u_cpu.REG_FILE._05409_ ),
    .X(\u_cpu.REG_FILE._05414_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10927_  (.A(\u_cpu.REG_FILE._05414_ ),
    .X(\u_cpu.REG_FILE._00782_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10928_  (.A0(\u_cpu.REG_FILE.rf[23][15] ),
    .A1(\u_cpu.REG_FILE._05250_ ),
    .S(\u_cpu.REG_FILE._05409_ ),
    .X(\u_cpu.REG_FILE._05415_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10929_  (.A(\u_cpu.REG_FILE._05415_ ),
    .X(\u_cpu.REG_FILE._00783_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10930_  (.A0(\u_cpu.REG_FILE.rf[23][16] ),
    .A1(\u_cpu.REG_FILE._05252_ ),
    .S(\u_cpu.REG_FILE._05409_ ),
    .X(\u_cpu.REG_FILE._05416_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10931_  (.A(\u_cpu.REG_FILE._05416_ ),
    .X(\u_cpu.REG_FILE._00784_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10932_  (.A0(\u_cpu.REG_FILE.rf[23][17] ),
    .A1(\u_cpu.REG_FILE._05254_ ),
    .S(\u_cpu.REG_FILE._05409_ ),
    .X(\u_cpu.REG_FILE._05417_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10933_  (.A(\u_cpu.REG_FILE._05417_ ),
    .X(\u_cpu.REG_FILE._00785_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10934_  (.A0(\u_cpu.REG_FILE.rf[23][18] ),
    .A1(\u_cpu.REG_FILE._05256_ ),
    .S(\u_cpu.REG_FILE._05409_ ),
    .X(\u_cpu.REG_FILE._05418_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10935_  (.A(\u_cpu.REG_FILE._05418_ ),
    .X(\u_cpu.REG_FILE._00786_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10936_  (.A0(\u_cpu.REG_FILE.rf[23][19] ),
    .A1(\u_cpu.REG_FILE._05258_ ),
    .S(\u_cpu.REG_FILE._05409_ ),
    .X(\u_cpu.REG_FILE._05419_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10937_  (.A(\u_cpu.REG_FILE._05419_ ),
    .X(\u_cpu.REG_FILE._00787_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10938_  (.A(\u_cpu.REG_FILE._05397_ ),
    .X(\u_cpu.REG_FILE._05420_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10939_  (.A0(\u_cpu.REG_FILE.rf[23][20] ),
    .A1(\u_cpu.REG_FILE._05260_ ),
    .S(\u_cpu.REG_FILE._05420_ ),
    .X(\u_cpu.REG_FILE._05421_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10940_  (.A(\u_cpu.REG_FILE._05421_ ),
    .X(\u_cpu.REG_FILE._00788_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10941_  (.A0(\u_cpu.REG_FILE.rf[23][21] ),
    .A1(\u_cpu.REG_FILE._05263_ ),
    .S(\u_cpu.REG_FILE._05420_ ),
    .X(\u_cpu.REG_FILE._05422_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10942_  (.A(\u_cpu.REG_FILE._05422_ ),
    .X(\u_cpu.REG_FILE._00789_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10943_  (.A0(\u_cpu.REG_FILE.rf[23][22] ),
    .A1(\u_cpu.REG_FILE._05265_ ),
    .S(\u_cpu.REG_FILE._05420_ ),
    .X(\u_cpu.REG_FILE._05423_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10944_  (.A(\u_cpu.REG_FILE._05423_ ),
    .X(\u_cpu.REG_FILE._00790_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10945_  (.A0(\u_cpu.REG_FILE.rf[23][23] ),
    .A1(\u_cpu.REG_FILE._05267_ ),
    .S(\u_cpu.REG_FILE._05420_ ),
    .X(\u_cpu.REG_FILE._05424_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10946_  (.A(\u_cpu.REG_FILE._05424_ ),
    .X(\u_cpu.REG_FILE._00791_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10947_  (.A0(\u_cpu.REG_FILE.rf[23][24] ),
    .A1(\u_cpu.REG_FILE._05269_ ),
    .S(\u_cpu.REG_FILE._05420_ ),
    .X(\u_cpu.REG_FILE._05425_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10948_  (.A(\u_cpu.REG_FILE._05425_ ),
    .X(\u_cpu.REG_FILE._00792_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10949_  (.A0(\u_cpu.REG_FILE.rf[23][25] ),
    .A1(\u_cpu.REG_FILE._05271_ ),
    .S(\u_cpu.REG_FILE._05420_ ),
    .X(\u_cpu.REG_FILE._05426_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10950_  (.A(\u_cpu.REG_FILE._05426_ ),
    .X(\u_cpu.REG_FILE._00793_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10951_  (.A0(\u_cpu.REG_FILE.rf[23][26] ),
    .A1(\u_cpu.REG_FILE._05273_ ),
    .S(\u_cpu.REG_FILE._05420_ ),
    .X(\u_cpu.REG_FILE._05427_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10952_  (.A(\u_cpu.REG_FILE._05427_ ),
    .X(\u_cpu.REG_FILE._00794_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10953_  (.A0(\u_cpu.REG_FILE.rf[23][27] ),
    .A1(\u_cpu.REG_FILE._05275_ ),
    .S(\u_cpu.REG_FILE._05420_ ),
    .X(\u_cpu.REG_FILE._05428_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10954_  (.A(\u_cpu.REG_FILE._05428_ ),
    .X(\u_cpu.REG_FILE._00795_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10955_  (.A0(\u_cpu.REG_FILE.rf[23][28] ),
    .A1(\u_cpu.REG_FILE._05277_ ),
    .S(\u_cpu.REG_FILE._05420_ ),
    .X(\u_cpu.REG_FILE._05429_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10956_  (.A(\u_cpu.REG_FILE._05429_ ),
    .X(\u_cpu.REG_FILE._00796_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10957_  (.A0(\u_cpu.REG_FILE.rf[23][29] ),
    .A1(\u_cpu.REG_FILE._05279_ ),
    .S(\u_cpu.REG_FILE._05420_ ),
    .X(\u_cpu.REG_FILE._05430_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10958_  (.A(\u_cpu.REG_FILE._05430_ ),
    .X(\u_cpu.REG_FILE._00797_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10959_  (.A0(\u_cpu.REG_FILE.rf[23][30] ),
    .A1(\u_cpu.REG_FILE._05281_ ),
    .S(\u_cpu.REG_FILE._05397_ ),
    .X(\u_cpu.REG_FILE._05431_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10960_  (.A(\u_cpu.REG_FILE._05431_ ),
    .X(\u_cpu.REG_FILE._00798_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10961_  (.A0(\u_cpu.REG_FILE.rf[23][31] ),
    .A1(\u_cpu.REG_FILE._05283_ ),
    .S(\u_cpu.REG_FILE._05397_ ),
    .X(\u_cpu.REG_FILE._05432_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10962_  (.A(\u_cpu.REG_FILE._05432_ ),
    .X(\u_cpu.REG_FILE._00799_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.REG_FILE._10963_  (.A_N(\u_cpu.REG_FILE._04425_ ),
    .B(\u_cpu.REG_FILE._04643_ ),
    .C(\u_cpu.REG_FILE._04424_ ),
    .D(\u_cpu.REG_FILE.a3[3] ),
    .X(\u_cpu.REG_FILE._05433_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10964_  (.A(\u_cpu.REG_FILE._05433_ ),
    .X(\u_cpu.REG_FILE._05434_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10965_  (.A(\u_cpu.REG_FILE._05434_ ),
    .X(\u_cpu.REG_FILE._05435_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10966_  (.A0(\u_cpu.REG_FILE.rf[24][0] ),
    .A1(\u_cpu.REG_FILE._05216_ ),
    .S(\u_cpu.REG_FILE._05435_ ),
    .X(\u_cpu.REG_FILE._05436_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10967_  (.A(\u_cpu.REG_FILE._05436_ ),
    .X(\u_cpu.REG_FILE._00800_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10968_  (.A0(\u_cpu.REG_FILE.rf[24][1] ),
    .A1(\u_cpu.REG_FILE._05221_ ),
    .S(\u_cpu.REG_FILE._05435_ ),
    .X(\u_cpu.REG_FILE._05437_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10969_  (.A(\u_cpu.REG_FILE._05437_ ),
    .X(\u_cpu.REG_FILE._00801_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10970_  (.A0(\u_cpu.REG_FILE.rf[24][2] ),
    .A1(\u_cpu.REG_FILE._05223_ ),
    .S(\u_cpu.REG_FILE._05435_ ),
    .X(\u_cpu.REG_FILE._05438_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10971_  (.A(\u_cpu.REG_FILE._05438_ ),
    .X(\u_cpu.REG_FILE._00802_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10972_  (.A0(\u_cpu.REG_FILE.rf[24][3] ),
    .A1(\u_cpu.REG_FILE._05225_ ),
    .S(\u_cpu.REG_FILE._05435_ ),
    .X(\u_cpu.REG_FILE._05439_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10973_  (.A(\u_cpu.REG_FILE._05439_ ),
    .X(\u_cpu.REG_FILE._00803_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10974_  (.A0(\u_cpu.REG_FILE.rf[24][4] ),
    .A1(\u_cpu.REG_FILE._05227_ ),
    .S(\u_cpu.REG_FILE._05435_ ),
    .X(\u_cpu.REG_FILE._05440_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10975_  (.A(\u_cpu.REG_FILE._05440_ ),
    .X(\u_cpu.REG_FILE._00804_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10976_  (.A0(\u_cpu.REG_FILE.rf[24][5] ),
    .A1(\u_cpu.REG_FILE._05229_ ),
    .S(\u_cpu.REG_FILE._05435_ ),
    .X(\u_cpu.REG_FILE._05441_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10977_  (.A(\u_cpu.REG_FILE._05441_ ),
    .X(\u_cpu.REG_FILE._00805_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10978_  (.A0(\u_cpu.REG_FILE.rf[24][6] ),
    .A1(\u_cpu.REG_FILE._05231_ ),
    .S(\u_cpu.REG_FILE._05435_ ),
    .X(\u_cpu.REG_FILE._05442_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10979_  (.A(\u_cpu.REG_FILE._05442_ ),
    .X(\u_cpu.REG_FILE._00806_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10980_  (.A0(\u_cpu.REG_FILE.rf[24][7] ),
    .A1(\u_cpu.REG_FILE._05233_ ),
    .S(\u_cpu.REG_FILE._05435_ ),
    .X(\u_cpu.REG_FILE._05443_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10981_  (.A(\u_cpu.REG_FILE._05443_ ),
    .X(\u_cpu.REG_FILE._00807_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10982_  (.A0(\u_cpu.REG_FILE.rf[24][8] ),
    .A1(\u_cpu.REG_FILE._05235_ ),
    .S(\u_cpu.REG_FILE._05435_ ),
    .X(\u_cpu.REG_FILE._05444_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10983_  (.A(\u_cpu.REG_FILE._05444_ ),
    .X(\u_cpu.REG_FILE._00808_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10984_  (.A0(\u_cpu.REG_FILE.rf[24][9] ),
    .A1(\u_cpu.REG_FILE._05237_ ),
    .S(\u_cpu.REG_FILE._05435_ ),
    .X(\u_cpu.REG_FILE._05445_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10985_  (.A(\u_cpu.REG_FILE._05445_ ),
    .X(\u_cpu.REG_FILE._00809_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10986_  (.A(\u_cpu.REG_FILE._05434_ ),
    .X(\u_cpu.REG_FILE._05446_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10987_  (.A0(\u_cpu.REG_FILE.rf[24][10] ),
    .A1(\u_cpu.REG_FILE._05239_ ),
    .S(\u_cpu.REG_FILE._05446_ ),
    .X(\u_cpu.REG_FILE._05447_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10988_  (.A(\u_cpu.REG_FILE._05447_ ),
    .X(\u_cpu.REG_FILE._00810_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10989_  (.A0(\u_cpu.REG_FILE.rf[24][11] ),
    .A1(\u_cpu.REG_FILE._05242_ ),
    .S(\u_cpu.REG_FILE._05446_ ),
    .X(\u_cpu.REG_FILE._05448_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10990_  (.A(\u_cpu.REG_FILE._05448_ ),
    .X(\u_cpu.REG_FILE._00811_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10991_  (.A0(\u_cpu.REG_FILE.rf[24][12] ),
    .A1(\u_cpu.REG_FILE._05244_ ),
    .S(\u_cpu.REG_FILE._05446_ ),
    .X(\u_cpu.REG_FILE._05449_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10992_  (.A(\u_cpu.REG_FILE._05449_ ),
    .X(\u_cpu.REG_FILE._00812_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10993_  (.A0(\u_cpu.REG_FILE.rf[24][13] ),
    .A1(\u_cpu.REG_FILE._05246_ ),
    .S(\u_cpu.REG_FILE._05446_ ),
    .X(\u_cpu.REG_FILE._05450_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10994_  (.A(\u_cpu.REG_FILE._05450_ ),
    .X(\u_cpu.REG_FILE._00813_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10995_  (.A0(\u_cpu.REG_FILE.rf[24][14] ),
    .A1(\u_cpu.REG_FILE._05248_ ),
    .S(\u_cpu.REG_FILE._05446_ ),
    .X(\u_cpu.REG_FILE._05451_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10996_  (.A(\u_cpu.REG_FILE._05451_ ),
    .X(\u_cpu.REG_FILE._00814_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10997_  (.A0(\u_cpu.REG_FILE.rf[24][15] ),
    .A1(\u_cpu.REG_FILE._05250_ ),
    .S(\u_cpu.REG_FILE._05446_ ),
    .X(\u_cpu.REG_FILE._05452_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._10998_  (.A(\u_cpu.REG_FILE._05452_ ),
    .X(\u_cpu.REG_FILE._00815_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._10999_  (.A0(\u_cpu.REG_FILE.rf[24][16] ),
    .A1(\u_cpu.REG_FILE._05252_ ),
    .S(\u_cpu.REG_FILE._05446_ ),
    .X(\u_cpu.REG_FILE._05453_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11000_  (.A(\u_cpu.REG_FILE._05453_ ),
    .X(\u_cpu.REG_FILE._00816_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11001_  (.A0(\u_cpu.REG_FILE.rf[24][17] ),
    .A1(\u_cpu.REG_FILE._05254_ ),
    .S(\u_cpu.REG_FILE._05446_ ),
    .X(\u_cpu.REG_FILE._05454_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11002_  (.A(\u_cpu.REG_FILE._05454_ ),
    .X(\u_cpu.REG_FILE._00817_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11003_  (.A0(\u_cpu.REG_FILE.rf[24][18] ),
    .A1(\u_cpu.REG_FILE._05256_ ),
    .S(\u_cpu.REG_FILE._05446_ ),
    .X(\u_cpu.REG_FILE._05455_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11004_  (.A(\u_cpu.REG_FILE._05455_ ),
    .X(\u_cpu.REG_FILE._00818_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11005_  (.A0(\u_cpu.REG_FILE.rf[24][19] ),
    .A1(\u_cpu.REG_FILE._05258_ ),
    .S(\u_cpu.REG_FILE._05446_ ),
    .X(\u_cpu.REG_FILE._05456_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11006_  (.A(\u_cpu.REG_FILE._05456_ ),
    .X(\u_cpu.REG_FILE._00819_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11007_  (.A(\u_cpu.REG_FILE._05434_ ),
    .X(\u_cpu.REG_FILE._05457_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11008_  (.A0(\u_cpu.REG_FILE.rf[24][20] ),
    .A1(\u_cpu.REG_FILE._05260_ ),
    .S(\u_cpu.REG_FILE._05457_ ),
    .X(\u_cpu.REG_FILE._05458_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11009_  (.A(\u_cpu.REG_FILE._05458_ ),
    .X(\u_cpu.REG_FILE._00820_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11010_  (.A0(\u_cpu.REG_FILE.rf[24][21] ),
    .A1(\u_cpu.REG_FILE._05263_ ),
    .S(\u_cpu.REG_FILE._05457_ ),
    .X(\u_cpu.REG_FILE._05459_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11011_  (.A(\u_cpu.REG_FILE._05459_ ),
    .X(\u_cpu.REG_FILE._00821_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11012_  (.A0(\u_cpu.REG_FILE.rf[24][22] ),
    .A1(\u_cpu.REG_FILE._05265_ ),
    .S(\u_cpu.REG_FILE._05457_ ),
    .X(\u_cpu.REG_FILE._05460_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11013_  (.A(\u_cpu.REG_FILE._05460_ ),
    .X(\u_cpu.REG_FILE._00822_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11014_  (.A0(\u_cpu.REG_FILE.rf[24][23] ),
    .A1(\u_cpu.REG_FILE._05267_ ),
    .S(\u_cpu.REG_FILE._05457_ ),
    .X(\u_cpu.REG_FILE._05461_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11015_  (.A(\u_cpu.REG_FILE._05461_ ),
    .X(\u_cpu.REG_FILE._00823_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11016_  (.A0(\u_cpu.REG_FILE.rf[24][24] ),
    .A1(\u_cpu.REG_FILE._05269_ ),
    .S(\u_cpu.REG_FILE._05457_ ),
    .X(\u_cpu.REG_FILE._05462_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11017_  (.A(\u_cpu.REG_FILE._05462_ ),
    .X(\u_cpu.REG_FILE._00824_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11018_  (.A0(\u_cpu.REG_FILE.rf[24][25] ),
    .A1(\u_cpu.REG_FILE._05271_ ),
    .S(\u_cpu.REG_FILE._05457_ ),
    .X(\u_cpu.REG_FILE._05463_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11019_  (.A(\u_cpu.REG_FILE._05463_ ),
    .X(\u_cpu.REG_FILE._00825_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11020_  (.A0(\u_cpu.REG_FILE.rf[24][26] ),
    .A1(\u_cpu.REG_FILE._05273_ ),
    .S(\u_cpu.REG_FILE._05457_ ),
    .X(\u_cpu.REG_FILE._05464_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11021_  (.A(\u_cpu.REG_FILE._05464_ ),
    .X(\u_cpu.REG_FILE._00826_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11022_  (.A0(\u_cpu.REG_FILE.rf[24][27] ),
    .A1(\u_cpu.REG_FILE._05275_ ),
    .S(\u_cpu.REG_FILE._05457_ ),
    .X(\u_cpu.REG_FILE._05465_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11023_  (.A(\u_cpu.REG_FILE._05465_ ),
    .X(\u_cpu.REG_FILE._00827_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11024_  (.A0(\u_cpu.REG_FILE.rf[24][28] ),
    .A1(\u_cpu.REG_FILE._05277_ ),
    .S(\u_cpu.REG_FILE._05457_ ),
    .X(\u_cpu.REG_FILE._05466_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11025_  (.A(\u_cpu.REG_FILE._05466_ ),
    .X(\u_cpu.REG_FILE._00828_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11026_  (.A0(\u_cpu.REG_FILE.rf[24][29] ),
    .A1(\u_cpu.REG_FILE._05279_ ),
    .S(\u_cpu.REG_FILE._05457_ ),
    .X(\u_cpu.REG_FILE._05467_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11027_  (.A(\u_cpu.REG_FILE._05467_ ),
    .X(\u_cpu.REG_FILE._00829_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11028_  (.A0(\u_cpu.REG_FILE.rf[24][30] ),
    .A1(\u_cpu.REG_FILE._05281_ ),
    .S(\u_cpu.REG_FILE._05434_ ),
    .X(\u_cpu.REG_FILE._05468_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11029_  (.A(\u_cpu.REG_FILE._05468_ ),
    .X(\u_cpu.REG_FILE._00830_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11030_  (.A0(\u_cpu.REG_FILE.rf[24][31] ),
    .A1(\u_cpu.REG_FILE._05283_ ),
    .S(\u_cpu.REG_FILE._05434_ ),
    .X(\u_cpu.REG_FILE._05469_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11031_  (.A(\u_cpu.REG_FILE._05469_ ),
    .X(\u_cpu.REG_FILE._00831_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.REG_FILE._11032_  (.A_N(\u_cpu.REG_FILE._04425_ ),
    .B(\u_cpu.REG_FILE._04423_ ),
    .C(\u_cpu.REG_FILE.a3[4] ),
    .D(\u_cpu.REG_FILE.a3[3] ),
    .X(\u_cpu.REG_FILE._05470_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11033_  (.A(\u_cpu.REG_FILE._05470_ ),
    .X(\u_cpu.REG_FILE._05471_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11034_  (.A(\u_cpu.REG_FILE._05471_ ),
    .X(\u_cpu.REG_FILE._05472_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11035_  (.A0(\u_cpu.REG_FILE.rf[25][0] ),
    .A1(\u_cpu.REG_FILE._05216_ ),
    .S(\u_cpu.REG_FILE._05472_ ),
    .X(\u_cpu.REG_FILE._05473_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11036_  (.A(\u_cpu.REG_FILE._05473_ ),
    .X(\u_cpu.REG_FILE._00832_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11037_  (.A0(\u_cpu.REG_FILE.rf[25][1] ),
    .A1(\u_cpu.REG_FILE._05221_ ),
    .S(\u_cpu.REG_FILE._05472_ ),
    .X(\u_cpu.REG_FILE._05474_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11038_  (.A(\u_cpu.REG_FILE._05474_ ),
    .X(\u_cpu.REG_FILE._00833_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11039_  (.A0(\u_cpu.REG_FILE.rf[25][2] ),
    .A1(\u_cpu.REG_FILE._05223_ ),
    .S(\u_cpu.REG_FILE._05472_ ),
    .X(\u_cpu.REG_FILE._05475_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11040_  (.A(\u_cpu.REG_FILE._05475_ ),
    .X(\u_cpu.REG_FILE._00834_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11041_  (.A0(\u_cpu.REG_FILE.rf[25][3] ),
    .A1(\u_cpu.REG_FILE._05225_ ),
    .S(\u_cpu.REG_FILE._05472_ ),
    .X(\u_cpu.REG_FILE._05476_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11042_  (.A(\u_cpu.REG_FILE._05476_ ),
    .X(\u_cpu.REG_FILE._00835_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11043_  (.A0(\u_cpu.REG_FILE.rf[25][4] ),
    .A1(\u_cpu.REG_FILE._05227_ ),
    .S(\u_cpu.REG_FILE._05472_ ),
    .X(\u_cpu.REG_FILE._05477_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11044_  (.A(\u_cpu.REG_FILE._05477_ ),
    .X(\u_cpu.REG_FILE._00836_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11045_  (.A0(\u_cpu.REG_FILE.rf[25][5] ),
    .A1(\u_cpu.REG_FILE._05229_ ),
    .S(\u_cpu.REG_FILE._05472_ ),
    .X(\u_cpu.REG_FILE._05478_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11046_  (.A(\u_cpu.REG_FILE._05478_ ),
    .X(\u_cpu.REG_FILE._00837_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11047_  (.A0(\u_cpu.REG_FILE.rf[25][6] ),
    .A1(\u_cpu.REG_FILE._05231_ ),
    .S(\u_cpu.REG_FILE._05472_ ),
    .X(\u_cpu.REG_FILE._05479_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11048_  (.A(\u_cpu.REG_FILE._05479_ ),
    .X(\u_cpu.REG_FILE._00838_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11049_  (.A0(\u_cpu.REG_FILE.rf[25][7] ),
    .A1(\u_cpu.REG_FILE._05233_ ),
    .S(\u_cpu.REG_FILE._05472_ ),
    .X(\u_cpu.REG_FILE._05480_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11050_  (.A(\u_cpu.REG_FILE._05480_ ),
    .X(\u_cpu.REG_FILE._00839_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11051_  (.A0(\u_cpu.REG_FILE.rf[25][8] ),
    .A1(\u_cpu.REG_FILE._05235_ ),
    .S(\u_cpu.REG_FILE._05472_ ),
    .X(\u_cpu.REG_FILE._05481_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11052_  (.A(\u_cpu.REG_FILE._05481_ ),
    .X(\u_cpu.REG_FILE._00840_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11053_  (.A0(\u_cpu.REG_FILE.rf[25][9] ),
    .A1(\u_cpu.REG_FILE._05237_ ),
    .S(\u_cpu.REG_FILE._05472_ ),
    .X(\u_cpu.REG_FILE._05482_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11054_  (.A(\u_cpu.REG_FILE._05482_ ),
    .X(\u_cpu.REG_FILE._00841_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11055_  (.A(\u_cpu.REG_FILE._05471_ ),
    .X(\u_cpu.REG_FILE._05483_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11056_  (.A0(\u_cpu.REG_FILE.rf[25][10] ),
    .A1(\u_cpu.REG_FILE._05239_ ),
    .S(\u_cpu.REG_FILE._05483_ ),
    .X(\u_cpu.REG_FILE._05484_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11057_  (.A(\u_cpu.REG_FILE._05484_ ),
    .X(\u_cpu.REG_FILE._00842_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11058_  (.A0(\u_cpu.REG_FILE.rf[25][11] ),
    .A1(\u_cpu.REG_FILE._05242_ ),
    .S(\u_cpu.REG_FILE._05483_ ),
    .X(\u_cpu.REG_FILE._05485_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11059_  (.A(\u_cpu.REG_FILE._05485_ ),
    .X(\u_cpu.REG_FILE._00843_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11060_  (.A0(\u_cpu.REG_FILE.rf[25][12] ),
    .A1(\u_cpu.REG_FILE._05244_ ),
    .S(\u_cpu.REG_FILE._05483_ ),
    .X(\u_cpu.REG_FILE._05486_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11061_  (.A(\u_cpu.REG_FILE._05486_ ),
    .X(\u_cpu.REG_FILE._00844_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11062_  (.A0(\u_cpu.REG_FILE.rf[25][13] ),
    .A1(\u_cpu.REG_FILE._05246_ ),
    .S(\u_cpu.REG_FILE._05483_ ),
    .X(\u_cpu.REG_FILE._05487_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11063_  (.A(\u_cpu.REG_FILE._05487_ ),
    .X(\u_cpu.REG_FILE._00845_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11064_  (.A0(\u_cpu.REG_FILE.rf[25][14] ),
    .A1(\u_cpu.REG_FILE._05248_ ),
    .S(\u_cpu.REG_FILE._05483_ ),
    .X(\u_cpu.REG_FILE._05488_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11065_  (.A(\u_cpu.REG_FILE._05488_ ),
    .X(\u_cpu.REG_FILE._00846_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11066_  (.A0(\u_cpu.REG_FILE.rf[25][15] ),
    .A1(\u_cpu.REG_FILE._05250_ ),
    .S(\u_cpu.REG_FILE._05483_ ),
    .X(\u_cpu.REG_FILE._05489_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11067_  (.A(\u_cpu.REG_FILE._05489_ ),
    .X(\u_cpu.REG_FILE._00847_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11068_  (.A0(\u_cpu.REG_FILE.rf[25][16] ),
    .A1(\u_cpu.REG_FILE._05252_ ),
    .S(\u_cpu.REG_FILE._05483_ ),
    .X(\u_cpu.REG_FILE._05490_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11069_  (.A(\u_cpu.REG_FILE._05490_ ),
    .X(\u_cpu.REG_FILE._00848_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11070_  (.A0(\u_cpu.REG_FILE.rf[25][17] ),
    .A1(\u_cpu.REG_FILE._05254_ ),
    .S(\u_cpu.REG_FILE._05483_ ),
    .X(\u_cpu.REG_FILE._05491_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11071_  (.A(\u_cpu.REG_FILE._05491_ ),
    .X(\u_cpu.REG_FILE._00849_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11072_  (.A0(\u_cpu.REG_FILE.rf[25][18] ),
    .A1(\u_cpu.REG_FILE._05256_ ),
    .S(\u_cpu.REG_FILE._05483_ ),
    .X(\u_cpu.REG_FILE._05492_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11073_  (.A(\u_cpu.REG_FILE._05492_ ),
    .X(\u_cpu.REG_FILE._00850_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11074_  (.A0(\u_cpu.REG_FILE.rf[25][19] ),
    .A1(\u_cpu.REG_FILE._05258_ ),
    .S(\u_cpu.REG_FILE._05483_ ),
    .X(\u_cpu.REG_FILE._05493_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11075_  (.A(\u_cpu.REG_FILE._05493_ ),
    .X(\u_cpu.REG_FILE._00851_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11076_  (.A(\u_cpu.REG_FILE._05471_ ),
    .X(\u_cpu.REG_FILE._05494_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11077_  (.A0(\u_cpu.REG_FILE.rf[25][20] ),
    .A1(\u_cpu.REG_FILE._05260_ ),
    .S(\u_cpu.REG_FILE._05494_ ),
    .X(\u_cpu.REG_FILE._05495_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11078_  (.A(\u_cpu.REG_FILE._05495_ ),
    .X(\u_cpu.REG_FILE._00852_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11079_  (.A0(\u_cpu.REG_FILE.rf[25][21] ),
    .A1(\u_cpu.REG_FILE._05263_ ),
    .S(\u_cpu.REG_FILE._05494_ ),
    .X(\u_cpu.REG_FILE._05496_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11080_  (.A(\u_cpu.REG_FILE._05496_ ),
    .X(\u_cpu.REG_FILE._00853_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11081_  (.A0(\u_cpu.REG_FILE.rf[25][22] ),
    .A1(\u_cpu.REG_FILE._05265_ ),
    .S(\u_cpu.REG_FILE._05494_ ),
    .X(\u_cpu.REG_FILE._05497_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11082_  (.A(\u_cpu.REG_FILE._05497_ ),
    .X(\u_cpu.REG_FILE._00854_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11083_  (.A0(\u_cpu.REG_FILE.rf[25][23] ),
    .A1(\u_cpu.REG_FILE._05267_ ),
    .S(\u_cpu.REG_FILE._05494_ ),
    .X(\u_cpu.REG_FILE._05498_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11084_  (.A(\u_cpu.REG_FILE._05498_ ),
    .X(\u_cpu.REG_FILE._00855_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11085_  (.A0(\u_cpu.REG_FILE.rf[25][24] ),
    .A1(\u_cpu.REG_FILE._05269_ ),
    .S(\u_cpu.REG_FILE._05494_ ),
    .X(\u_cpu.REG_FILE._05499_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11086_  (.A(\u_cpu.REG_FILE._05499_ ),
    .X(\u_cpu.REG_FILE._00856_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11087_  (.A0(\u_cpu.REG_FILE.rf[25][25] ),
    .A1(\u_cpu.REG_FILE._05271_ ),
    .S(\u_cpu.REG_FILE._05494_ ),
    .X(\u_cpu.REG_FILE._05500_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11088_  (.A(\u_cpu.REG_FILE._05500_ ),
    .X(\u_cpu.REG_FILE._00857_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11089_  (.A0(\u_cpu.REG_FILE.rf[25][26] ),
    .A1(\u_cpu.REG_FILE._05273_ ),
    .S(\u_cpu.REG_FILE._05494_ ),
    .X(\u_cpu.REG_FILE._05501_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11090_  (.A(\u_cpu.REG_FILE._05501_ ),
    .X(\u_cpu.REG_FILE._00858_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11091_  (.A0(\u_cpu.REG_FILE.rf[25][27] ),
    .A1(\u_cpu.REG_FILE._05275_ ),
    .S(\u_cpu.REG_FILE._05494_ ),
    .X(\u_cpu.REG_FILE._05502_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11092_  (.A(\u_cpu.REG_FILE._05502_ ),
    .X(\u_cpu.REG_FILE._00859_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11093_  (.A0(\u_cpu.REG_FILE.rf[25][28] ),
    .A1(\u_cpu.REG_FILE._05277_ ),
    .S(\u_cpu.REG_FILE._05494_ ),
    .X(\u_cpu.REG_FILE._05503_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11094_  (.A(\u_cpu.REG_FILE._05503_ ),
    .X(\u_cpu.REG_FILE._00860_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11095_  (.A0(\u_cpu.REG_FILE.rf[25][29] ),
    .A1(\u_cpu.REG_FILE._05279_ ),
    .S(\u_cpu.REG_FILE._05494_ ),
    .X(\u_cpu.REG_FILE._05504_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11096_  (.A(\u_cpu.REG_FILE._05504_ ),
    .X(\u_cpu.REG_FILE._00861_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11097_  (.A0(\u_cpu.REG_FILE.rf[25][30] ),
    .A1(\u_cpu.REG_FILE._05281_ ),
    .S(\u_cpu.REG_FILE._05471_ ),
    .X(\u_cpu.REG_FILE._05505_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11098_  (.A(\u_cpu.REG_FILE._05505_ ),
    .X(\u_cpu.REG_FILE._00862_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11099_  (.A0(\u_cpu.REG_FILE.rf[25][31] ),
    .A1(\u_cpu.REG_FILE._05283_ ),
    .S(\u_cpu.REG_FILE._05471_ ),
    .X(\u_cpu.REG_FILE._05506_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11100_  (.A(\u_cpu.REG_FILE._05506_ ),
    .X(\u_cpu.REG_FILE._00863_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.REG_FILE._11101_  (.A_N(\u_cpu.REG_FILE._04425_ ),
    .B(\u_cpu.REG_FILE._04747_ ),
    .C(\u_cpu.REG_FILE.a3[4] ),
    .D(\u_cpu.REG_FILE.a3[3] ),
    .X(\u_cpu.REG_FILE._05507_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11102_  (.A(\u_cpu.REG_FILE._05507_ ),
    .X(\u_cpu.REG_FILE._05508_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11103_  (.A(\u_cpu.REG_FILE._05508_ ),
    .X(\u_cpu.REG_FILE._05509_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11104_  (.A0(\u_cpu.REG_FILE.rf[26][0] ),
    .A1(\u_cpu.REG_FILE._05216_ ),
    .S(\u_cpu.REG_FILE._05509_ ),
    .X(\u_cpu.REG_FILE._05510_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11105_  (.A(\u_cpu.REG_FILE._05510_ ),
    .X(\u_cpu.REG_FILE._00864_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11106_  (.A0(\u_cpu.REG_FILE.rf[26][1] ),
    .A1(\u_cpu.REG_FILE._05221_ ),
    .S(\u_cpu.REG_FILE._05509_ ),
    .X(\u_cpu.REG_FILE._05511_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11107_  (.A(\u_cpu.REG_FILE._05511_ ),
    .X(\u_cpu.REG_FILE._00865_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11108_  (.A0(\u_cpu.REG_FILE.rf[26][2] ),
    .A1(\u_cpu.REG_FILE._05223_ ),
    .S(\u_cpu.REG_FILE._05509_ ),
    .X(\u_cpu.REG_FILE._05512_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11109_  (.A(\u_cpu.REG_FILE._05512_ ),
    .X(\u_cpu.REG_FILE._00866_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11110_  (.A0(\u_cpu.REG_FILE.rf[26][3] ),
    .A1(\u_cpu.REG_FILE._05225_ ),
    .S(\u_cpu.REG_FILE._05509_ ),
    .X(\u_cpu.REG_FILE._05513_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11111_  (.A(\u_cpu.REG_FILE._05513_ ),
    .X(\u_cpu.REG_FILE._00867_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11112_  (.A0(\u_cpu.REG_FILE.rf[26][4] ),
    .A1(\u_cpu.REG_FILE._05227_ ),
    .S(\u_cpu.REG_FILE._05509_ ),
    .X(\u_cpu.REG_FILE._05514_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11113_  (.A(\u_cpu.REG_FILE._05514_ ),
    .X(\u_cpu.REG_FILE._00868_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11114_  (.A0(\u_cpu.REG_FILE.rf[26][5] ),
    .A1(\u_cpu.REG_FILE._05229_ ),
    .S(\u_cpu.REG_FILE._05509_ ),
    .X(\u_cpu.REG_FILE._05515_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11115_  (.A(\u_cpu.REG_FILE._05515_ ),
    .X(\u_cpu.REG_FILE._00869_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11116_  (.A0(\u_cpu.REG_FILE.rf[26][6] ),
    .A1(\u_cpu.REG_FILE._05231_ ),
    .S(\u_cpu.REG_FILE._05509_ ),
    .X(\u_cpu.REG_FILE._05516_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11117_  (.A(\u_cpu.REG_FILE._05516_ ),
    .X(\u_cpu.REG_FILE._00870_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11118_  (.A0(\u_cpu.REG_FILE.rf[26][7] ),
    .A1(\u_cpu.REG_FILE._05233_ ),
    .S(\u_cpu.REG_FILE._05509_ ),
    .X(\u_cpu.REG_FILE._05517_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11119_  (.A(\u_cpu.REG_FILE._05517_ ),
    .X(\u_cpu.REG_FILE._00871_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11120_  (.A0(\u_cpu.REG_FILE.rf[26][8] ),
    .A1(\u_cpu.REG_FILE._05235_ ),
    .S(\u_cpu.REG_FILE._05509_ ),
    .X(\u_cpu.REG_FILE._05518_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11121_  (.A(\u_cpu.REG_FILE._05518_ ),
    .X(\u_cpu.REG_FILE._00872_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11122_  (.A0(\u_cpu.REG_FILE.rf[26][9] ),
    .A1(\u_cpu.REG_FILE._05237_ ),
    .S(\u_cpu.REG_FILE._05509_ ),
    .X(\u_cpu.REG_FILE._05519_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11123_  (.A(\u_cpu.REG_FILE._05519_ ),
    .X(\u_cpu.REG_FILE._00873_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11124_  (.A(\u_cpu.REG_FILE._05508_ ),
    .X(\u_cpu.REG_FILE._05520_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11125_  (.A0(\u_cpu.REG_FILE.rf[26][10] ),
    .A1(\u_cpu.REG_FILE._05239_ ),
    .S(\u_cpu.REG_FILE._05520_ ),
    .X(\u_cpu.REG_FILE._05521_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11126_  (.A(\u_cpu.REG_FILE._05521_ ),
    .X(\u_cpu.REG_FILE._00874_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11127_  (.A0(\u_cpu.REG_FILE.rf[26][11] ),
    .A1(\u_cpu.REG_FILE._05242_ ),
    .S(\u_cpu.REG_FILE._05520_ ),
    .X(\u_cpu.REG_FILE._05522_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11128_  (.A(\u_cpu.REG_FILE._05522_ ),
    .X(\u_cpu.REG_FILE._00875_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11129_  (.A0(\u_cpu.REG_FILE.rf[26][12] ),
    .A1(\u_cpu.REG_FILE._05244_ ),
    .S(\u_cpu.REG_FILE._05520_ ),
    .X(\u_cpu.REG_FILE._05523_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11130_  (.A(\u_cpu.REG_FILE._05523_ ),
    .X(\u_cpu.REG_FILE._00876_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11131_  (.A0(\u_cpu.REG_FILE.rf[26][13] ),
    .A1(\u_cpu.REG_FILE._05246_ ),
    .S(\u_cpu.REG_FILE._05520_ ),
    .X(\u_cpu.REG_FILE._05524_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11132_  (.A(\u_cpu.REG_FILE._05524_ ),
    .X(\u_cpu.REG_FILE._00877_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11133_  (.A0(\u_cpu.REG_FILE.rf[26][14] ),
    .A1(\u_cpu.REG_FILE._05248_ ),
    .S(\u_cpu.REG_FILE._05520_ ),
    .X(\u_cpu.REG_FILE._05525_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11134_  (.A(\u_cpu.REG_FILE._05525_ ),
    .X(\u_cpu.REG_FILE._00878_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11135_  (.A0(\u_cpu.REG_FILE.rf[26][15] ),
    .A1(\u_cpu.REG_FILE._05250_ ),
    .S(\u_cpu.REG_FILE._05520_ ),
    .X(\u_cpu.REG_FILE._05526_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11136_  (.A(\u_cpu.REG_FILE._05526_ ),
    .X(\u_cpu.REG_FILE._00879_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11137_  (.A0(\u_cpu.REG_FILE.rf[26][16] ),
    .A1(\u_cpu.REG_FILE._05252_ ),
    .S(\u_cpu.REG_FILE._05520_ ),
    .X(\u_cpu.REG_FILE._05527_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11138_  (.A(\u_cpu.REG_FILE._05527_ ),
    .X(\u_cpu.REG_FILE._00880_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11139_  (.A0(\u_cpu.REG_FILE.rf[26][17] ),
    .A1(\u_cpu.REG_FILE._05254_ ),
    .S(\u_cpu.REG_FILE._05520_ ),
    .X(\u_cpu.REG_FILE._05528_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11140_  (.A(\u_cpu.REG_FILE._05528_ ),
    .X(\u_cpu.REG_FILE._00881_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11141_  (.A0(\u_cpu.REG_FILE.rf[26][18] ),
    .A1(\u_cpu.REG_FILE._05256_ ),
    .S(\u_cpu.REG_FILE._05520_ ),
    .X(\u_cpu.REG_FILE._05529_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11142_  (.A(\u_cpu.REG_FILE._05529_ ),
    .X(\u_cpu.REG_FILE._00882_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11143_  (.A0(\u_cpu.REG_FILE.rf[26][19] ),
    .A1(\u_cpu.REG_FILE._05258_ ),
    .S(\u_cpu.REG_FILE._05520_ ),
    .X(\u_cpu.REG_FILE._05530_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11144_  (.A(\u_cpu.REG_FILE._05530_ ),
    .X(\u_cpu.REG_FILE._00883_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11145_  (.A(\u_cpu.REG_FILE._05508_ ),
    .X(\u_cpu.REG_FILE._05531_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11146_  (.A0(\u_cpu.REG_FILE.rf[26][20] ),
    .A1(\u_cpu.REG_FILE._05260_ ),
    .S(\u_cpu.REG_FILE._05531_ ),
    .X(\u_cpu.REG_FILE._05532_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11147_  (.A(\u_cpu.REG_FILE._05532_ ),
    .X(\u_cpu.REG_FILE._00884_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11148_  (.A0(\u_cpu.REG_FILE.rf[26][21] ),
    .A1(\u_cpu.REG_FILE._05263_ ),
    .S(\u_cpu.REG_FILE._05531_ ),
    .X(\u_cpu.REG_FILE._05533_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11149_  (.A(\u_cpu.REG_FILE._05533_ ),
    .X(\u_cpu.REG_FILE._00885_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11150_  (.A0(\u_cpu.REG_FILE.rf[26][22] ),
    .A1(\u_cpu.REG_FILE._05265_ ),
    .S(\u_cpu.REG_FILE._05531_ ),
    .X(\u_cpu.REG_FILE._05534_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11151_  (.A(\u_cpu.REG_FILE._05534_ ),
    .X(\u_cpu.REG_FILE._00886_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11152_  (.A0(\u_cpu.REG_FILE.rf[26][23] ),
    .A1(\u_cpu.REG_FILE._05267_ ),
    .S(\u_cpu.REG_FILE._05531_ ),
    .X(\u_cpu.REG_FILE._05535_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11153_  (.A(\u_cpu.REG_FILE._05535_ ),
    .X(\u_cpu.REG_FILE._00887_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11154_  (.A0(\u_cpu.REG_FILE.rf[26][24] ),
    .A1(\u_cpu.REG_FILE._05269_ ),
    .S(\u_cpu.REG_FILE._05531_ ),
    .X(\u_cpu.REG_FILE._05536_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11155_  (.A(\u_cpu.REG_FILE._05536_ ),
    .X(\u_cpu.REG_FILE._00888_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11156_  (.A0(\u_cpu.REG_FILE.rf[26][25] ),
    .A1(\u_cpu.REG_FILE._05271_ ),
    .S(\u_cpu.REG_FILE._05531_ ),
    .X(\u_cpu.REG_FILE._05537_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11157_  (.A(\u_cpu.REG_FILE._05537_ ),
    .X(\u_cpu.REG_FILE._00889_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11158_  (.A0(\u_cpu.REG_FILE.rf[26][26] ),
    .A1(\u_cpu.REG_FILE._05273_ ),
    .S(\u_cpu.REG_FILE._05531_ ),
    .X(\u_cpu.REG_FILE._05538_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11159_  (.A(\u_cpu.REG_FILE._05538_ ),
    .X(\u_cpu.REG_FILE._00890_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11160_  (.A0(\u_cpu.REG_FILE.rf[26][27] ),
    .A1(\u_cpu.REG_FILE._05275_ ),
    .S(\u_cpu.REG_FILE._05531_ ),
    .X(\u_cpu.REG_FILE._05539_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11161_  (.A(\u_cpu.REG_FILE._05539_ ),
    .X(\u_cpu.REG_FILE._00891_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11162_  (.A0(\u_cpu.REG_FILE.rf[26][28] ),
    .A1(\u_cpu.REG_FILE._05277_ ),
    .S(\u_cpu.REG_FILE._05531_ ),
    .X(\u_cpu.REG_FILE._05540_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11163_  (.A(\u_cpu.REG_FILE._05540_ ),
    .X(\u_cpu.REG_FILE._00892_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11164_  (.A0(\u_cpu.REG_FILE.rf[26][29] ),
    .A1(\u_cpu.REG_FILE._05279_ ),
    .S(\u_cpu.REG_FILE._05531_ ),
    .X(\u_cpu.REG_FILE._05541_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11165_  (.A(\u_cpu.REG_FILE._05541_ ),
    .X(\u_cpu.REG_FILE._00893_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11166_  (.A0(\u_cpu.REG_FILE.rf[26][30] ),
    .A1(\u_cpu.REG_FILE._05281_ ),
    .S(\u_cpu.REG_FILE._05508_ ),
    .X(\u_cpu.REG_FILE._05542_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11167_  (.A(\u_cpu.REG_FILE._05542_ ),
    .X(\u_cpu.REG_FILE._00894_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11168_  (.A0(\u_cpu.REG_FILE.rf[26][31] ),
    .A1(\u_cpu.REG_FILE._05283_ ),
    .S(\u_cpu.REG_FILE._05508_ ),
    .X(\u_cpu.REG_FILE._05543_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11169_  (.A(\u_cpu.REG_FILE._05543_ ),
    .X(\u_cpu.REG_FILE._00895_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.REG_FILE._11170_  (.A_N(\u_cpu.REG_FILE._04425_ ),
    .B(\u_cpu.REG_FILE._04495_ ),
    .C(\u_cpu.REG_FILE.a3[4] ),
    .D(\u_cpu.REG_FILE.a3[3] ),
    .X(\u_cpu.REG_FILE._05544_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11171_  (.A(\u_cpu.REG_FILE._05544_ ),
    .X(\u_cpu.REG_FILE._05545_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11172_  (.A(\u_cpu.REG_FILE._05545_ ),
    .X(\u_cpu.REG_FILE._05546_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11173_  (.A0(\u_cpu.REG_FILE.rf[27][0] ),
    .A1(\u_cpu.REG_FILE._05216_ ),
    .S(\u_cpu.REG_FILE._05546_ ),
    .X(\u_cpu.REG_FILE._05547_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11174_  (.A(\u_cpu.REG_FILE._05547_ ),
    .X(\u_cpu.REG_FILE._00896_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11175_  (.A0(\u_cpu.REG_FILE.rf[27][1] ),
    .A1(\u_cpu.REG_FILE._05221_ ),
    .S(\u_cpu.REG_FILE._05546_ ),
    .X(\u_cpu.REG_FILE._05548_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11176_  (.A(\u_cpu.REG_FILE._05548_ ),
    .X(\u_cpu.REG_FILE._00897_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11177_  (.A0(\u_cpu.REG_FILE.rf[27][2] ),
    .A1(\u_cpu.REG_FILE._05223_ ),
    .S(\u_cpu.REG_FILE._05546_ ),
    .X(\u_cpu.REG_FILE._05549_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11178_  (.A(\u_cpu.REG_FILE._05549_ ),
    .X(\u_cpu.REG_FILE._00898_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11179_  (.A0(\u_cpu.REG_FILE.rf[27][3] ),
    .A1(\u_cpu.REG_FILE._05225_ ),
    .S(\u_cpu.REG_FILE._05546_ ),
    .X(\u_cpu.REG_FILE._05550_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11180_  (.A(\u_cpu.REG_FILE._05550_ ),
    .X(\u_cpu.REG_FILE._00899_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11181_  (.A0(\u_cpu.REG_FILE.rf[27][4] ),
    .A1(\u_cpu.REG_FILE._05227_ ),
    .S(\u_cpu.REG_FILE._05546_ ),
    .X(\u_cpu.REG_FILE._05551_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11182_  (.A(\u_cpu.REG_FILE._05551_ ),
    .X(\u_cpu.REG_FILE._00900_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11183_  (.A0(\u_cpu.REG_FILE.rf[27][5] ),
    .A1(\u_cpu.REG_FILE._05229_ ),
    .S(\u_cpu.REG_FILE._05546_ ),
    .X(\u_cpu.REG_FILE._05552_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11184_  (.A(\u_cpu.REG_FILE._05552_ ),
    .X(\u_cpu.REG_FILE._00901_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11185_  (.A0(\u_cpu.REG_FILE.rf[27][6] ),
    .A1(\u_cpu.REG_FILE._05231_ ),
    .S(\u_cpu.REG_FILE._05546_ ),
    .X(\u_cpu.REG_FILE._05553_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11186_  (.A(\u_cpu.REG_FILE._05553_ ),
    .X(\u_cpu.REG_FILE._00902_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11187_  (.A0(\u_cpu.REG_FILE.rf[27][7] ),
    .A1(\u_cpu.REG_FILE._05233_ ),
    .S(\u_cpu.REG_FILE._05546_ ),
    .X(\u_cpu.REG_FILE._05554_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11188_  (.A(\u_cpu.REG_FILE._05554_ ),
    .X(\u_cpu.REG_FILE._00903_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11189_  (.A0(\u_cpu.REG_FILE.rf[27][8] ),
    .A1(\u_cpu.REG_FILE._05235_ ),
    .S(\u_cpu.REG_FILE._05546_ ),
    .X(\u_cpu.REG_FILE._05555_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11190_  (.A(\u_cpu.REG_FILE._05555_ ),
    .X(\u_cpu.REG_FILE._00904_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11191_  (.A0(\u_cpu.REG_FILE.rf[27][9] ),
    .A1(\u_cpu.REG_FILE._05237_ ),
    .S(\u_cpu.REG_FILE._05546_ ),
    .X(\u_cpu.REG_FILE._05556_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11192_  (.A(\u_cpu.REG_FILE._05556_ ),
    .X(\u_cpu.REG_FILE._00905_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11193_  (.A(\u_cpu.REG_FILE._05545_ ),
    .X(\u_cpu.REG_FILE._05557_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11194_  (.A0(\u_cpu.REG_FILE.rf[27][10] ),
    .A1(\u_cpu.REG_FILE._05239_ ),
    .S(\u_cpu.REG_FILE._05557_ ),
    .X(\u_cpu.REG_FILE._05558_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11195_  (.A(\u_cpu.REG_FILE._05558_ ),
    .X(\u_cpu.REG_FILE._00906_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11196_  (.A0(\u_cpu.REG_FILE.rf[27][11] ),
    .A1(\u_cpu.REG_FILE._05242_ ),
    .S(\u_cpu.REG_FILE._05557_ ),
    .X(\u_cpu.REG_FILE._05559_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11197_  (.A(\u_cpu.REG_FILE._05559_ ),
    .X(\u_cpu.REG_FILE._00907_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11198_  (.A0(\u_cpu.REG_FILE.rf[27][12] ),
    .A1(\u_cpu.REG_FILE._05244_ ),
    .S(\u_cpu.REG_FILE._05557_ ),
    .X(\u_cpu.REG_FILE._05560_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11199_  (.A(\u_cpu.REG_FILE._05560_ ),
    .X(\u_cpu.REG_FILE._00908_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11200_  (.A0(\u_cpu.REG_FILE.rf[27][13] ),
    .A1(\u_cpu.REG_FILE._05246_ ),
    .S(\u_cpu.REG_FILE._05557_ ),
    .X(\u_cpu.REG_FILE._05561_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11201_  (.A(\u_cpu.REG_FILE._05561_ ),
    .X(\u_cpu.REG_FILE._00909_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11202_  (.A0(\u_cpu.REG_FILE.rf[27][14] ),
    .A1(\u_cpu.REG_FILE._05248_ ),
    .S(\u_cpu.REG_FILE._05557_ ),
    .X(\u_cpu.REG_FILE._05562_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11203_  (.A(\u_cpu.REG_FILE._05562_ ),
    .X(\u_cpu.REG_FILE._00910_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11204_  (.A0(\u_cpu.REG_FILE.rf[27][15] ),
    .A1(\u_cpu.REG_FILE._05250_ ),
    .S(\u_cpu.REG_FILE._05557_ ),
    .X(\u_cpu.REG_FILE._05563_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11205_  (.A(\u_cpu.REG_FILE._05563_ ),
    .X(\u_cpu.REG_FILE._00911_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11206_  (.A0(\u_cpu.REG_FILE.rf[27][16] ),
    .A1(\u_cpu.REG_FILE._05252_ ),
    .S(\u_cpu.REG_FILE._05557_ ),
    .X(\u_cpu.REG_FILE._05564_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11207_  (.A(\u_cpu.REG_FILE._05564_ ),
    .X(\u_cpu.REG_FILE._00912_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11208_  (.A0(\u_cpu.REG_FILE.rf[27][17] ),
    .A1(\u_cpu.REG_FILE._05254_ ),
    .S(\u_cpu.REG_FILE._05557_ ),
    .X(\u_cpu.REG_FILE._05565_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11209_  (.A(\u_cpu.REG_FILE._05565_ ),
    .X(\u_cpu.REG_FILE._00913_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11210_  (.A0(\u_cpu.REG_FILE.rf[27][18] ),
    .A1(\u_cpu.REG_FILE._05256_ ),
    .S(\u_cpu.REG_FILE._05557_ ),
    .X(\u_cpu.REG_FILE._05566_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11211_  (.A(\u_cpu.REG_FILE._05566_ ),
    .X(\u_cpu.REG_FILE._00914_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11212_  (.A0(\u_cpu.REG_FILE.rf[27][19] ),
    .A1(\u_cpu.REG_FILE._05258_ ),
    .S(\u_cpu.REG_FILE._05557_ ),
    .X(\u_cpu.REG_FILE._05567_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11213_  (.A(\u_cpu.REG_FILE._05567_ ),
    .X(\u_cpu.REG_FILE._00915_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11214_  (.A(\u_cpu.REG_FILE._05545_ ),
    .X(\u_cpu.REG_FILE._05568_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11215_  (.A0(\u_cpu.REG_FILE.rf[27][20] ),
    .A1(\u_cpu.REG_FILE._05260_ ),
    .S(\u_cpu.REG_FILE._05568_ ),
    .X(\u_cpu.REG_FILE._05569_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11216_  (.A(\u_cpu.REG_FILE._05569_ ),
    .X(\u_cpu.REG_FILE._00916_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11217_  (.A0(\u_cpu.REG_FILE.rf[27][21] ),
    .A1(\u_cpu.REG_FILE._05263_ ),
    .S(\u_cpu.REG_FILE._05568_ ),
    .X(\u_cpu.REG_FILE._05570_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11218_  (.A(\u_cpu.REG_FILE._05570_ ),
    .X(\u_cpu.REG_FILE._00917_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11219_  (.A0(\u_cpu.REG_FILE.rf[27][22] ),
    .A1(\u_cpu.REG_FILE._05265_ ),
    .S(\u_cpu.REG_FILE._05568_ ),
    .X(\u_cpu.REG_FILE._05571_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11220_  (.A(\u_cpu.REG_FILE._05571_ ),
    .X(\u_cpu.REG_FILE._00918_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11221_  (.A0(\u_cpu.REG_FILE.rf[27][23] ),
    .A1(\u_cpu.REG_FILE._05267_ ),
    .S(\u_cpu.REG_FILE._05568_ ),
    .X(\u_cpu.REG_FILE._05572_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11222_  (.A(\u_cpu.REG_FILE._05572_ ),
    .X(\u_cpu.REG_FILE._00919_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11223_  (.A0(\u_cpu.REG_FILE.rf[27][24] ),
    .A1(\u_cpu.REG_FILE._05269_ ),
    .S(\u_cpu.REG_FILE._05568_ ),
    .X(\u_cpu.REG_FILE._05573_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11224_  (.A(\u_cpu.REG_FILE._05573_ ),
    .X(\u_cpu.REG_FILE._00920_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11225_  (.A0(\u_cpu.REG_FILE.rf[27][25] ),
    .A1(\u_cpu.REG_FILE._05271_ ),
    .S(\u_cpu.REG_FILE._05568_ ),
    .X(\u_cpu.REG_FILE._05574_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11226_  (.A(\u_cpu.REG_FILE._05574_ ),
    .X(\u_cpu.REG_FILE._00921_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11227_  (.A0(\u_cpu.REG_FILE.rf[27][26] ),
    .A1(\u_cpu.REG_FILE._05273_ ),
    .S(\u_cpu.REG_FILE._05568_ ),
    .X(\u_cpu.REG_FILE._05575_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11228_  (.A(\u_cpu.REG_FILE._05575_ ),
    .X(\u_cpu.REG_FILE._00922_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11229_  (.A0(\u_cpu.REG_FILE.rf[27][27] ),
    .A1(\u_cpu.REG_FILE._05275_ ),
    .S(\u_cpu.REG_FILE._05568_ ),
    .X(\u_cpu.REG_FILE._05576_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11230_  (.A(\u_cpu.REG_FILE._05576_ ),
    .X(\u_cpu.REG_FILE._00923_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11231_  (.A0(\u_cpu.REG_FILE.rf[27][28] ),
    .A1(\u_cpu.REG_FILE._05277_ ),
    .S(\u_cpu.REG_FILE._05568_ ),
    .X(\u_cpu.REG_FILE._05577_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11232_  (.A(\u_cpu.REG_FILE._05577_ ),
    .X(\u_cpu.REG_FILE._00924_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11233_  (.A0(\u_cpu.REG_FILE.rf[27][29] ),
    .A1(\u_cpu.REG_FILE._05279_ ),
    .S(\u_cpu.REG_FILE._05568_ ),
    .X(\u_cpu.REG_FILE._05578_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11234_  (.A(\u_cpu.REG_FILE._05578_ ),
    .X(\u_cpu.REG_FILE._00925_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11235_  (.A0(\u_cpu.REG_FILE.rf[27][30] ),
    .A1(\u_cpu.REG_FILE._05281_ ),
    .S(\u_cpu.REG_FILE._05545_ ),
    .X(\u_cpu.REG_FILE._05579_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11236_  (.A(\u_cpu.REG_FILE._05579_ ),
    .X(\u_cpu.REG_FILE._00926_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11237_  (.A0(\u_cpu.REG_FILE.rf[27][31] ),
    .A1(\u_cpu.REG_FILE._05283_ ),
    .S(\u_cpu.REG_FILE._05545_ ),
    .X(\u_cpu.REG_FILE._05580_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11238_  (.A(\u_cpu.REG_FILE._05580_ ),
    .X(\u_cpu.REG_FILE._00927_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu.REG_FILE._11239_  (.A(\u_cpu.REG_FILE._04496_ ),
    .B(\u_cpu.REG_FILE._04422_ ),
    .C(\u_cpu.REG_FILE._04494_ ),
    .D(\u_cpu.REG_FILE._04643_ ),
    .Y(\u_cpu.REG_FILE._05581_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11240_  (.A(\u_cpu.REG_FILE._05581_ ),
    .X(\u_cpu.REG_FILE._05582_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11241_  (.A0(\u_cpu.REG_FILE._04420_ ),
    .A1(\u_cpu.REG_FILE.rf[28][0] ),
    .S(\u_cpu.REG_FILE._05582_ ),
    .X(\u_cpu.REG_FILE._05583_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11242_  (.A(\u_cpu.REG_FILE._05583_ ),
    .X(\u_cpu.REG_FILE._00928_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11243_  (.A0(\u_cpu.REG_FILE._04430_ ),
    .A1(\u_cpu.REG_FILE.rf[28][1] ),
    .S(\u_cpu.REG_FILE._05582_ ),
    .X(\u_cpu.REG_FILE._05584_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11244_  (.A(\u_cpu.REG_FILE._05584_ ),
    .X(\u_cpu.REG_FILE._00929_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11245_  (.A0(\u_cpu.REG_FILE._04432_ ),
    .A1(\u_cpu.REG_FILE.rf[28][2] ),
    .S(\u_cpu.REG_FILE._05582_ ),
    .X(\u_cpu.REG_FILE._05585_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11246_  (.A(\u_cpu.REG_FILE._05585_ ),
    .X(\u_cpu.REG_FILE._00930_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11247_  (.A0(\u_cpu.REG_FILE._04434_ ),
    .A1(\u_cpu.REG_FILE.rf[28][3] ),
    .S(\u_cpu.REG_FILE._05582_ ),
    .X(\u_cpu.REG_FILE._05586_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11248_  (.A(\u_cpu.REG_FILE._05586_ ),
    .X(\u_cpu.REG_FILE._00931_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11249_  (.A0(\u_cpu.REG_FILE._04436_ ),
    .A1(\u_cpu.REG_FILE.rf[28][4] ),
    .S(\u_cpu.REG_FILE._05582_ ),
    .X(\u_cpu.REG_FILE._05587_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11250_  (.A(\u_cpu.REG_FILE._05587_ ),
    .X(\u_cpu.REG_FILE._00932_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11251_  (.A0(\u_cpu.REG_FILE._04438_ ),
    .A1(\u_cpu.REG_FILE.rf[28][5] ),
    .S(\u_cpu.REG_FILE._05582_ ),
    .X(\u_cpu.REG_FILE._05588_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11252_  (.A(\u_cpu.REG_FILE._05588_ ),
    .X(\u_cpu.REG_FILE._00933_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11253_  (.A0(\u_cpu.REG_FILE._04440_ ),
    .A1(\u_cpu.REG_FILE.rf[28][6] ),
    .S(\u_cpu.REG_FILE._05582_ ),
    .X(\u_cpu.REG_FILE._05589_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11254_  (.A(\u_cpu.REG_FILE._05589_ ),
    .X(\u_cpu.REG_FILE._00934_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11255_  (.A0(\u_cpu.REG_FILE._04442_ ),
    .A1(\u_cpu.REG_FILE.rf[28][7] ),
    .S(\u_cpu.REG_FILE._05582_ ),
    .X(\u_cpu.REG_FILE._05590_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11256_  (.A(\u_cpu.REG_FILE._05590_ ),
    .X(\u_cpu.REG_FILE._00935_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11257_  (.A0(\u_cpu.REG_FILE._04444_ ),
    .A1(\u_cpu.REG_FILE.rf[28][8] ),
    .S(\u_cpu.REG_FILE._05582_ ),
    .X(\u_cpu.REG_FILE._05591_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11258_  (.A(\u_cpu.REG_FILE._05591_ ),
    .X(\u_cpu.REG_FILE._00936_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11259_  (.A0(\u_cpu.REG_FILE._04446_ ),
    .A1(\u_cpu.REG_FILE.rf[28][9] ),
    .S(\u_cpu.REG_FILE._05582_ ),
    .X(\u_cpu.REG_FILE._05592_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11260_  (.A(\u_cpu.REG_FILE._05592_ ),
    .X(\u_cpu.REG_FILE._00937_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11261_  (.A(\u_cpu.REG_FILE._05581_ ),
    .X(\u_cpu.REG_FILE._05593_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11262_  (.A0(\u_cpu.REG_FILE._04448_ ),
    .A1(\u_cpu.REG_FILE.rf[28][10] ),
    .S(\u_cpu.REG_FILE._05593_ ),
    .X(\u_cpu.REG_FILE._05594_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11263_  (.A(\u_cpu.REG_FILE._05594_ ),
    .X(\u_cpu.REG_FILE._00938_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11264_  (.A0(\u_cpu.REG_FILE._04451_ ),
    .A1(\u_cpu.REG_FILE.rf[28][11] ),
    .S(\u_cpu.REG_FILE._05593_ ),
    .X(\u_cpu.REG_FILE._05595_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11265_  (.A(\u_cpu.REG_FILE._05595_ ),
    .X(\u_cpu.REG_FILE._00939_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11266_  (.A0(\u_cpu.REG_FILE._04453_ ),
    .A1(\u_cpu.REG_FILE.rf[28][12] ),
    .S(\u_cpu.REG_FILE._05593_ ),
    .X(\u_cpu.REG_FILE._05596_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11267_  (.A(\u_cpu.REG_FILE._05596_ ),
    .X(\u_cpu.REG_FILE._00940_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11268_  (.A0(\u_cpu.REG_FILE._04455_ ),
    .A1(\u_cpu.REG_FILE.rf[28][13] ),
    .S(\u_cpu.REG_FILE._05593_ ),
    .X(\u_cpu.REG_FILE._05597_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11269_  (.A(\u_cpu.REG_FILE._05597_ ),
    .X(\u_cpu.REG_FILE._00941_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11270_  (.A0(\u_cpu.REG_FILE._04457_ ),
    .A1(\u_cpu.REG_FILE.rf[28][14] ),
    .S(\u_cpu.REG_FILE._05593_ ),
    .X(\u_cpu.REG_FILE._05598_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11271_  (.A(\u_cpu.REG_FILE._05598_ ),
    .X(\u_cpu.REG_FILE._00942_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11272_  (.A0(\u_cpu.REG_FILE._04459_ ),
    .A1(\u_cpu.REG_FILE.rf[28][15] ),
    .S(\u_cpu.REG_FILE._05593_ ),
    .X(\u_cpu.REG_FILE._05599_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11273_  (.A(\u_cpu.REG_FILE._05599_ ),
    .X(\u_cpu.REG_FILE._00943_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11274_  (.A0(\u_cpu.REG_FILE._04461_ ),
    .A1(\u_cpu.REG_FILE.rf[28][16] ),
    .S(\u_cpu.REG_FILE._05593_ ),
    .X(\u_cpu.REG_FILE._05600_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11275_  (.A(\u_cpu.REG_FILE._05600_ ),
    .X(\u_cpu.REG_FILE._00944_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11276_  (.A0(\u_cpu.REG_FILE._04463_ ),
    .A1(\u_cpu.REG_FILE.rf[28][17] ),
    .S(\u_cpu.REG_FILE._05593_ ),
    .X(\u_cpu.REG_FILE._05601_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11277_  (.A(\u_cpu.REG_FILE._05601_ ),
    .X(\u_cpu.REG_FILE._00945_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11278_  (.A0(\u_cpu.REG_FILE._04465_ ),
    .A1(\u_cpu.REG_FILE.rf[28][18] ),
    .S(\u_cpu.REG_FILE._05593_ ),
    .X(\u_cpu.REG_FILE._05602_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11279_  (.A(\u_cpu.REG_FILE._05602_ ),
    .X(\u_cpu.REG_FILE._00946_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11280_  (.A0(\u_cpu.REG_FILE._04467_ ),
    .A1(\u_cpu.REG_FILE.rf[28][19] ),
    .S(\u_cpu.REG_FILE._05593_ ),
    .X(\u_cpu.REG_FILE._05603_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11281_  (.A(\u_cpu.REG_FILE._05603_ ),
    .X(\u_cpu.REG_FILE._00947_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11282_  (.A(\u_cpu.REG_FILE._05581_ ),
    .X(\u_cpu.REG_FILE._05604_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11283_  (.A0(\u_cpu.REG_FILE._04469_ ),
    .A1(\u_cpu.REG_FILE.rf[28][20] ),
    .S(\u_cpu.REG_FILE._05604_ ),
    .X(\u_cpu.REG_FILE._05605_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11284_  (.A(\u_cpu.REG_FILE._05605_ ),
    .X(\u_cpu.REG_FILE._00948_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11285_  (.A0(\u_cpu.REG_FILE._04472_ ),
    .A1(\u_cpu.REG_FILE.rf[28][21] ),
    .S(\u_cpu.REG_FILE._05604_ ),
    .X(\u_cpu.REG_FILE._05606_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11286_  (.A(\u_cpu.REG_FILE._05606_ ),
    .X(\u_cpu.REG_FILE._00949_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11287_  (.A0(\u_cpu.REG_FILE._04474_ ),
    .A1(\u_cpu.REG_FILE.rf[28][22] ),
    .S(\u_cpu.REG_FILE._05604_ ),
    .X(\u_cpu.REG_FILE._05607_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11288_  (.A(\u_cpu.REG_FILE._05607_ ),
    .X(\u_cpu.REG_FILE._00950_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11289_  (.A0(\u_cpu.REG_FILE._04476_ ),
    .A1(\u_cpu.REG_FILE.rf[28][23] ),
    .S(\u_cpu.REG_FILE._05604_ ),
    .X(\u_cpu.REG_FILE._05608_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11290_  (.A(\u_cpu.REG_FILE._05608_ ),
    .X(\u_cpu.REG_FILE._00951_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11291_  (.A0(\u_cpu.REG_FILE._04478_ ),
    .A1(\u_cpu.REG_FILE.rf[28][24] ),
    .S(\u_cpu.REG_FILE._05604_ ),
    .X(\u_cpu.REG_FILE._05609_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11292_  (.A(\u_cpu.REG_FILE._05609_ ),
    .X(\u_cpu.REG_FILE._00952_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11293_  (.A0(\u_cpu.REG_FILE._04480_ ),
    .A1(\u_cpu.REG_FILE.rf[28][25] ),
    .S(\u_cpu.REG_FILE._05604_ ),
    .X(\u_cpu.REG_FILE._05610_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11294_  (.A(\u_cpu.REG_FILE._05610_ ),
    .X(\u_cpu.REG_FILE._00953_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11295_  (.A0(\u_cpu.REG_FILE._04482_ ),
    .A1(\u_cpu.REG_FILE.rf[28][26] ),
    .S(\u_cpu.REG_FILE._05604_ ),
    .X(\u_cpu.REG_FILE._05611_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11296_  (.A(\u_cpu.REG_FILE._05611_ ),
    .X(\u_cpu.REG_FILE._00954_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11297_  (.A0(\u_cpu.REG_FILE._04484_ ),
    .A1(\u_cpu.REG_FILE.rf[28][27] ),
    .S(\u_cpu.REG_FILE._05604_ ),
    .X(\u_cpu.REG_FILE._05612_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11298_  (.A(\u_cpu.REG_FILE._05612_ ),
    .X(\u_cpu.REG_FILE._00955_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11299_  (.A0(\u_cpu.REG_FILE._04486_ ),
    .A1(\u_cpu.REG_FILE.rf[28][28] ),
    .S(\u_cpu.REG_FILE._05604_ ),
    .X(\u_cpu.REG_FILE._05613_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11300_  (.A(\u_cpu.REG_FILE._05613_ ),
    .X(\u_cpu.REG_FILE._00956_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11301_  (.A0(\u_cpu.REG_FILE._04488_ ),
    .A1(\u_cpu.REG_FILE.rf[28][29] ),
    .S(\u_cpu.REG_FILE._05604_ ),
    .X(\u_cpu.REG_FILE._05614_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11302_  (.A(\u_cpu.REG_FILE._05614_ ),
    .X(\u_cpu.REG_FILE._00957_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11303_  (.A0(\u_cpu.REG_FILE._04490_ ),
    .A1(\u_cpu.REG_FILE.rf[28][30] ),
    .S(\u_cpu.REG_FILE._05581_ ),
    .X(\u_cpu.REG_FILE._05615_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11304_  (.A(\u_cpu.REG_FILE._05615_ ),
    .X(\u_cpu.REG_FILE._00958_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11305_  (.A0(\u_cpu.REG_FILE._04492_ ),
    .A1(\u_cpu.REG_FILE.rf[28][31] ),
    .S(\u_cpu.REG_FILE._05581_ ),
    .X(\u_cpu.REG_FILE._05616_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11306_  (.A(\u_cpu.REG_FILE._05616_ ),
    .X(\u_cpu.REG_FILE._00959_ ));
 sky130_fd_sc_hd__and4b_2 \u_cpu.REG_FILE._11307_  (.A_N(\u_cpu.REG_FILE.a3[0] ),
    .B(\u_cpu.REG_FILE.we3 ),
    .C(\u_cpu.REG_FILE._04605_ ),
    .D(\u_cpu.REG_FILE.a3[1] ),
    .X(\u_cpu.REG_FILE._05617_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11308_  (.A(\u_cpu.REG_FILE._05617_ ),
    .X(\u_cpu.REG_FILE._05618_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11309_  (.A(\u_cpu.REG_FILE._05618_ ),
    .X(\u_cpu.REG_FILE._05619_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11310_  (.A0(\u_cpu.REG_FILE.rf[2][0] ),
    .A1(\u_cpu.REG_FILE._05216_ ),
    .S(\u_cpu.REG_FILE._05619_ ),
    .X(\u_cpu.REG_FILE._05620_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11311_  (.A(\u_cpu.REG_FILE._05620_ ),
    .X(\u_cpu.REG_FILE._00960_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11312_  (.A0(\u_cpu.REG_FILE.rf[2][1] ),
    .A1(\u_cpu.REG_FILE._05221_ ),
    .S(\u_cpu.REG_FILE._05619_ ),
    .X(\u_cpu.REG_FILE._05621_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11313_  (.A(\u_cpu.REG_FILE._05621_ ),
    .X(\u_cpu.REG_FILE._00961_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11314_  (.A0(\u_cpu.REG_FILE.rf[2][2] ),
    .A1(\u_cpu.REG_FILE._05223_ ),
    .S(\u_cpu.REG_FILE._05619_ ),
    .X(\u_cpu.REG_FILE._05622_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11315_  (.A(\u_cpu.REG_FILE._05622_ ),
    .X(\u_cpu.REG_FILE._00962_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11316_  (.A0(\u_cpu.REG_FILE.rf[2][3] ),
    .A1(\u_cpu.REG_FILE._05225_ ),
    .S(\u_cpu.REG_FILE._05619_ ),
    .X(\u_cpu.REG_FILE._05623_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11317_  (.A(\u_cpu.REG_FILE._05623_ ),
    .X(\u_cpu.REG_FILE._00963_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11318_  (.A0(\u_cpu.REG_FILE.rf[2][4] ),
    .A1(\u_cpu.REG_FILE._05227_ ),
    .S(\u_cpu.REG_FILE._05619_ ),
    .X(\u_cpu.REG_FILE._05624_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11319_  (.A(\u_cpu.REG_FILE._05624_ ),
    .X(\u_cpu.REG_FILE._00964_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11320_  (.A0(\u_cpu.REG_FILE.rf[2][5] ),
    .A1(\u_cpu.REG_FILE._05229_ ),
    .S(\u_cpu.REG_FILE._05619_ ),
    .X(\u_cpu.REG_FILE._05625_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11321_  (.A(\u_cpu.REG_FILE._05625_ ),
    .X(\u_cpu.REG_FILE._00965_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11322_  (.A0(\u_cpu.REG_FILE.rf[2][6] ),
    .A1(\u_cpu.REG_FILE._05231_ ),
    .S(\u_cpu.REG_FILE._05619_ ),
    .X(\u_cpu.REG_FILE._05626_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11323_  (.A(\u_cpu.REG_FILE._05626_ ),
    .X(\u_cpu.REG_FILE._00966_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11324_  (.A0(\u_cpu.REG_FILE.rf[2][7] ),
    .A1(\u_cpu.REG_FILE._05233_ ),
    .S(\u_cpu.REG_FILE._05619_ ),
    .X(\u_cpu.REG_FILE._05627_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11325_  (.A(\u_cpu.REG_FILE._05627_ ),
    .X(\u_cpu.REG_FILE._00967_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11326_  (.A0(\u_cpu.REG_FILE.rf[2][8] ),
    .A1(\u_cpu.REG_FILE._05235_ ),
    .S(\u_cpu.REG_FILE._05619_ ),
    .X(\u_cpu.REG_FILE._05628_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11327_  (.A(\u_cpu.REG_FILE._05628_ ),
    .X(\u_cpu.REG_FILE._00968_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11328_  (.A0(\u_cpu.REG_FILE.rf[2][9] ),
    .A1(\u_cpu.REG_FILE._05237_ ),
    .S(\u_cpu.REG_FILE._05619_ ),
    .X(\u_cpu.REG_FILE._05629_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11329_  (.A(\u_cpu.REG_FILE._05629_ ),
    .X(\u_cpu.REG_FILE._00969_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11330_  (.A(\u_cpu.REG_FILE._05618_ ),
    .X(\u_cpu.REG_FILE._05630_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11331_  (.A0(\u_cpu.REG_FILE.rf[2][10] ),
    .A1(\u_cpu.REG_FILE._05239_ ),
    .S(\u_cpu.REG_FILE._05630_ ),
    .X(\u_cpu.REG_FILE._05631_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11332_  (.A(\u_cpu.REG_FILE._05631_ ),
    .X(\u_cpu.REG_FILE._00970_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11333_  (.A0(\u_cpu.REG_FILE.rf[2][11] ),
    .A1(\u_cpu.REG_FILE._05242_ ),
    .S(\u_cpu.REG_FILE._05630_ ),
    .X(\u_cpu.REG_FILE._05632_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11334_  (.A(\u_cpu.REG_FILE._05632_ ),
    .X(\u_cpu.REG_FILE._00971_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11335_  (.A0(\u_cpu.REG_FILE.rf[2][12] ),
    .A1(\u_cpu.REG_FILE._05244_ ),
    .S(\u_cpu.REG_FILE._05630_ ),
    .X(\u_cpu.REG_FILE._05633_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11336_  (.A(\u_cpu.REG_FILE._05633_ ),
    .X(\u_cpu.REG_FILE._00972_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11337_  (.A0(\u_cpu.REG_FILE.rf[2][13] ),
    .A1(\u_cpu.REG_FILE._05246_ ),
    .S(\u_cpu.REG_FILE._05630_ ),
    .X(\u_cpu.REG_FILE._05634_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11338_  (.A(\u_cpu.REG_FILE._05634_ ),
    .X(\u_cpu.REG_FILE._00973_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11339_  (.A0(\u_cpu.REG_FILE.rf[2][14] ),
    .A1(\u_cpu.REG_FILE._05248_ ),
    .S(\u_cpu.REG_FILE._05630_ ),
    .X(\u_cpu.REG_FILE._05635_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11340_  (.A(\u_cpu.REG_FILE._05635_ ),
    .X(\u_cpu.REG_FILE._00974_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11341_  (.A0(\u_cpu.REG_FILE.rf[2][15] ),
    .A1(\u_cpu.REG_FILE._05250_ ),
    .S(\u_cpu.REG_FILE._05630_ ),
    .X(\u_cpu.REG_FILE._05636_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11342_  (.A(\u_cpu.REG_FILE._05636_ ),
    .X(\u_cpu.REG_FILE._00975_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11343_  (.A0(\u_cpu.REG_FILE.rf[2][16] ),
    .A1(\u_cpu.REG_FILE._05252_ ),
    .S(\u_cpu.REG_FILE._05630_ ),
    .X(\u_cpu.REG_FILE._05637_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11344_  (.A(\u_cpu.REG_FILE._05637_ ),
    .X(\u_cpu.REG_FILE._00976_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11345_  (.A0(\u_cpu.REG_FILE.rf[2][17] ),
    .A1(\u_cpu.REG_FILE._05254_ ),
    .S(\u_cpu.REG_FILE._05630_ ),
    .X(\u_cpu.REG_FILE._05638_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11346_  (.A(\u_cpu.REG_FILE._05638_ ),
    .X(\u_cpu.REG_FILE._00977_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11347_  (.A0(\u_cpu.REG_FILE.rf[2][18] ),
    .A1(\u_cpu.REG_FILE._05256_ ),
    .S(\u_cpu.REG_FILE._05630_ ),
    .X(\u_cpu.REG_FILE._05639_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11348_  (.A(\u_cpu.REG_FILE._05639_ ),
    .X(\u_cpu.REG_FILE._00978_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11349_  (.A0(\u_cpu.REG_FILE.rf[2][19] ),
    .A1(\u_cpu.REG_FILE._05258_ ),
    .S(\u_cpu.REG_FILE._05630_ ),
    .X(\u_cpu.REG_FILE._05640_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11350_  (.A(\u_cpu.REG_FILE._05640_ ),
    .X(\u_cpu.REG_FILE._00979_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11351_  (.A(\u_cpu.REG_FILE._05618_ ),
    .X(\u_cpu.REG_FILE._05641_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11352_  (.A0(\u_cpu.REG_FILE.rf[2][20] ),
    .A1(\u_cpu.REG_FILE._05260_ ),
    .S(\u_cpu.REG_FILE._05641_ ),
    .X(\u_cpu.REG_FILE._05642_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11353_  (.A(\u_cpu.REG_FILE._05642_ ),
    .X(\u_cpu.REG_FILE._00980_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11354_  (.A0(\u_cpu.REG_FILE.rf[2][21] ),
    .A1(\u_cpu.REG_FILE._05263_ ),
    .S(\u_cpu.REG_FILE._05641_ ),
    .X(\u_cpu.REG_FILE._05643_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11355_  (.A(\u_cpu.REG_FILE._05643_ ),
    .X(\u_cpu.REG_FILE._00981_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11356_  (.A0(\u_cpu.REG_FILE.rf[2][22] ),
    .A1(\u_cpu.REG_FILE._05265_ ),
    .S(\u_cpu.REG_FILE._05641_ ),
    .X(\u_cpu.REG_FILE._05644_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11357_  (.A(\u_cpu.REG_FILE._05644_ ),
    .X(\u_cpu.REG_FILE._00982_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11358_  (.A0(\u_cpu.REG_FILE.rf[2][23] ),
    .A1(\u_cpu.REG_FILE._05267_ ),
    .S(\u_cpu.REG_FILE._05641_ ),
    .X(\u_cpu.REG_FILE._05645_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11359_  (.A(\u_cpu.REG_FILE._05645_ ),
    .X(\u_cpu.REG_FILE._00983_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11360_  (.A0(\u_cpu.REG_FILE.rf[2][24] ),
    .A1(\u_cpu.REG_FILE._05269_ ),
    .S(\u_cpu.REG_FILE._05641_ ),
    .X(\u_cpu.REG_FILE._05646_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11361_  (.A(\u_cpu.REG_FILE._05646_ ),
    .X(\u_cpu.REG_FILE._00984_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11362_  (.A0(\u_cpu.REG_FILE.rf[2][25] ),
    .A1(\u_cpu.REG_FILE._05271_ ),
    .S(\u_cpu.REG_FILE._05641_ ),
    .X(\u_cpu.REG_FILE._05647_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11363_  (.A(\u_cpu.REG_FILE._05647_ ),
    .X(\u_cpu.REG_FILE._00985_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11364_  (.A0(\u_cpu.REG_FILE.rf[2][26] ),
    .A1(\u_cpu.REG_FILE._05273_ ),
    .S(\u_cpu.REG_FILE._05641_ ),
    .X(\u_cpu.REG_FILE._05648_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11365_  (.A(\u_cpu.REG_FILE._05648_ ),
    .X(\u_cpu.REG_FILE._00986_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11366_  (.A0(\u_cpu.REG_FILE.rf[2][27] ),
    .A1(\u_cpu.REG_FILE._05275_ ),
    .S(\u_cpu.REG_FILE._05641_ ),
    .X(\u_cpu.REG_FILE._05649_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11367_  (.A(\u_cpu.REG_FILE._05649_ ),
    .X(\u_cpu.REG_FILE._00987_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11368_  (.A0(\u_cpu.REG_FILE.rf[2][28] ),
    .A1(\u_cpu.REG_FILE._05277_ ),
    .S(\u_cpu.REG_FILE._05641_ ),
    .X(\u_cpu.REG_FILE._05650_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11369_  (.A(\u_cpu.REG_FILE._05650_ ),
    .X(\u_cpu.REG_FILE._00988_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11370_  (.A0(\u_cpu.REG_FILE.rf[2][29] ),
    .A1(\u_cpu.REG_FILE._05279_ ),
    .S(\u_cpu.REG_FILE._05641_ ),
    .X(\u_cpu.REG_FILE._05651_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11371_  (.A(\u_cpu.REG_FILE._05651_ ),
    .X(\u_cpu.REG_FILE._00989_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11372_  (.A0(\u_cpu.REG_FILE.rf[2][30] ),
    .A1(\u_cpu.REG_FILE._05281_ ),
    .S(\u_cpu.REG_FILE._05618_ ),
    .X(\u_cpu.REG_FILE._05652_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11373_  (.A(\u_cpu.REG_FILE._05652_ ),
    .X(\u_cpu.REG_FILE._00990_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11374_  (.A0(\u_cpu.REG_FILE.rf[2][31] ),
    .A1(\u_cpu.REG_FILE._05283_ ),
    .S(\u_cpu.REG_FILE._05618_ ),
    .X(\u_cpu.REG_FILE._05653_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11375_  (.A(\u_cpu.REG_FILE._05653_ ),
    .X(\u_cpu.REG_FILE._00991_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu.REG_FILE._11376_  (.A(\u_cpu.REG_FILE._04496_ ),
    .B(\u_cpu.REG_FILE._04422_ ),
    .C(\u_cpu.REG_FILE._04494_ ),
    .D(\u_cpu.REG_FILE._04747_ ),
    .X(\u_cpu.REG_FILE._05654_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11377_  (.A(\u_cpu.REG_FILE._05654_ ),
    .X(\u_cpu.REG_FILE._05655_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11378_  (.A0(\u_cpu.REG_FILE.rf[30][0] ),
    .A1(\u_cpu.REG_FILE.wd3[0] ),
    .S(\u_cpu.REG_FILE._05655_ ),
    .X(\u_cpu.REG_FILE._05656_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11379_  (.A(\u_cpu.REG_FILE._05656_ ),
    .X(\u_cpu.REG_FILE._00992_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11380_  (.A0(\u_cpu.REG_FILE.rf[30][1] ),
    .A1(\u_cpu.REG_FILE.wd3[1] ),
    .S(\u_cpu.REG_FILE._05655_ ),
    .X(\u_cpu.REG_FILE._05657_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11381_  (.A(\u_cpu.REG_FILE._05657_ ),
    .X(\u_cpu.REG_FILE._00993_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11382_  (.A0(\u_cpu.REG_FILE.rf[30][2] ),
    .A1(\u_cpu.REG_FILE.wd3[2] ),
    .S(\u_cpu.REG_FILE._05655_ ),
    .X(\u_cpu.REG_FILE._05658_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11383_  (.A(\u_cpu.REG_FILE._05658_ ),
    .X(\u_cpu.REG_FILE._00994_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11384_  (.A0(\u_cpu.REG_FILE.rf[30][3] ),
    .A1(\u_cpu.REG_FILE.wd3[3] ),
    .S(\u_cpu.REG_FILE._05655_ ),
    .X(\u_cpu.REG_FILE._05659_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11385_  (.A(\u_cpu.REG_FILE._05659_ ),
    .X(\u_cpu.REG_FILE._00995_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11386_  (.A0(\u_cpu.REG_FILE.rf[30][4] ),
    .A1(\u_cpu.REG_FILE.wd3[4] ),
    .S(\u_cpu.REG_FILE._05655_ ),
    .X(\u_cpu.REG_FILE._05660_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11387_  (.A(\u_cpu.REG_FILE._05660_ ),
    .X(\u_cpu.REG_FILE._00996_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11388_  (.A0(\u_cpu.REG_FILE.rf[30][5] ),
    .A1(\u_cpu.REG_FILE.wd3[5] ),
    .S(\u_cpu.REG_FILE._05655_ ),
    .X(\u_cpu.REG_FILE._05661_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11389_  (.A(\u_cpu.REG_FILE._05661_ ),
    .X(\u_cpu.REG_FILE._00997_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11390_  (.A0(\u_cpu.REG_FILE.rf[30][6] ),
    .A1(\u_cpu.REG_FILE.wd3[6] ),
    .S(\u_cpu.REG_FILE._05655_ ),
    .X(\u_cpu.REG_FILE._05662_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11391_  (.A(\u_cpu.REG_FILE._05662_ ),
    .X(\u_cpu.REG_FILE._00998_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11392_  (.A0(\u_cpu.REG_FILE.rf[30][7] ),
    .A1(\u_cpu.REG_FILE.wd3[7] ),
    .S(\u_cpu.REG_FILE._05655_ ),
    .X(\u_cpu.REG_FILE._05663_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11393_  (.A(\u_cpu.REG_FILE._05663_ ),
    .X(\u_cpu.REG_FILE._00999_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11394_  (.A0(\u_cpu.REG_FILE.rf[30][8] ),
    .A1(\u_cpu.REG_FILE.wd3[8] ),
    .S(\u_cpu.REG_FILE._05655_ ),
    .X(\u_cpu.REG_FILE._05664_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11395_  (.A(\u_cpu.REG_FILE._05664_ ),
    .X(\u_cpu.REG_FILE._01000_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11396_  (.A0(\u_cpu.REG_FILE.rf[30][9] ),
    .A1(\u_cpu.REG_FILE.wd3[9] ),
    .S(\u_cpu.REG_FILE._05655_ ),
    .X(\u_cpu.REG_FILE._05665_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11397_  (.A(\u_cpu.REG_FILE._05665_ ),
    .X(\u_cpu.REG_FILE._01001_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11398_  (.A(\u_cpu.REG_FILE._05654_ ),
    .X(\u_cpu.REG_FILE._05666_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11399_  (.A0(\u_cpu.REG_FILE.rf[30][10] ),
    .A1(\u_cpu.REG_FILE.wd3[10] ),
    .S(\u_cpu.REG_FILE._05666_ ),
    .X(\u_cpu.REG_FILE._05667_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11400_  (.A(\u_cpu.REG_FILE._05667_ ),
    .X(\u_cpu.REG_FILE._01002_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11401_  (.A0(\u_cpu.REG_FILE.rf[30][11] ),
    .A1(\u_cpu.REG_FILE.wd3[11] ),
    .S(\u_cpu.REG_FILE._05666_ ),
    .X(\u_cpu.REG_FILE._05668_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11402_  (.A(\u_cpu.REG_FILE._05668_ ),
    .X(\u_cpu.REG_FILE._01003_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11403_  (.A0(\u_cpu.REG_FILE.rf[30][12] ),
    .A1(\u_cpu.REG_FILE.wd3[12] ),
    .S(\u_cpu.REG_FILE._05666_ ),
    .X(\u_cpu.REG_FILE._05669_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11404_  (.A(\u_cpu.REG_FILE._05669_ ),
    .X(\u_cpu.REG_FILE._01004_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11405_  (.A0(\u_cpu.REG_FILE.rf[30][13] ),
    .A1(\u_cpu.REG_FILE.wd3[13] ),
    .S(\u_cpu.REG_FILE._05666_ ),
    .X(\u_cpu.REG_FILE._05670_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11406_  (.A(\u_cpu.REG_FILE._05670_ ),
    .X(\u_cpu.REG_FILE._01005_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11407_  (.A0(\u_cpu.REG_FILE.rf[30][14] ),
    .A1(\u_cpu.REG_FILE.wd3[14] ),
    .S(\u_cpu.REG_FILE._05666_ ),
    .X(\u_cpu.REG_FILE._05671_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11408_  (.A(\u_cpu.REG_FILE._05671_ ),
    .X(\u_cpu.REG_FILE._01006_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11409_  (.A0(\u_cpu.REG_FILE.rf[30][15] ),
    .A1(\u_cpu.REG_FILE.wd3[15] ),
    .S(\u_cpu.REG_FILE._05666_ ),
    .X(\u_cpu.REG_FILE._05672_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11410_  (.A(\u_cpu.REG_FILE._05672_ ),
    .X(\u_cpu.REG_FILE._01007_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11411_  (.A0(\u_cpu.REG_FILE.rf[30][16] ),
    .A1(\u_cpu.REG_FILE.wd3[16] ),
    .S(\u_cpu.REG_FILE._05666_ ),
    .X(\u_cpu.REG_FILE._05673_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11412_  (.A(\u_cpu.REG_FILE._05673_ ),
    .X(\u_cpu.REG_FILE._01008_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11413_  (.A0(\u_cpu.REG_FILE.rf[30][17] ),
    .A1(\u_cpu.REG_FILE.wd3[17] ),
    .S(\u_cpu.REG_FILE._05666_ ),
    .X(\u_cpu.REG_FILE._05674_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11414_  (.A(\u_cpu.REG_FILE._05674_ ),
    .X(\u_cpu.REG_FILE._01009_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11415_  (.A0(\u_cpu.REG_FILE.rf[30][18] ),
    .A1(\u_cpu.REG_FILE.wd3[18] ),
    .S(\u_cpu.REG_FILE._05666_ ),
    .X(\u_cpu.REG_FILE._05675_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11416_  (.A(\u_cpu.REG_FILE._05675_ ),
    .X(\u_cpu.REG_FILE._01010_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11417_  (.A0(\u_cpu.REG_FILE.rf[30][19] ),
    .A1(\u_cpu.REG_FILE.wd3[19] ),
    .S(\u_cpu.REG_FILE._05666_ ),
    .X(\u_cpu.REG_FILE._05676_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11418_  (.A(\u_cpu.REG_FILE._05676_ ),
    .X(\u_cpu.REG_FILE._01011_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11419_  (.A(\u_cpu.REG_FILE._05654_ ),
    .X(\u_cpu.REG_FILE._05677_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11420_  (.A0(\u_cpu.REG_FILE.rf[30][20] ),
    .A1(\u_cpu.REG_FILE.wd3[20] ),
    .S(\u_cpu.REG_FILE._05677_ ),
    .X(\u_cpu.REG_FILE._05678_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11421_  (.A(\u_cpu.REG_FILE._05678_ ),
    .X(\u_cpu.REG_FILE._01012_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11422_  (.A0(\u_cpu.REG_FILE.rf[30][21] ),
    .A1(\u_cpu.REG_FILE.wd3[21] ),
    .S(\u_cpu.REG_FILE._05677_ ),
    .X(\u_cpu.REG_FILE._05679_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11423_  (.A(\u_cpu.REG_FILE._05679_ ),
    .X(\u_cpu.REG_FILE._01013_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11424_  (.A0(\u_cpu.REG_FILE.rf[30][22] ),
    .A1(\u_cpu.REG_FILE.wd3[22] ),
    .S(\u_cpu.REG_FILE._05677_ ),
    .X(\u_cpu.REG_FILE._05680_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11425_  (.A(\u_cpu.REG_FILE._05680_ ),
    .X(\u_cpu.REG_FILE._01014_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11426_  (.A0(\u_cpu.REG_FILE.rf[30][23] ),
    .A1(\u_cpu.REG_FILE.wd3[23] ),
    .S(\u_cpu.REG_FILE._05677_ ),
    .X(\u_cpu.REG_FILE._05681_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11427_  (.A(\u_cpu.REG_FILE._05681_ ),
    .X(\u_cpu.REG_FILE._01015_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11428_  (.A0(\u_cpu.REG_FILE.rf[30][24] ),
    .A1(\u_cpu.REG_FILE.wd3[24] ),
    .S(\u_cpu.REG_FILE._05677_ ),
    .X(\u_cpu.REG_FILE._05682_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11429_  (.A(\u_cpu.REG_FILE._05682_ ),
    .X(\u_cpu.REG_FILE._01016_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11430_  (.A0(\u_cpu.REG_FILE.rf[30][25] ),
    .A1(\u_cpu.REG_FILE.wd3[25] ),
    .S(\u_cpu.REG_FILE._05677_ ),
    .X(\u_cpu.REG_FILE._05683_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11431_  (.A(\u_cpu.REG_FILE._05683_ ),
    .X(\u_cpu.REG_FILE._01017_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11432_  (.A0(\u_cpu.REG_FILE.rf[30][26] ),
    .A1(\u_cpu.REG_FILE.wd3[26] ),
    .S(\u_cpu.REG_FILE._05677_ ),
    .X(\u_cpu.REG_FILE._05684_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11433_  (.A(\u_cpu.REG_FILE._05684_ ),
    .X(\u_cpu.REG_FILE._01018_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11434_  (.A0(\u_cpu.REG_FILE.rf[30][27] ),
    .A1(\u_cpu.REG_FILE.wd3[27] ),
    .S(\u_cpu.REG_FILE._05677_ ),
    .X(\u_cpu.REG_FILE._05685_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11435_  (.A(\u_cpu.REG_FILE._05685_ ),
    .X(\u_cpu.REG_FILE._01019_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11436_  (.A0(\u_cpu.REG_FILE.rf[30][28] ),
    .A1(\u_cpu.REG_FILE.wd3[28] ),
    .S(\u_cpu.REG_FILE._05677_ ),
    .X(\u_cpu.REG_FILE._05686_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11437_  (.A(\u_cpu.REG_FILE._05686_ ),
    .X(\u_cpu.REG_FILE._01020_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11438_  (.A0(\u_cpu.REG_FILE.rf[30][29] ),
    .A1(\u_cpu.REG_FILE.wd3[29] ),
    .S(\u_cpu.REG_FILE._05677_ ),
    .X(\u_cpu.REG_FILE._05687_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11439_  (.A(\u_cpu.REG_FILE._05687_ ),
    .X(\u_cpu.REG_FILE._01021_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11440_  (.A0(\u_cpu.REG_FILE.rf[30][30] ),
    .A1(\u_cpu.REG_FILE.wd3[30] ),
    .S(\u_cpu.REG_FILE._05654_ ),
    .X(\u_cpu.REG_FILE._05688_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11441_  (.A(\u_cpu.REG_FILE._05688_ ),
    .X(\u_cpu.REG_FILE._01022_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu.REG_FILE._11442_  (.A0(\u_cpu.REG_FILE.rf[30][31] ),
    .A1(\u_cpu.REG_FILE.wd3[31] ),
    .S(\u_cpu.REG_FILE._05654_ ),
    .X(\u_cpu.REG_FILE._05689_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu.REG_FILE._11443_  (.A(\u_cpu.REG_FILE._05689_ ),
    .X(\u_cpu.REG_FILE._01023_ ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11444_  (.CLK(clknet_leaf_124_wb_clk_i),
    .D(\u_cpu.REG_FILE._00000_ ),
    .Q(\u_cpu.REG_FILE.rf[9][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11445_  (.CLK(clknet_leaf_125_wb_clk_i),
    .D(\u_cpu.REG_FILE._00001_ ),
    .Q(\u_cpu.REG_FILE.rf[9][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11446_  (.CLK(clknet_leaf_122_wb_clk_i),
    .D(\u_cpu.REG_FILE._00002_ ),
    .Q(\u_cpu.REG_FILE.rf[9][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11447_  (.CLK(clknet_leaf_115_wb_clk_i),
    .D(\u_cpu.REG_FILE._00003_ ),
    .Q(\u_cpu.REG_FILE.rf[9][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11448_  (.CLK(clknet_leaf_122_wb_clk_i),
    .D(\u_cpu.REG_FILE._00004_ ),
    .Q(\u_cpu.REG_FILE.rf[9][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11449_  (.CLK(clknet_leaf_100_wb_clk_i),
    .D(\u_cpu.REG_FILE._00005_ ),
    .Q(\u_cpu.REG_FILE.rf[9][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11450_  (.CLK(clknet_leaf_108_wb_clk_i),
    .D(\u_cpu.REG_FILE._00006_ ),
    .Q(\u_cpu.REG_FILE.rf[9][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11451_  (.CLK(clknet_leaf_115_wb_clk_i),
    .D(\u_cpu.REG_FILE._00007_ ),
    .Q(\u_cpu.REG_FILE.rf[9][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11452_  (.CLK(clknet_leaf_98_wb_clk_i),
    .D(\u_cpu.REG_FILE._00008_ ),
    .Q(\u_cpu.REG_FILE.rf[9][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11453_  (.CLK(clknet_leaf_114_wb_clk_i),
    .D(\u_cpu.REG_FILE._00009_ ),
    .Q(\u_cpu.REG_FILE.rf[9][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11454_  (.CLK(clknet_leaf_96_wb_clk_i),
    .D(\u_cpu.REG_FILE._00010_ ),
    .Q(\u_cpu.REG_FILE.rf[9][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11455_  (.CLK(clknet_leaf_102_wb_clk_i),
    .D(\u_cpu.REG_FILE._00011_ ),
    .Q(\u_cpu.REG_FILE.rf[9][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11456_  (.CLK(clknet_leaf_95_wb_clk_i),
    .D(\u_cpu.REG_FILE._00012_ ),
    .Q(\u_cpu.REG_FILE.rf[9][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11457_  (.CLK(clknet_leaf_94_wb_clk_i),
    .D(\u_cpu.REG_FILE._00013_ ),
    .Q(\u_cpu.REG_FILE.rf[9][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11458_  (.CLK(clknet_leaf_91_wb_clk_i),
    .D(\u_cpu.REG_FILE._00014_ ),
    .Q(\u_cpu.REG_FILE.rf[9][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11459_  (.CLK(clknet_leaf_102_wb_clk_i),
    .D(\u_cpu.REG_FILE._00015_ ),
    .Q(\u_cpu.REG_FILE.rf[9][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11460_  (.CLK(clknet_leaf_107_wb_clk_i),
    .D(\u_cpu.REG_FILE._00016_ ),
    .Q(\u_cpu.REG_FILE.rf[9][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11461_  (.CLK(clknet_leaf_104_wb_clk_i),
    .D(\u_cpu.REG_FILE._00017_ ),
    .Q(\u_cpu.REG_FILE.rf[9][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11462_  (.CLK(clknet_leaf_105_wb_clk_i),
    .D(\u_cpu.REG_FILE._00018_ ),
    .Q(\u_cpu.REG_FILE.rf[9][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11463_  (.CLK(clknet_leaf_107_wb_clk_i),
    .D(\u_cpu.REG_FILE._00019_ ),
    .Q(\u_cpu.REG_FILE.rf[9][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11464_  (.CLK(clknet_leaf_80_wb_clk_i),
    .D(\u_cpu.REG_FILE._00020_ ),
    .Q(\u_cpu.REG_FILE.rf[9][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11465_  (.CLK(clknet_leaf_82_wb_clk_i),
    .D(\u_cpu.REG_FILE._00021_ ),
    .Q(\u_cpu.REG_FILE.rf[9][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11466_  (.CLK(clknet_leaf_79_wb_clk_i),
    .D(\u_cpu.REG_FILE._00022_ ),
    .Q(\u_cpu.REG_FILE.rf[9][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11467_  (.CLK(clknet_leaf_79_wb_clk_i),
    .D(\u_cpu.REG_FILE._00023_ ),
    .Q(\u_cpu.REG_FILE.rf[9][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11468_  (.CLK(clknet_leaf_83_wb_clk_i),
    .D(\u_cpu.REG_FILE._00024_ ),
    .Q(\u_cpu.REG_FILE.rf[9][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11469_  (.CLK(clknet_leaf_83_wb_clk_i),
    .D(\u_cpu.REG_FILE._00025_ ),
    .Q(\u_cpu.REG_FILE.rf[9][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11470_  (.CLK(clknet_leaf_84_wb_clk_i),
    .D(\u_cpu.REG_FILE._00026_ ),
    .Q(\u_cpu.REG_FILE.rf[9][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11471_  (.CLK(clknet_leaf_86_wb_clk_i),
    .D(\u_cpu.REG_FILE._00027_ ),
    .Q(\u_cpu.REG_FILE.rf[9][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11472_  (.CLK(clknet_leaf_81_wb_clk_i),
    .D(\u_cpu.REG_FILE._00028_ ),
    .Q(\u_cpu.REG_FILE.rf[9][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11473_  (.CLK(clknet_leaf_69_wb_clk_i),
    .D(\u_cpu.REG_FILE._00029_ ),
    .Q(\u_cpu.REG_FILE.rf[9][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11474_  (.CLK(clknet_leaf_113_wb_clk_i),
    .D(\u_cpu.REG_FILE._00030_ ),
    .Q(\u_cpu.REG_FILE.rf[9][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11475_  (.CLK(clknet_leaf_75_wb_clk_i),
    .D(\u_cpu.REG_FILE._00031_ ),
    .Q(\u_cpu.REG_FILE.rf[9][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11476_  (.CLK(clknet_leaf_3_wb_clk_i),
    .D(\u_cpu.REG_FILE._00032_ ),
    .Q(\u_cpu.REG_FILE.rf[19][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11477_  (.CLK(clknet_leaf_3_wb_clk_i),
    .D(\u_cpu.REG_FILE._00033_ ),
    .Q(\u_cpu.REG_FILE.rf[19][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11478_  (.CLK(clknet_leaf_7_wb_clk_i),
    .D(\u_cpu.REG_FILE._00034_ ),
    .Q(\u_cpu.REG_FILE.rf[19][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11479_  (.CLK(clknet_leaf_113_wb_clk_i),
    .D(\u_cpu.REG_FILE._00035_ ),
    .Q(\u_cpu.REG_FILE.rf[19][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11480_  (.CLK(clknet_leaf_4_wb_clk_i),
    .D(\u_cpu.REG_FILE._00036_ ),
    .Q(\u_cpu.REG_FILE.rf[19][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11481_  (.CLK(clknet_leaf_5_wb_clk_i),
    .D(\u_cpu.REG_FILE._00037_ ),
    .Q(\u_cpu.REG_FILE.rf[19][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11482_  (.CLK(clknet_leaf_3_wb_clk_i),
    .D(\u_cpu.REG_FILE._00038_ ),
    .Q(\u_cpu.REG_FILE.rf[19][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11483_  (.CLK(clknet_leaf_117_wb_clk_i),
    .D(\u_cpu.REG_FILE._00039_ ),
    .Q(\u_cpu.REG_FILE.rf[19][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11484_  (.CLK(clknet_leaf_3_wb_clk_i),
    .D(\u_cpu.REG_FILE._00040_ ),
    .Q(\u_cpu.REG_FILE.rf[19][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11485_  (.CLK(clknet_leaf_6_wb_clk_i),
    .D(\u_cpu.REG_FILE._00041_ ),
    .Q(\u_cpu.REG_FILE.rf[19][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11486_  (.CLK(clknet_leaf_118_wb_clk_i),
    .D(\u_cpu.REG_FILE._00042_ ),
    .Q(\u_cpu.REG_FILE.rf[19][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11487_  (.CLK(clknet_leaf_38_wb_clk_i),
    .D(\u_cpu.REG_FILE._00043_ ),
    .Q(\u_cpu.REG_FILE.rf[19][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11488_  (.CLK(clknet_leaf_118_wb_clk_i),
    .D(\u_cpu.REG_FILE._00044_ ),
    .Q(\u_cpu.REG_FILE.rf[19][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11489_  (.CLK(clknet_leaf_118_wb_clk_i),
    .D(\u_cpu.REG_FILE._00045_ ),
    .Q(\u_cpu.REG_FILE.rf[19][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11490_  (.CLK(clknet_leaf_118_wb_clk_i),
    .D(\u_cpu.REG_FILE._00046_ ),
    .Q(\u_cpu.REG_FILE.rf[19][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11491_  (.CLK(clknet_leaf_37_wb_clk_i),
    .D(\u_cpu.REG_FILE._00047_ ),
    .Q(\u_cpu.REG_FILE.rf[19][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11492_  (.CLK(clknet_leaf_39_wb_clk_i),
    .D(\u_cpu.REG_FILE._00048_ ),
    .Q(\u_cpu.REG_FILE.rf[19][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11493_  (.CLK(clknet_leaf_36_wb_clk_i),
    .D(\u_cpu.REG_FILE._00049_ ),
    .Q(\u_cpu.REG_FILE.rf[19][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11494_  (.CLK(clknet_leaf_35_wb_clk_i),
    .D(\u_cpu.REG_FILE._00050_ ),
    .Q(\u_cpu.REG_FILE.rf[19][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11495_  (.CLK(clknet_leaf_41_wb_clk_i),
    .D(\u_cpu.REG_FILE._00051_ ),
    .Q(\u_cpu.REG_FILE.rf[19][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11496_  (.CLK(clknet_leaf_44_wb_clk_i),
    .D(\u_cpu.REG_FILE._00052_ ),
    .Q(\u_cpu.REG_FILE.rf[19][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11497_  (.CLK(clknet_leaf_46_wb_clk_i),
    .D(\u_cpu.REG_FILE._00053_ ),
    .Q(\u_cpu.REG_FILE.rf[19][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11498_  (.CLK(clknet_leaf_77_wb_clk_i),
    .D(\u_cpu.REG_FILE._00054_ ),
    .Q(\u_cpu.REG_FILE.rf[19][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11499_  (.CLK(clknet_leaf_46_wb_clk_i),
    .D(\u_cpu.REG_FILE._00055_ ),
    .Q(\u_cpu.REG_FILE.rf[19][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11500_  (.CLK(clknet_leaf_51_wb_clk_i),
    .D(\u_cpu.REG_FILE._00056_ ),
    .Q(\u_cpu.REG_FILE.rf[19][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11501_  (.CLK(clknet_leaf_111_wb_clk_i),
    .D(\u_cpu.REG_FILE._00057_ ),
    .Q(\u_cpu.REG_FILE.rf[19][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11502_  (.CLK(clknet_leaf_51_wb_clk_i),
    .D(\u_cpu.REG_FILE._00058_ ),
    .Q(\u_cpu.REG_FILE.rf[19][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11503_  (.CLK(clknet_leaf_46_wb_clk_i),
    .D(\u_cpu.REG_FILE._00059_ ),
    .Q(\u_cpu.REG_FILE.rf[19][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11504_  (.CLK(clknet_leaf_51_wb_clk_i),
    .D(\u_cpu.REG_FILE._00060_ ),
    .Q(\u_cpu.REG_FILE.rf[19][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11505_  (.CLK(clknet_leaf_111_wb_clk_i),
    .D(\u_cpu.REG_FILE._00061_ ),
    .Q(\u_cpu.REG_FILE.rf[19][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11506_  (.CLK(clknet_leaf_41_wb_clk_i),
    .D(\u_cpu.REG_FILE._00062_ ),
    .Q(\u_cpu.REG_FILE.rf[19][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11507_  (.CLK(clknet_leaf_112_wb_clk_i),
    .D(\u_cpu.REG_FILE._00063_ ),
    .Q(\u_cpu.REG_FILE.rf[19][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11508_  (.CLK(clknet_leaf_2_wb_clk_i),
    .D(\u_cpu.REG_FILE._00064_ ),
    .Q(\u_cpu.REG_FILE.rf[29][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11509_  (.CLK(clknet_leaf_2_wb_clk_i),
    .D(\u_cpu.REG_FILE._00065_ ),
    .Q(\u_cpu.REG_FILE.rf[29][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11510_  (.CLK(clknet_leaf_5_wb_clk_i),
    .D(\u_cpu.REG_FILE._00066_ ),
    .Q(\u_cpu.REG_FILE.rf[29][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11511_  (.CLK(clknet_leaf_10_wb_clk_i),
    .D(\u_cpu.REG_FILE._00067_ ),
    .Q(\u_cpu.REG_FILE.rf[29][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11512_  (.CLK(clknet_leaf_4_wb_clk_i),
    .D(\u_cpu.REG_FILE._00068_ ),
    .Q(\u_cpu.REG_FILE.rf[29][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11513_  (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\u_cpu.REG_FILE._00069_ ),
    .Q(\u_cpu.REG_FILE.rf[29][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11514_  (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\u_cpu.REG_FILE._00070_ ),
    .Q(\u_cpu.REG_FILE.rf[29][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11515_  (.CLK(clknet_leaf_5_wb_clk_i),
    .D(\u_cpu.REG_FILE._00071_ ),
    .Q(\u_cpu.REG_FILE.rf[29][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11516_  (.CLK(clknet_leaf_4_wb_clk_i),
    .D(\u_cpu.REG_FILE._00072_ ),
    .Q(\u_cpu.REG_FILE.rf[29][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11517_  (.CLK(clknet_leaf_6_wb_clk_i),
    .D(\u_cpu.REG_FILE._00073_ ),
    .Q(\u_cpu.REG_FILE.rf[29][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11518_  (.CLK(clknet_leaf_3_wb_clk_i),
    .D(\u_cpu.REG_FILE._00074_ ),
    .Q(\u_cpu.REG_FILE.rf[29][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11519_  (.CLK(clknet_leaf_39_wb_clk_i),
    .D(\u_cpu.REG_FILE._00075_ ),
    .Q(\u_cpu.REG_FILE.rf[29][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11520_  (.CLK(clknet_leaf_118_wb_clk_i),
    .D(\u_cpu.REG_FILE._00076_ ),
    .Q(\u_cpu.REG_FILE.rf[29][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11521_  (.CLK(clknet_leaf_118_wb_clk_i),
    .D(\u_cpu.REG_FILE._00077_ ),
    .Q(\u_cpu.REG_FILE.rf[29][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11522_  (.CLK(clknet_leaf_117_wb_clk_i),
    .D(\u_cpu.REG_FILE._00078_ ),
    .Q(\u_cpu.REG_FILE.rf[29][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11523_  (.CLK(clknet_leaf_37_wb_clk_i),
    .D(\u_cpu.REG_FILE._00079_ ),
    .Q(\u_cpu.REG_FILE.rf[29][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11524_  (.CLK(clknet_leaf_34_wb_clk_i),
    .D(\u_cpu.REG_FILE._00080_ ),
    .Q(\u_cpu.REG_FILE.rf[29][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11525_  (.CLK(clknet_leaf_37_wb_clk_i),
    .D(\u_cpu.REG_FILE._00081_ ),
    .Q(\u_cpu.REG_FILE.rf[29][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11526_  (.CLK(clknet_leaf_35_wb_clk_i),
    .D(\u_cpu.REG_FILE._00082_ ),
    .Q(\u_cpu.REG_FILE.rf[29][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11527_  (.CLK(clknet_leaf_33_wb_clk_i),
    .D(\u_cpu.REG_FILE._00083_ ),
    .Q(\u_cpu.REG_FILE.rf[29][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11528_  (.CLK(clknet_leaf_50_wb_clk_i),
    .D(\u_cpu.REG_FILE._00084_ ),
    .Q(\u_cpu.REG_FILE.rf[29][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11529_  (.CLK(clknet_leaf_76_wb_clk_i),
    .D(\u_cpu.REG_FILE._00085_ ),
    .Q(\u_cpu.REG_FILE.rf[29][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11530_  (.CLK(clknet_leaf_45_wb_clk_i),
    .D(\u_cpu.REG_FILE._00086_ ),
    .Q(\u_cpu.REG_FILE.rf[29][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11531_  (.CLK(clknet_leaf_48_wb_clk_i),
    .D(\u_cpu.REG_FILE._00087_ ),
    .Q(\u_cpu.REG_FILE.rf[29][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11532_  (.CLK(clknet_leaf_52_wb_clk_i),
    .D(\u_cpu.REG_FILE._00088_ ),
    .Q(\u_cpu.REG_FILE.rf[29][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11533_  (.CLK(clknet_leaf_43_wb_clk_i),
    .D(\u_cpu.REG_FILE._00089_ ),
    .Q(\u_cpu.REG_FILE.rf[29][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11534_  (.CLK(clknet_leaf_50_wb_clk_i),
    .D(\u_cpu.REG_FILE._00090_ ),
    .Q(\u_cpu.REG_FILE.rf[29][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11535_  (.CLK(clknet_leaf_34_wb_clk_i),
    .D(\u_cpu.REG_FILE._00091_ ),
    .Q(\u_cpu.REG_FILE.rf[29][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11536_  (.CLK(clknet_leaf_51_wb_clk_i),
    .D(\u_cpu.REG_FILE._00092_ ),
    .Q(\u_cpu.REG_FILE.rf[29][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11537_  (.CLK(clknet_leaf_43_wb_clk_i),
    .D(\u_cpu.REG_FILE._00093_ ),
    .Q(\u_cpu.REG_FILE.rf[29][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11538_  (.CLK(clknet_leaf_42_wb_clk_i),
    .D(\u_cpu.REG_FILE._00094_ ),
    .Q(\u_cpu.REG_FILE.rf[29][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11539_  (.CLK(clknet_leaf_42_wb_clk_i),
    .D(\u_cpu.REG_FILE._00095_ ),
    .Q(\u_cpu.REG_FILE.rf[29][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11540_  (.CLK(clknet_leaf_2_wb_clk_i),
    .D(\u_cpu.REG_FILE._00096_ ),
    .Q(\u_cpu.REG_FILE.rf[31][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11541_  (.CLK(clknet_leaf_2_wb_clk_i),
    .D(\u_cpu.REG_FILE._00097_ ),
    .Q(\u_cpu.REG_FILE.rf[31][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11542_  (.CLK(clknet_leaf_4_wb_clk_i),
    .D(\u_cpu.REG_FILE._00098_ ),
    .Q(\u_cpu.REG_FILE.rf[31][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11543_  (.CLK(clknet_leaf_9_wb_clk_i),
    .D(\u_cpu.REG_FILE._00099_ ),
    .Q(\u_cpu.REG_FILE.rf[31][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11544_  (.CLK(clknet_leaf_4_wb_clk_i),
    .D(\u_cpu.REG_FILE._00100_ ),
    .Q(\u_cpu.REG_FILE.rf[31][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11545_  (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\u_cpu.REG_FILE._00101_ ),
    .Q(\u_cpu.REG_FILE.rf[31][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11546_  (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\u_cpu.REG_FILE._00102_ ),
    .Q(\u_cpu.REG_FILE.rf[31][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11547_  (.CLK(clknet_leaf_8_wb_clk_i),
    .D(\u_cpu.REG_FILE._00103_ ),
    .Q(\u_cpu.REG_FILE.rf[31][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11548_  (.CLK(clknet_leaf_117_wb_clk_i),
    .D(\u_cpu.REG_FILE._00104_ ),
    .Q(\u_cpu.REG_FILE.rf[31][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11549_  (.CLK(clknet_leaf_6_wb_clk_i),
    .D(\u_cpu.REG_FILE._00105_ ),
    .Q(\u_cpu.REG_FILE.rf[31][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11550_  (.CLK(clknet_leaf_3_wb_clk_i),
    .D(\u_cpu.REG_FILE._00106_ ),
    .Q(\u_cpu.REG_FILE.rf[31][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11551_  (.CLK(clknet_leaf_39_wb_clk_i),
    .D(\u_cpu.REG_FILE._00107_ ),
    .Q(\u_cpu.REG_FILE.rf[31][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11552_  (.CLK(clknet_leaf_117_wb_clk_i),
    .D(\u_cpu.REG_FILE._00108_ ),
    .Q(\u_cpu.REG_FILE.rf[31][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11553_  (.CLK(clknet_leaf_4_wb_clk_i),
    .D(\u_cpu.REG_FILE._00109_ ),
    .Q(\u_cpu.REG_FILE.rf[31][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11554_  (.CLK(clknet_leaf_117_wb_clk_i),
    .D(\u_cpu.REG_FILE._00110_ ),
    .Q(\u_cpu.REG_FILE.rf[31][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11555_  (.CLK(clknet_leaf_27_wb_clk_i),
    .D(\u_cpu.REG_FILE._00111_ ),
    .Q(\u_cpu.REG_FILE.rf[31][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11556_  (.CLK(clknet_leaf_34_wb_clk_i),
    .D(\u_cpu.REG_FILE._00112_ ),
    .Q(\u_cpu.REG_FILE.rf[31][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11557_  (.CLK(clknet_leaf_37_wb_clk_i),
    .D(\u_cpu.REG_FILE._00113_ ),
    .Q(\u_cpu.REG_FILE.rf[31][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11558_  (.CLK(clknet_leaf_35_wb_clk_i),
    .D(\u_cpu.REG_FILE._00114_ ),
    .Q(\u_cpu.REG_FILE.rf[31][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11559_  (.CLK(clknet_leaf_32_wb_clk_i),
    .D(\u_cpu.REG_FILE._00115_ ),
    .Q(\u_cpu.REG_FILE.rf[31][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11560_  (.CLK(clknet_leaf_50_wb_clk_i),
    .D(\u_cpu.REG_FILE._00116_ ),
    .Q(\u_cpu.REG_FILE.rf[31][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11561_  (.CLK(clknet_leaf_43_wb_clk_i),
    .D(\u_cpu.REG_FILE._00117_ ),
    .Q(\u_cpu.REG_FILE.rf[31][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11562_  (.CLK(clknet_leaf_45_wb_clk_i),
    .D(\u_cpu.REG_FILE._00118_ ),
    .Q(\u_cpu.REG_FILE.rf[31][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11563_  (.CLK(clknet_leaf_48_wb_clk_i),
    .D(\u_cpu.REG_FILE._00119_ ),
    .Q(\u_cpu.REG_FILE.rf[31][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11564_  (.CLK(clknet_leaf_52_wb_clk_i),
    .D(\u_cpu.REG_FILE._00120_ ),
    .Q(\u_cpu.REG_FILE.rf[31][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11565_  (.CLK(clknet_leaf_40_wb_clk_i),
    .D(\u_cpu.REG_FILE._00121_ ),
    .Q(\u_cpu.REG_FILE.rf[31][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11566_  (.CLK(clknet_leaf_50_wb_clk_i),
    .D(\u_cpu.REG_FILE._00122_ ),
    .Q(\u_cpu.REG_FILE.rf[31][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11567_  (.CLK(clknet_leaf_34_wb_clk_i),
    .D(\u_cpu.REG_FILE._00123_ ),
    .Q(\u_cpu.REG_FILE.rf[31][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11568_  (.CLK(clknet_leaf_52_wb_clk_i),
    .D(\u_cpu.REG_FILE._00124_ ),
    .Q(\u_cpu.REG_FILE.rf[31][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11569_  (.CLK(clknet_leaf_43_wb_clk_i),
    .D(\u_cpu.REG_FILE._00125_ ),
    .Q(\u_cpu.REG_FILE.rf[31][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11570_  (.CLK(clknet_leaf_42_wb_clk_i),
    .D(\u_cpu.REG_FILE._00126_ ),
    .Q(\u_cpu.REG_FILE.rf[31][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11571_  (.CLK(clknet_leaf_41_wb_clk_i),
    .D(\u_cpu.REG_FILE._00127_ ),
    .Q(\u_cpu.REG_FILE.rf[31][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11572_  (.CLK(clknet_leaf_126_wb_clk_i),
    .D(\u_cpu.REG_FILE._00128_ ),
    .Q(\u_cpu.REG_FILE.rf[3][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11573_  (.CLK(clknet_leaf_127_wb_clk_i),
    .D(\u_cpu.REG_FILE._00129_ ),
    .Q(\u_cpu.REG_FILE.rf[3][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11574_  (.CLK(clknet_leaf_120_wb_clk_i),
    .D(\u_cpu.REG_FILE._00130_ ),
    .Q(\u_cpu.REG_FILE.rf[3][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11575_  (.CLK(clknet_leaf_117_wb_clk_i),
    .D(\u_cpu.REG_FILE._00131_ ),
    .Q(\u_cpu.REG_FILE.rf[3][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11576_  (.CLK(clknet_leaf_120_wb_clk_i),
    .D(\u_cpu.REG_FILE._00132_ ),
    .Q(\u_cpu.REG_FILE.rf[3][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11577_  (.CLK(clknet_leaf_122_wb_clk_i),
    .D(\u_cpu.REG_FILE._00133_ ),
    .Q(\u_cpu.REG_FILE.rf[3][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11578_  (.CLK(clknet_leaf_127_wb_clk_i),
    .D(\u_cpu.REG_FILE._00134_ ),
    .Q(\u_cpu.REG_FILE.rf[3][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11579_  (.CLK(clknet_leaf_7_wb_clk_i),
    .D(\u_cpu.REG_FILE._00135_ ),
    .Q(\u_cpu.REG_FILE.rf[3][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11580_  (.CLK(clknet_leaf_124_wb_clk_i),
    .D(\u_cpu.REG_FILE._00136_ ),
    .Q(\u_cpu.REG_FILE.rf[3][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11581_  (.CLK(clknet_leaf_8_wb_clk_i),
    .D(\u_cpu.REG_FILE._00137_ ),
    .Q(\u_cpu.REG_FILE.rf[3][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11582_  (.CLK(clknet_leaf_99_wb_clk_i),
    .D(\u_cpu.REG_FILE._00138_ ),
    .Q(\u_cpu.REG_FILE.rf[3][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11583_  (.CLK(clknet_leaf_111_wb_clk_i),
    .D(\u_cpu.REG_FILE._00139_ ),
    .Q(\u_cpu.REG_FILE.rf[3][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11584_  (.CLK(clknet_leaf_93_wb_clk_i),
    .D(\u_cpu.REG_FILE._00140_ ),
    .Q(\u_cpu.REG_FILE.rf[3][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11585_  (.CLK(clknet_leaf_94_wb_clk_i),
    .D(\u_cpu.REG_FILE._00141_ ),
    .Q(\u_cpu.REG_FILE.rf[3][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11586_  (.CLK(clknet_leaf_91_wb_clk_i),
    .D(\u_cpu.REG_FILE._00142_ ),
    .Q(\u_cpu.REG_FILE.rf[3][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11587_  (.CLK(clknet_leaf_102_wb_clk_i),
    .D(\u_cpu.REG_FILE._00143_ ),
    .Q(\u_cpu.REG_FILE.rf[3][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11588_  (.CLK(clknet_leaf_108_wb_clk_i),
    .D(\u_cpu.REG_FILE._00144_ ),
    .Q(\u_cpu.REG_FILE.rf[3][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11589_  (.CLK(clknet_leaf_105_wb_clk_i),
    .D(\u_cpu.REG_FILE._00145_ ),
    .Q(\u_cpu.REG_FILE.rf[3][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11590_  (.CLK(clknet_leaf_49_wb_clk_i),
    .D(\u_cpu.REG_FILE._00146_ ),
    .Q(\u_cpu.REG_FILE.rf[3][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11591_  (.CLK(clknet_leaf_43_wb_clk_i),
    .D(\u_cpu.REG_FILE._00147_ ),
    .Q(\u_cpu.REG_FILE.rf[3][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11592_  (.CLK(clknet_leaf_75_wb_clk_i),
    .D(\u_cpu.REG_FILE._00148_ ),
    .Q(\u_cpu.REG_FILE.rf[3][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11593_  (.CLK(clknet_leaf_73_wb_clk_i),
    .D(\u_cpu.REG_FILE._00149_ ),
    .Q(\u_cpu.REG_FILE.rf[3][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11594_  (.CLK(clknet_leaf_47_wb_clk_i),
    .D(\u_cpu.REG_FILE._00150_ ),
    .Q(\u_cpu.REG_FILE.rf[3][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11595_  (.CLK(clknet_leaf_73_wb_clk_i),
    .D(\u_cpu.REG_FILE._00151_ ),
    .Q(\u_cpu.REG_FILE.rf[3][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11596_  (.CLK(clknet_leaf_72_wb_clk_i),
    .D(\u_cpu.REG_FILE._00152_ ),
    .Q(\u_cpu.REG_FILE.rf[3][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11597_  (.CLK(clknet_leaf_74_wb_clk_i),
    .D(\u_cpu.REG_FILE._00153_ ),
    .Q(\u_cpu.REG_FILE.rf[3][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11598_  (.CLK(clknet_leaf_49_wb_clk_i),
    .D(\u_cpu.REG_FILE._00154_ ),
    .Q(\u_cpu.REG_FILE.rf[3][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11599_  (.CLK(clknet_leaf_49_wb_clk_i),
    .D(\u_cpu.REG_FILE._00155_ ),
    .Q(\u_cpu.REG_FILE.rf[3][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11600_  (.CLK(clknet_leaf_74_wb_clk_i),
    .D(\u_cpu.REG_FILE._00156_ ),
    .Q(\u_cpu.REG_FILE.rf[3][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11601_  (.CLK(clknet_leaf_74_wb_clk_i),
    .D(\u_cpu.REG_FILE._00157_ ),
    .Q(\u_cpu.REG_FILE.rf[3][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11602_  (.CLK(clknet_leaf_9_wb_clk_i),
    .D(\u_cpu.REG_FILE._00158_ ),
    .Q(\u_cpu.REG_FILE.rf[3][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11603_  (.CLK(clknet_leaf_73_wb_clk_i),
    .D(\u_cpu.REG_FILE._00159_ ),
    .Q(\u_cpu.REG_FILE.rf[3][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11604_  (.CLK(clknet_leaf_124_wb_clk_i),
    .D(\u_cpu.REG_FILE._00160_ ),
    .Q(\u_cpu.REG_FILE.rf[4][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11605_  (.CLK(clknet_leaf_126_wb_clk_i),
    .D(\u_cpu.REG_FILE._00161_ ),
    .Q(\u_cpu.REG_FILE.rf[4][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11606_  (.CLK(clknet_leaf_123_wb_clk_i),
    .D(\u_cpu.REG_FILE._00162_ ),
    .Q(\u_cpu.REG_FILE.rf[4][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11607_  (.CLK(clknet_leaf_114_wb_clk_i),
    .D(\u_cpu.REG_FILE._00163_ ),
    .Q(\u_cpu.REG_FILE.rf[4][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11608_  (.CLK(clknet_leaf_122_wb_clk_i),
    .D(\u_cpu.REG_FILE._00164_ ),
    .Q(\u_cpu.REG_FILE.rf[4][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11609_  (.CLK(clknet_leaf_100_wb_clk_i),
    .D(\u_cpu.REG_FILE._00165_ ),
    .Q(\u_cpu.REG_FILE.rf[4][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11610_  (.CLK(clknet_leaf_99_wb_clk_i),
    .D(\u_cpu.REG_FILE._00166_ ),
    .Q(\u_cpu.REG_FILE.rf[4][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11611_  (.CLK(clknet_leaf_113_wb_clk_i),
    .D(\u_cpu.REG_FILE._00167_ ),
    .Q(\u_cpu.REG_FILE.rf[4][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11612_  (.CLK(clknet_leaf_96_wb_clk_i),
    .D(\u_cpu.REG_FILE._00168_ ),
    .Q(\u_cpu.REG_FILE.rf[4][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11613_  (.CLK(clknet_leaf_112_wb_clk_i),
    .D(\u_cpu.REG_FILE._00169_ ),
    .Q(\u_cpu.REG_FILE.rf[4][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11614_  (.CLK(clknet_leaf_96_wb_clk_i),
    .D(\u_cpu.REG_FILE._00170_ ),
    .Q(\u_cpu.REG_FILE.rf[4][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11615_  (.CLK(clknet_leaf_78_wb_clk_i),
    .D(\u_cpu.REG_FILE._00171_ ),
    .Q(\u_cpu.REG_FILE.rf[4][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11616_  (.CLK(clknet_leaf_93_wb_clk_i),
    .D(\u_cpu.REG_FILE._00172_ ),
    .Q(\u_cpu.REG_FILE.rf[4][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11617_  (.CLK(clknet_leaf_94_wb_clk_i),
    .D(\u_cpu.REG_FILE._00173_ ),
    .Q(\u_cpu.REG_FILE.rf[4][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11618_  (.CLK(clknet_leaf_91_wb_clk_i),
    .D(\u_cpu.REG_FILE._00174_ ),
    .Q(\u_cpu.REG_FILE.rf[4][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11619_  (.CLK(clknet_leaf_103_wb_clk_i),
    .D(\u_cpu.REG_FILE._00175_ ),
    .Q(\u_cpu.REG_FILE.rf[4][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11620_  (.CLK(clknet_leaf_107_wb_clk_i),
    .D(\u_cpu.REG_FILE._00176_ ),
    .Q(\u_cpu.REG_FILE.rf[4][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11621_  (.CLK(clknet_leaf_103_wb_clk_i),
    .D(\u_cpu.REG_FILE._00177_ ),
    .Q(\u_cpu.REG_FILE.rf[4][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11622_  (.CLK(clknet_leaf_90_wb_clk_i),
    .D(\u_cpu.REG_FILE._00178_ ),
    .Q(\u_cpu.REG_FILE.rf[4][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11623_  (.CLK(clknet_leaf_78_wb_clk_i),
    .D(\u_cpu.REG_FILE._00179_ ),
    .Q(\u_cpu.REG_FILE.rf[4][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11624_  (.CLK(clknet_leaf_75_wb_clk_i),
    .D(\u_cpu.REG_FILE._00180_ ),
    .Q(\u_cpu.REG_FILE.rf[4][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11625_  (.CLK(clknet_leaf_73_wb_clk_i),
    .D(\u_cpu.REG_FILE._00181_ ),
    .Q(\u_cpu.REG_FILE.rf[4][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11626_  (.CLK(clknet_leaf_72_wb_clk_i),
    .D(\u_cpu.REG_FILE._00182_ ),
    .Q(\u_cpu.REG_FILE.rf[4][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11627_  (.CLK(clknet_leaf_73_wb_clk_i),
    .D(\u_cpu.REG_FILE._00183_ ),
    .Q(\u_cpu.REG_FILE.rf[4][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11628_  (.CLK(clknet_leaf_70_wb_clk_i),
    .D(\u_cpu.REG_FILE._00184_ ),
    .Q(\u_cpu.REG_FILE.rf[4][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11629_  (.CLK(clknet_leaf_70_wb_clk_i),
    .D(\u_cpu.REG_FILE._00185_ ),
    .Q(\u_cpu.REG_FILE.rf[4][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11630_  (.CLK(clknet_leaf_71_wb_clk_i),
    .D(\u_cpu.REG_FILE._00186_ ),
    .Q(\u_cpu.REG_FILE.rf[4][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11631_  (.CLK(clknet_leaf_70_wb_clk_i),
    .D(\u_cpu.REG_FILE._00187_ ),
    .Q(\u_cpu.REG_FILE.rf[4][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11632_  (.CLK(clknet_leaf_69_wb_clk_i),
    .D(\u_cpu.REG_FILE._00188_ ),
    .Q(\u_cpu.REG_FILE.rf[4][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11633_  (.CLK(clknet_leaf_69_wb_clk_i),
    .D(\u_cpu.REG_FILE._00189_ ),
    .Q(\u_cpu.REG_FILE.rf[4][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11634_  (.CLK(clknet_leaf_111_wb_clk_i),
    .D(\u_cpu.REG_FILE._00190_ ),
    .Q(\u_cpu.REG_FILE.rf[4][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11635_  (.CLK(clknet_leaf_74_wb_clk_i),
    .D(\u_cpu.REG_FILE._00191_ ),
    .Q(\u_cpu.REG_FILE.rf[4][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11636_  (.CLK(clknet_leaf_126_wb_clk_i),
    .D(\u_cpu.REG_FILE._00192_ ),
    .Q(\u_cpu.REG_FILE.rf[5][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11637_  (.CLK(clknet_leaf_126_wb_clk_i),
    .D(\u_cpu.REG_FILE._00193_ ),
    .Q(\u_cpu.REG_FILE.rf[5][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11638_  (.CLK(clknet_leaf_123_wb_clk_i),
    .D(\u_cpu.REG_FILE._00194_ ),
    .Q(\u_cpu.REG_FILE.rf[5][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11639_  (.CLK(clknet_leaf_117_wb_clk_i),
    .D(\u_cpu.REG_FILE._00195_ ),
    .Q(\u_cpu.REG_FILE.rf[5][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11640_  (.CLK(clknet_leaf_120_wb_clk_i),
    .D(\u_cpu.REG_FILE._00196_ ),
    .Q(\u_cpu.REG_FILE.rf[5][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11641_  (.CLK(clknet_leaf_100_wb_clk_i),
    .D(\u_cpu.REG_FILE._00197_ ),
    .Q(\u_cpu.REG_FILE.rf[5][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11642_  (.CLK(clknet_leaf_98_wb_clk_i),
    .D(\u_cpu.REG_FILE._00198_ ),
    .Q(\u_cpu.REG_FILE.rf[5][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11643_  (.CLK(clknet_leaf_114_wb_clk_i),
    .D(\u_cpu.REG_FILE._00199_ ),
    .Q(\u_cpu.REG_FILE.rf[5][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11644_  (.CLK(clknet_leaf_98_wb_clk_i),
    .D(\u_cpu.REG_FILE._00200_ ),
    .Q(\u_cpu.REG_FILE.rf[5][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11645_  (.CLK(clknet_leaf_113_wb_clk_i),
    .D(\u_cpu.REG_FILE._00201_ ),
    .Q(\u_cpu.REG_FILE.rf[5][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11646_  (.CLK(clknet_leaf_99_wb_clk_i),
    .D(\u_cpu.REG_FILE._00202_ ),
    .Q(\u_cpu.REG_FILE.rf[5][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11647_  (.CLK(clknet_leaf_78_wb_clk_i),
    .D(\u_cpu.REG_FILE._00203_ ),
    .Q(\u_cpu.REG_FILE.rf[5][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11648_  (.CLK(clknet_leaf_95_wb_clk_i),
    .D(\u_cpu.REG_FILE._00204_ ),
    .Q(\u_cpu.REG_FILE.rf[5][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11649_  (.CLK(clknet_leaf_94_wb_clk_i),
    .D(\u_cpu.REG_FILE._00205_ ),
    .Q(\u_cpu.REG_FILE.rf[5][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11650_  (.CLK(clknet_leaf_91_wb_clk_i),
    .D(\u_cpu.REG_FILE._00206_ ),
    .Q(\u_cpu.REG_FILE.rf[5][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11651_  (.CLK(clknet_leaf_102_wb_clk_i),
    .D(\u_cpu.REG_FILE._00207_ ),
    .Q(\u_cpu.REG_FILE.rf[5][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11652_  (.CLK(clknet_leaf_109_wb_clk_i),
    .D(\u_cpu.REG_FILE._00208_ ),
    .Q(\u_cpu.REG_FILE.rf[5][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11653_  (.CLK(clknet_leaf_103_wb_clk_i),
    .D(\u_cpu.REG_FILE._00209_ ),
    .Q(\u_cpu.REG_FILE.rf[5][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11654_  (.CLK(clknet_leaf_90_wb_clk_i),
    .D(\u_cpu.REG_FILE._00210_ ),
    .Q(\u_cpu.REG_FILE.rf[5][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11655_  (.CLK(clknet_leaf_110_wb_clk_i),
    .D(\u_cpu.REG_FILE._00211_ ),
    .Q(\u_cpu.REG_FILE.rf[5][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11656_  (.CLK(clknet_leaf_75_wb_clk_i),
    .D(\u_cpu.REG_FILE._00212_ ),
    .Q(\u_cpu.REG_FILE.rf[5][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11657_  (.CLK(clknet_leaf_73_wb_clk_i),
    .D(\u_cpu.REG_FILE._00213_ ),
    .Q(\u_cpu.REG_FILE.rf[5][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11658_  (.CLK(clknet_leaf_72_wb_clk_i),
    .D(\u_cpu.REG_FILE._00214_ ),
    .Q(\u_cpu.REG_FILE.rf[5][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11659_  (.CLK(clknet_leaf_76_wb_clk_i),
    .D(\u_cpu.REG_FILE._00215_ ),
    .Q(\u_cpu.REG_FILE.rf[5][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11660_  (.CLK(clknet_leaf_74_wb_clk_i),
    .D(\u_cpu.REG_FILE._00216_ ),
    .Q(\u_cpu.REG_FILE.rf[5][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11661_  (.CLK(clknet_leaf_69_wb_clk_i),
    .D(\u_cpu.REG_FILE._00217_ ),
    .Q(\u_cpu.REG_FILE.rf[5][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11662_  (.CLK(clknet_leaf_71_wb_clk_i),
    .D(\u_cpu.REG_FILE._00218_ ),
    .Q(\u_cpu.REG_FILE.rf[5][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11663_  (.CLK(clknet_leaf_71_wb_clk_i),
    .D(\u_cpu.REG_FILE._00219_ ),
    .Q(\u_cpu.REG_FILE.rf[5][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11664_  (.CLK(clknet_leaf_74_wb_clk_i),
    .D(\u_cpu.REG_FILE._00220_ ),
    .Q(\u_cpu.REG_FILE.rf[5][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11665_  (.CLK(clknet_leaf_69_wb_clk_i),
    .D(\u_cpu.REG_FILE._00221_ ),
    .Q(\u_cpu.REG_FILE.rf[5][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11666_  (.CLK(clknet_leaf_112_wb_clk_i),
    .D(\u_cpu.REG_FILE._00222_ ),
    .Q(\u_cpu.REG_FILE.rf[5][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11667_  (.CLK(clknet_leaf_74_wb_clk_i),
    .D(\u_cpu.REG_FILE._00223_ ),
    .Q(\u_cpu.REG_FILE.rf[5][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11668_  (.CLK(clknet_leaf_123_wb_clk_i),
    .D(\u_cpu.REG_FILE._00224_ ),
    .Q(\u_cpu.REG_FILE.rf[6][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11669_  (.CLK(clknet_leaf_123_wb_clk_i),
    .D(\u_cpu.REG_FILE._00225_ ),
    .Q(\u_cpu.REG_FILE.rf[6][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11670_  (.CLK(clknet_leaf_123_wb_clk_i),
    .D(\u_cpu.REG_FILE._00226_ ),
    .Q(\u_cpu.REG_FILE.rf[6][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11671_  (.CLK(clknet_leaf_121_wb_clk_i),
    .D(\u_cpu.REG_FILE._00227_ ),
    .Q(\u_cpu.REG_FILE.rf[6][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11672_  (.CLK(clknet_leaf_121_wb_clk_i),
    .D(\u_cpu.REG_FILE._00228_ ),
    .Q(\u_cpu.REG_FILE.rf[6][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11673_  (.CLK(clknet_leaf_101_wb_clk_i),
    .D(\u_cpu.REG_FILE._00229_ ),
    .Q(\u_cpu.REG_FILE.rf[6][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11674_  (.CLK(clknet_leaf_122_wb_clk_i),
    .D(\u_cpu.REG_FILE._00230_ ),
    .Q(\u_cpu.REG_FILE.rf[6][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11675_  (.CLK(clknet_leaf_113_wb_clk_i),
    .D(\u_cpu.REG_FILE._00231_ ),
    .Q(\u_cpu.REG_FILE.rf[6][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11676_  (.CLK(clknet_leaf_99_wb_clk_i),
    .D(\u_cpu.REG_FILE._00232_ ),
    .Q(\u_cpu.REG_FILE.rf[6][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11677_  (.CLK(clknet_leaf_113_wb_clk_i),
    .D(\u_cpu.REG_FILE._00233_ ),
    .Q(\u_cpu.REG_FILE.rf[6][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11678_  (.CLK(clknet_leaf_96_wb_clk_i),
    .D(\u_cpu.REG_FILE._00234_ ),
    .Q(\u_cpu.REG_FILE.rf[6][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11679_  (.CLK(clknet_leaf_78_wb_clk_i),
    .D(\u_cpu.REG_FILE._00235_ ),
    .Q(\u_cpu.REG_FILE.rf[6][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11680_  (.CLK(clknet_leaf_93_wb_clk_i),
    .D(\u_cpu.REG_FILE._00236_ ),
    .Q(\u_cpu.REG_FILE.rf[6][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11681_  (.CLK(clknet_leaf_92_wb_clk_i),
    .D(\u_cpu.REG_FILE._00237_ ),
    .Q(\u_cpu.REG_FILE.rf[6][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11682_  (.CLK(clknet_leaf_92_wb_clk_i),
    .D(\u_cpu.REG_FILE._00238_ ),
    .Q(\u_cpu.REG_FILE.rf[6][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11683_  (.CLK(clknet_leaf_103_wb_clk_i),
    .D(\u_cpu.REG_FILE._00239_ ),
    .Q(\u_cpu.REG_FILE.rf[6][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11684_  (.CLK(clknet_leaf_109_wb_clk_i),
    .D(\u_cpu.REG_FILE._00240_ ),
    .Q(\u_cpu.REG_FILE.rf[6][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11685_  (.CLK(clknet_leaf_103_wb_clk_i),
    .D(\u_cpu.REG_FILE._00241_ ),
    .Q(\u_cpu.REG_FILE.rf[6][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11686_  (.CLK(clknet_leaf_105_wb_clk_i),
    .D(\u_cpu.REG_FILE._00242_ ),
    .Q(\u_cpu.REG_FILE.rf[6][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11687_  (.CLK(clknet_leaf_110_wb_clk_i),
    .D(\u_cpu.REG_FILE._00243_ ),
    .Q(\u_cpu.REG_FILE.rf[6][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11688_  (.CLK(clknet_leaf_75_wb_clk_i),
    .D(\u_cpu.REG_FILE._00244_ ),
    .Q(\u_cpu.REG_FILE.rf[6][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11689_  (.CLK(clknet_leaf_73_wb_clk_i),
    .D(\u_cpu.REG_FILE._00245_ ),
    .Q(\u_cpu.REG_FILE.rf[6][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11690_  (.CLK(clknet_leaf_72_wb_clk_i),
    .D(\u_cpu.REG_FILE._00246_ ),
    .Q(\u_cpu.REG_FILE.rf[6][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11691_  (.CLK(clknet_leaf_75_wb_clk_i),
    .D(\u_cpu.REG_FILE._00247_ ),
    .Q(\u_cpu.REG_FILE.rf[6][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11692_  (.CLK(clknet_leaf_70_wb_clk_i),
    .D(\u_cpu.REG_FILE._00248_ ),
    .Q(\u_cpu.REG_FILE.rf[6][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11693_  (.CLK(clknet_leaf_70_wb_clk_i),
    .D(\u_cpu.REG_FILE._00249_ ),
    .Q(\u_cpu.REG_FILE.rf[6][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11694_  (.CLK(clknet_leaf_70_wb_clk_i),
    .D(\u_cpu.REG_FILE._00250_ ),
    .Q(\u_cpu.REG_FILE.rf[6][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11695_  (.CLK(clknet_leaf_70_wb_clk_i),
    .D(\u_cpu.REG_FILE._00251_ ),
    .Q(\u_cpu.REG_FILE.rf[6][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11696_  (.CLK(clknet_leaf_69_wb_clk_i),
    .D(\u_cpu.REG_FILE._00252_ ),
    .Q(\u_cpu.REG_FILE.rf[6][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11697_  (.CLK(clknet_leaf_68_wb_clk_i),
    .D(\u_cpu.REG_FILE._00253_ ),
    .Q(\u_cpu.REG_FILE.rf[6][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11698_  (.CLK(clknet_leaf_111_wb_clk_i),
    .D(\u_cpu.REG_FILE._00254_ ),
    .Q(\u_cpu.REG_FILE.rf[6][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11699_  (.CLK(clknet_leaf_75_wb_clk_i),
    .D(\u_cpu.REG_FILE._00255_ ),
    .Q(\u_cpu.REG_FILE.rf[6][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11700_  (.CLK(clknet_leaf_126_wb_clk_i),
    .D(\u_cpu.REG_FILE._00256_ ),
    .Q(\u_cpu.REG_FILE.rf[7][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11701_  (.CLK(clknet_leaf_126_wb_clk_i),
    .D(\u_cpu.REG_FILE._00257_ ),
    .Q(\u_cpu.REG_FILE.rf[7][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11702_  (.CLK(clknet_leaf_123_wb_clk_i),
    .D(\u_cpu.REG_FILE._00258_ ),
    .Q(\u_cpu.REG_FILE.rf[7][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11703_  (.CLK(clknet_leaf_121_wb_clk_i),
    .D(\u_cpu.REG_FILE._00259_ ),
    .Q(\u_cpu.REG_FILE.rf[7][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11704_  (.CLK(clknet_leaf_121_wb_clk_i),
    .D(\u_cpu.REG_FILE._00260_ ),
    .Q(\u_cpu.REG_FILE.rf[7][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11705_  (.CLK(clknet_leaf_100_wb_clk_i),
    .D(\u_cpu.REG_FILE._00261_ ),
    .Q(\u_cpu.REG_FILE.rf[7][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11706_  (.CLK(clknet_leaf_124_wb_clk_i),
    .D(\u_cpu.REG_FILE._00262_ ),
    .Q(\u_cpu.REG_FILE.rf[7][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11707_  (.CLK(clknet_leaf_113_wb_clk_i),
    .D(\u_cpu.REG_FILE._00263_ ),
    .Q(\u_cpu.REG_FILE.rf[7][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11708_  (.CLK(clknet_leaf_97_wb_clk_i),
    .D(\u_cpu.REG_FILE._00264_ ),
    .Q(\u_cpu.REG_FILE.rf[7][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11709_  (.CLK(clknet_leaf_113_wb_clk_i),
    .D(\u_cpu.REG_FILE._00265_ ),
    .Q(\u_cpu.REG_FILE.rf[7][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11710_  (.CLK(clknet_leaf_96_wb_clk_i),
    .D(\u_cpu.REG_FILE._00266_ ),
    .Q(\u_cpu.REG_FILE.rf[7][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11711_  (.CLK(clknet_leaf_110_wb_clk_i),
    .D(\u_cpu.REG_FILE._00267_ ),
    .Q(\u_cpu.REG_FILE.rf[7][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11712_  (.CLK(clknet_leaf_93_wb_clk_i),
    .D(\u_cpu.REG_FILE._00268_ ),
    .Q(\u_cpu.REG_FILE.rf[7][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11713_  (.CLK(clknet_leaf_94_wb_clk_i),
    .D(\u_cpu.REG_FILE._00269_ ),
    .Q(\u_cpu.REG_FILE.rf[7][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11714_  (.CLK(clknet_leaf_92_wb_clk_i),
    .D(\u_cpu.REG_FILE._00270_ ),
    .Q(\u_cpu.REG_FILE.rf[7][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11715_  (.CLK(clknet_leaf_103_wb_clk_i),
    .D(\u_cpu.REG_FILE._00271_ ),
    .Q(\u_cpu.REG_FILE.rf[7][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11716_  (.CLK(clknet_leaf_109_wb_clk_i),
    .D(\u_cpu.REG_FILE._00272_ ),
    .Q(\u_cpu.REG_FILE.rf[7][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11717_  (.CLK(clknet_leaf_103_wb_clk_i),
    .D(\u_cpu.REG_FILE._00273_ ),
    .Q(\u_cpu.REG_FILE.rf[7][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11718_  (.CLK(clknet_leaf_83_wb_clk_i),
    .D(\u_cpu.REG_FILE._00274_ ),
    .Q(\u_cpu.REG_FILE.rf[7][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11719_  (.CLK(clknet_leaf_110_wb_clk_i),
    .D(\u_cpu.REG_FILE._00275_ ),
    .Q(\u_cpu.REG_FILE.rf[7][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11720_  (.CLK(clknet_leaf_75_wb_clk_i),
    .D(\u_cpu.REG_FILE._00276_ ),
    .Q(\u_cpu.REG_FILE.rf[7][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11721_  (.CLK(clknet_leaf_73_wb_clk_i),
    .D(\u_cpu.REG_FILE._00277_ ),
    .Q(\u_cpu.REG_FILE.rf[7][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11722_  (.CLK(clknet_leaf_72_wb_clk_i),
    .D(\u_cpu.REG_FILE._00278_ ),
    .Q(\u_cpu.REG_FILE.rf[7][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11723_  (.CLK(clknet_leaf_75_wb_clk_i),
    .D(\u_cpu.REG_FILE._00279_ ),
    .Q(\u_cpu.REG_FILE.rf[7][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11724_  (.CLK(clknet_leaf_71_wb_clk_i),
    .D(\u_cpu.REG_FILE._00280_ ),
    .Q(\u_cpu.REG_FILE.rf[7][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11725_  (.CLK(clknet_leaf_70_wb_clk_i),
    .D(\u_cpu.REG_FILE._00281_ ),
    .Q(\u_cpu.REG_FILE.rf[7][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11726_  (.CLK(clknet_leaf_70_wb_clk_i),
    .D(\u_cpu.REG_FILE._00282_ ),
    .Q(\u_cpu.REG_FILE.rf[7][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11727_  (.CLK(clknet_leaf_70_wb_clk_i),
    .D(\u_cpu.REG_FILE._00283_ ),
    .Q(\u_cpu.REG_FILE.rf[7][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11728_  (.CLK(clknet_leaf_69_wb_clk_i),
    .D(\u_cpu.REG_FILE._00284_ ),
    .Q(\u_cpu.REG_FILE.rf[7][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11729_  (.CLK(clknet_leaf_68_wb_clk_i),
    .D(\u_cpu.REG_FILE._00285_ ),
    .Q(\u_cpu.REG_FILE.rf[7][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11730_  (.CLK(clknet_leaf_111_wb_clk_i),
    .D(\u_cpu.REG_FILE._00286_ ),
    .Q(\u_cpu.REG_FILE.rf[7][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11731_  (.CLK(clknet_leaf_75_wb_clk_i),
    .D(\u_cpu.REG_FILE._00287_ ),
    .Q(\u_cpu.REG_FILE.rf[7][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11732_  (.CLK(clknet_leaf_125_wb_clk_i),
    .D(\u_cpu.REG_FILE._00288_ ),
    .Q(\u_cpu.REG_FILE.rf[8][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11733_  (.CLK(clknet_leaf_98_wb_clk_i),
    .D(\u_cpu.REG_FILE._00289_ ),
    .Q(\u_cpu.REG_FILE.rf[8][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11734_  (.CLK(clknet_leaf_124_wb_clk_i),
    .D(\u_cpu.REG_FILE._00290_ ),
    .Q(\u_cpu.REG_FILE.rf[8][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11735_  (.CLK(clknet_leaf_116_wb_clk_i),
    .D(\u_cpu.REG_FILE._00291_ ),
    .Q(\u_cpu.REG_FILE.rf[8][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11736_  (.CLK(clknet_leaf_122_wb_clk_i),
    .D(\u_cpu.REG_FILE._00292_ ),
    .Q(\u_cpu.REG_FILE.rf[8][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11737_  (.CLK(clknet_leaf_99_wb_clk_i),
    .D(\u_cpu.REG_FILE._00293_ ),
    .Q(\u_cpu.REG_FILE.rf[8][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11738_  (.CLK(clknet_leaf_101_wb_clk_i),
    .D(\u_cpu.REG_FILE._00294_ ),
    .Q(\u_cpu.REG_FILE.rf[8][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11739_  (.CLK(clknet_leaf_115_wb_clk_i),
    .D(\u_cpu.REG_FILE._00295_ ),
    .Q(\u_cpu.REG_FILE.rf[8][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11740_  (.CLK(clknet_leaf_97_wb_clk_i),
    .D(\u_cpu.REG_FILE._00296_ ),
    .Q(\u_cpu.REG_FILE.rf[8][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11741_  (.CLK(clknet_leaf_115_wb_clk_i),
    .D(\u_cpu.REG_FILE._00297_ ),
    .Q(\u_cpu.REG_FILE.rf[8][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11742_  (.CLK(clknet_leaf_96_wb_clk_i),
    .D(\u_cpu.REG_FILE._00298_ ),
    .Q(\u_cpu.REG_FILE.rf[8][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11743_  (.CLK(clknet_leaf_107_wb_clk_i),
    .D(\u_cpu.REG_FILE._00299_ ),
    .Q(\u_cpu.REG_FILE.rf[8][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11744_  (.CLK(clknet_leaf_95_wb_clk_i),
    .D(\u_cpu.REG_FILE._00300_ ),
    .Q(\u_cpu.REG_FILE.rf[8][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11745_  (.CLK(clknet_leaf_94_wb_clk_i),
    .D(\u_cpu.REG_FILE._00301_ ),
    .Q(\u_cpu.REG_FILE.rf[8][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11746_  (.CLK(clknet_leaf_104_wb_clk_i),
    .D(\u_cpu.REG_FILE._00302_ ),
    .Q(\u_cpu.REG_FILE.rf[8][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11747_  (.CLK(clknet_leaf_103_wb_clk_i),
    .D(\u_cpu.REG_FILE._00303_ ),
    .Q(\u_cpu.REG_FILE.rf[8][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11748_  (.CLK(clknet_leaf_107_wb_clk_i),
    .D(\u_cpu.REG_FILE._00304_ ),
    .Q(\u_cpu.REG_FILE.rf[8][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11749_  (.CLK(clknet_leaf_91_wb_clk_i),
    .D(\u_cpu.REG_FILE._00305_ ),
    .Q(\u_cpu.REG_FILE.rf[8][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11750_  (.CLK(clknet_leaf_105_wb_clk_i),
    .D(\u_cpu.REG_FILE._00306_ ),
    .Q(\u_cpu.REG_FILE.rf[8][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11751_  (.CLK(clknet_leaf_107_wb_clk_i),
    .D(\u_cpu.REG_FILE._00307_ ),
    .Q(\u_cpu.REG_FILE.rf[8][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11752_  (.CLK(clknet_leaf_75_wb_clk_i),
    .D(\u_cpu.REG_FILE._00308_ ),
    .Q(\u_cpu.REG_FILE.rf[8][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11753_  (.CLK(clknet_leaf_82_wb_clk_i),
    .D(\u_cpu.REG_FILE._00309_ ),
    .Q(\u_cpu.REG_FILE.rf[8][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11754_  (.CLK(clknet_leaf_81_wb_clk_i),
    .D(\u_cpu.REG_FILE._00310_ ),
    .Q(\u_cpu.REG_FILE.rf[8][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11755_  (.CLK(clknet_leaf_79_wb_clk_i),
    .D(\u_cpu.REG_FILE._00311_ ),
    .Q(\u_cpu.REG_FILE.rf[8][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11756_  (.CLK(clknet_leaf_83_wb_clk_i),
    .D(\u_cpu.REG_FILE._00312_ ),
    .Q(\u_cpu.REG_FILE.rf[8][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11757_  (.CLK(clknet_leaf_84_wb_clk_i),
    .D(\u_cpu.REG_FILE._00313_ ),
    .Q(\u_cpu.REG_FILE.rf[8][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11758_  (.CLK(clknet_leaf_84_wb_clk_i),
    .D(\u_cpu.REG_FILE._00314_ ),
    .Q(\u_cpu.REG_FILE.rf[8][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11759_  (.CLK(clknet_leaf_86_wb_clk_i),
    .D(\u_cpu.REG_FILE._00315_ ),
    .Q(\u_cpu.REG_FILE.rf[8][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11760_  (.CLK(clknet_leaf_85_wb_clk_i),
    .D(\u_cpu.REG_FILE._00316_ ),
    .Q(\u_cpu.REG_FILE.rf[8][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11761_  (.CLK(clknet_leaf_86_wb_clk_i),
    .D(\u_cpu.REG_FILE._00317_ ),
    .Q(\u_cpu.REG_FILE.rf[8][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11762_  (.CLK(clknet_leaf_114_wb_clk_i),
    .D(\u_cpu.REG_FILE._00318_ ),
    .Q(\u_cpu.REG_FILE.rf[8][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11763_  (.CLK(clknet_leaf_75_wb_clk_i),
    .D(\u_cpu.REG_FILE._00319_ ),
    .Q(\u_cpu.REG_FILE.rf[8][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11764_  (.CLK(clknet_leaf_126_wb_clk_i),
    .D(\u_cpu.REG_FILE._00320_ ),
    .Q(\u_cpu.REG_FILE.rf[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11765_  (.CLK(clknet_leaf_126_wb_clk_i),
    .D(\u_cpu.REG_FILE._00321_ ),
    .Q(\u_cpu.REG_FILE.rf[0][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11766_  (.CLK(clknet_leaf_120_wb_clk_i),
    .D(\u_cpu.REG_FILE._00322_ ),
    .Q(\u_cpu.REG_FILE.rf[0][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11767_  (.CLK(clknet_leaf_121_wb_clk_i),
    .D(\u_cpu.REG_FILE._00323_ ),
    .Q(\u_cpu.REG_FILE.rf[0][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11768_  (.CLK(clknet_leaf_120_wb_clk_i),
    .D(\u_cpu.REG_FILE._00324_ ),
    .Q(\u_cpu.REG_FILE.rf[0][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11769_  (.CLK(clknet_leaf_122_wb_clk_i),
    .D(\u_cpu.REG_FILE._00325_ ),
    .Q(\u_cpu.REG_FILE.rf[0][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11770_  (.CLK(clknet_leaf_126_wb_clk_i),
    .D(\u_cpu.REG_FILE._00326_ ),
    .Q(\u_cpu.REG_FILE.rf[0][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11771_  (.CLK(clknet_leaf_8_wb_clk_i),
    .D(\u_cpu.REG_FILE._00327_ ),
    .Q(\u_cpu.REG_FILE.rf[0][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11772_  (.CLK(clknet_leaf_99_wb_clk_i),
    .D(\u_cpu.REG_FILE._00328_ ),
    .Q(\u_cpu.REG_FILE.rf[0][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11773_  (.CLK(clknet_leaf_9_wb_clk_i),
    .D(\u_cpu.REG_FILE._00329_ ),
    .Q(\u_cpu.REG_FILE.rf[0][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11774_  (.CLK(clknet_leaf_96_wb_clk_i),
    .D(\u_cpu.REG_FILE._00330_ ),
    .Q(\u_cpu.REG_FILE.rf[0][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11775_  (.CLK(clknet_leaf_110_wb_clk_i),
    .D(\u_cpu.REG_FILE._00331_ ),
    .Q(\u_cpu.REG_FILE.rf[0][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11776_  (.CLK(clknet_leaf_93_wb_clk_i),
    .D(\u_cpu.REG_FILE._00332_ ),
    .Q(\u_cpu.REG_FILE.rf[0][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11777_  (.CLK(clknet_leaf_92_wb_clk_i),
    .D(\u_cpu.REG_FILE._00333_ ),
    .Q(\u_cpu.REG_FILE.rf[0][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11778_  (.CLK(clknet_leaf_91_wb_clk_i),
    .D(\u_cpu.REG_FILE._00334_ ),
    .Q(\u_cpu.REG_FILE.rf[0][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11779_  (.CLK(clknet_leaf_102_wb_clk_i),
    .D(\u_cpu.REG_FILE._00335_ ),
    .Q(\u_cpu.REG_FILE.rf[0][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11780_  (.CLK(clknet_leaf_110_wb_clk_i),
    .D(\u_cpu.REG_FILE._00336_ ),
    .Q(\u_cpu.REG_FILE.rf[0][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11781_  (.CLK(clknet_leaf_104_wb_clk_i),
    .D(\u_cpu.REG_FILE._00337_ ),
    .Q(\u_cpu.REG_FILE.rf[0][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11782_  (.CLK(clknet_leaf_71_wb_clk_i),
    .D(\u_cpu.REG_FILE._00338_ ),
    .Q(\u_cpu.REG_FILE.rf[0][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11783_  (.CLK(clknet_leaf_44_wb_clk_i),
    .D(\u_cpu.REG_FILE._00339_ ),
    .Q(\u_cpu.REG_FILE.rf[0][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11784_  (.CLK(clknet_leaf_76_wb_clk_i),
    .D(\u_cpu.REG_FILE._00340_ ),
    .Q(\u_cpu.REG_FILE.rf[0][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11785_  (.CLK(clknet_leaf_73_wb_clk_i),
    .D(\u_cpu.REG_FILE._00341_ ),
    .Q(\u_cpu.REG_FILE.rf[0][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11786_  (.CLK(clknet_leaf_72_wb_clk_i),
    .D(\u_cpu.REG_FILE._00342_ ),
    .Q(\u_cpu.REG_FILE.rf[0][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11787_  (.CLK(clknet_leaf_75_wb_clk_i),
    .D(\u_cpu.REG_FILE._00343_ ),
    .Q(\u_cpu.REG_FILE.rf[0][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11788_  (.CLK(clknet_leaf_71_wb_clk_i),
    .D(\u_cpu.REG_FILE._00344_ ),
    .Q(\u_cpu.REG_FILE.rf[0][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11789_  (.CLK(clknet_leaf_70_wb_clk_i),
    .D(\u_cpu.REG_FILE._00345_ ),
    .Q(\u_cpu.REG_FILE.rf[0][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11790_  (.CLK(clknet_leaf_71_wb_clk_i),
    .D(\u_cpu.REG_FILE._00346_ ),
    .Q(\u_cpu.REG_FILE.rf[0][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11791_  (.CLK(clknet_leaf_71_wb_clk_i),
    .D(\u_cpu.REG_FILE._00347_ ),
    .Q(\u_cpu.REG_FILE.rf[0][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11792_  (.CLK(clknet_leaf_80_wb_clk_i),
    .D(\u_cpu.REG_FILE._00348_ ),
    .Q(\u_cpu.REG_FILE.rf[0][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11793_  (.CLK(clknet_leaf_69_wb_clk_i),
    .D(\u_cpu.REG_FILE._00349_ ),
    .Q(\u_cpu.REG_FILE.rf[0][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11794_  (.CLK(clknet_leaf_112_wb_clk_i),
    .D(\u_cpu.REG_FILE._00350_ ),
    .Q(\u_cpu.REG_FILE.rf[0][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11795_  (.CLK(clknet_leaf_74_wb_clk_i),
    .D(\u_cpu.REG_FILE._00351_ ),
    .Q(\u_cpu.REG_FILE.rf[0][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11796_  (.CLK(clknet_leaf_125_wb_clk_i),
    .D(\u_cpu.REG_FILE._00352_ ),
    .Q(\u_cpu.REG_FILE.rf[10][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11797_  (.CLK(clknet_leaf_98_wb_clk_i),
    .D(\u_cpu.REG_FILE._00353_ ),
    .Q(\u_cpu.REG_FILE.rf[10][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11798_  (.CLK(clknet_leaf_124_wb_clk_i),
    .D(\u_cpu.REG_FILE._00354_ ),
    .Q(\u_cpu.REG_FILE.rf[10][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11799_  (.CLK(clknet_leaf_121_wb_clk_i),
    .D(\u_cpu.REG_FILE._00355_ ),
    .Q(\u_cpu.REG_FILE.rf[10][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11800_  (.CLK(clknet_leaf_122_wb_clk_i),
    .D(\u_cpu.REG_FILE._00356_ ),
    .Q(\u_cpu.REG_FILE.rf[10][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11801_  (.CLK(clknet_leaf_100_wb_clk_i),
    .D(\u_cpu.REG_FILE._00357_ ),
    .Q(\u_cpu.REG_FILE.rf[10][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11802_  (.CLK(clknet_leaf_101_wb_clk_i),
    .D(\u_cpu.REG_FILE._00358_ ),
    .Q(\u_cpu.REG_FILE.rf[10][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11803_  (.CLK(clknet_leaf_115_wb_clk_i),
    .D(\u_cpu.REG_FILE._00359_ ),
    .Q(\u_cpu.REG_FILE.rf[10][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11804_  (.CLK(clknet_leaf_97_wb_clk_i),
    .D(\u_cpu.REG_FILE._00360_ ),
    .Q(\u_cpu.REG_FILE.rf[10][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11805_  (.CLK(clknet_leaf_115_wb_clk_i),
    .D(\u_cpu.REG_FILE._00361_ ),
    .Q(\u_cpu.REG_FILE.rf[10][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11806_  (.CLK(clknet_leaf_97_wb_clk_i),
    .D(\u_cpu.REG_FILE._00362_ ),
    .Q(\u_cpu.REG_FILE.rf[10][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11807_  (.CLK(clknet_leaf_107_wb_clk_i),
    .D(\u_cpu.REG_FILE._00363_ ),
    .Q(\u_cpu.REG_FILE.rf[10][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11808_  (.CLK(clknet_leaf_95_wb_clk_i),
    .D(\u_cpu.REG_FILE._00364_ ),
    .Q(\u_cpu.REG_FILE.rf[10][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11809_  (.CLK(clknet_leaf_94_wb_clk_i),
    .D(\u_cpu.REG_FILE._00365_ ),
    .Q(\u_cpu.REG_FILE.rf[10][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11810_  (.CLK(clknet_leaf_104_wb_clk_i),
    .D(\u_cpu.REG_FILE._00366_ ),
    .Q(\u_cpu.REG_FILE.rf[10][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11811_  (.CLK(clknet_leaf_103_wb_clk_i),
    .D(\u_cpu.REG_FILE._00367_ ),
    .Q(\u_cpu.REG_FILE.rf[10][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11812_  (.CLK(clknet_leaf_107_wb_clk_i),
    .D(\u_cpu.REG_FILE._00368_ ),
    .Q(\u_cpu.REG_FILE.rf[10][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11813_  (.CLK(clknet_leaf_92_wb_clk_i),
    .D(\u_cpu.REG_FILE._00369_ ),
    .Q(\u_cpu.REG_FILE.rf[10][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11814_  (.CLK(clknet_leaf_105_wb_clk_i),
    .D(\u_cpu.REG_FILE._00370_ ),
    .Q(\u_cpu.REG_FILE.rf[10][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11815_  (.CLK(clknet_leaf_106_wb_clk_i),
    .D(\u_cpu.REG_FILE._00371_ ),
    .Q(\u_cpu.REG_FILE.rf[10][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11816_  (.CLK(clknet_leaf_80_wb_clk_i),
    .D(\u_cpu.REG_FILE._00372_ ),
    .Q(\u_cpu.REG_FILE.rf[10][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11817_  (.CLK(clknet_leaf_82_wb_clk_i),
    .D(\u_cpu.REG_FILE._00373_ ),
    .Q(\u_cpu.REG_FILE.rf[10][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11818_  (.CLK(clknet_leaf_81_wb_clk_i),
    .D(\u_cpu.REG_FILE._00374_ ),
    .Q(\u_cpu.REG_FILE.rf[10][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11819_  (.CLK(clknet_leaf_80_wb_clk_i),
    .D(\u_cpu.REG_FILE._00375_ ),
    .Q(\u_cpu.REG_FILE.rf[10][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11820_  (.CLK(clknet_leaf_82_wb_clk_i),
    .D(\u_cpu.REG_FILE._00376_ ),
    .Q(\u_cpu.REG_FILE.rf[10][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11821_  (.CLK(clknet_leaf_84_wb_clk_i),
    .D(\u_cpu.REG_FILE._00377_ ),
    .Q(\u_cpu.REG_FILE.rf[10][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11822_  (.CLK(clknet_leaf_84_wb_clk_i),
    .D(\u_cpu.REG_FILE._00378_ ),
    .Q(\u_cpu.REG_FILE.rf[10][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11823_  (.CLK(clknet_leaf_86_wb_clk_i),
    .D(\u_cpu.REG_FILE._00379_ ),
    .Q(\u_cpu.REG_FILE.rf[10][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11824_  (.CLK(clknet_leaf_81_wb_clk_i),
    .D(\u_cpu.REG_FILE._00380_ ),
    .Q(\u_cpu.REG_FILE.rf[10][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11825_  (.CLK(clknet_leaf_86_wb_clk_i),
    .D(\u_cpu.REG_FILE._00381_ ),
    .Q(\u_cpu.REG_FILE.rf[10][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11826_  (.CLK(clknet_leaf_113_wb_clk_i),
    .D(\u_cpu.REG_FILE._00382_ ),
    .Q(\u_cpu.REG_FILE.rf[10][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11827_  (.CLK(clknet_leaf_80_wb_clk_i),
    .D(\u_cpu.REG_FILE._00383_ ),
    .Q(\u_cpu.REG_FILE.rf[10][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11828_  (.CLK(clknet_leaf_124_wb_clk_i),
    .D(\u_cpu.REG_FILE._00384_ ),
    .Q(\u_cpu.REG_FILE.rf[11][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11829_  (.CLK(clknet_leaf_124_wb_clk_i),
    .D(\u_cpu.REG_FILE._00385_ ),
    .Q(\u_cpu.REG_FILE.rf[11][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11830_  (.CLK(clknet_leaf_124_wb_clk_i),
    .D(\u_cpu.REG_FILE._00386_ ),
    .Q(\u_cpu.REG_FILE.rf[11][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11831_  (.CLK(clknet_leaf_116_wb_clk_i),
    .D(\u_cpu.REG_FILE._00387_ ),
    .Q(\u_cpu.REG_FILE.rf[11][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11832_  (.CLK(clknet_leaf_123_wb_clk_i),
    .D(\u_cpu.REG_FILE._00388_ ),
    .Q(\u_cpu.REG_FILE.rf[11][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11833_  (.CLK(clknet_leaf_100_wb_clk_i),
    .D(\u_cpu.REG_FILE._00389_ ),
    .Q(\u_cpu.REG_FILE.rf[11][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11834_  (.CLK(clknet_leaf_108_wb_clk_i),
    .D(\u_cpu.REG_FILE._00390_ ),
    .Q(\u_cpu.REG_FILE.rf[11][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11835_  (.CLK(clknet_leaf_115_wb_clk_i),
    .D(\u_cpu.REG_FILE._00391_ ),
    .Q(\u_cpu.REG_FILE.rf[11][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11836_  (.CLK(clknet_leaf_98_wb_clk_i),
    .D(\u_cpu.REG_FILE._00392_ ),
    .Q(\u_cpu.REG_FILE.rf[11][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11837_  (.CLK(clknet_leaf_114_wb_clk_i),
    .D(\u_cpu.REG_FILE._00393_ ),
    .Q(\u_cpu.REG_FILE.rf[11][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11838_  (.CLK(clknet_leaf_96_wb_clk_i),
    .D(\u_cpu.REG_FILE._00394_ ),
    .Q(\u_cpu.REG_FILE.rf[11][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11839_  (.CLK(clknet_leaf_107_wb_clk_i),
    .D(\u_cpu.REG_FILE._00395_ ),
    .Q(\u_cpu.REG_FILE.rf[11][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11840_  (.CLK(clknet_leaf_96_wb_clk_i),
    .D(\u_cpu.REG_FILE._00396_ ),
    .Q(\u_cpu.REG_FILE.rf[11][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11841_  (.CLK(clknet_leaf_95_wb_clk_i),
    .D(\u_cpu.REG_FILE._00397_ ),
    .Q(\u_cpu.REG_FILE.rf[11][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11842_  (.CLK(clknet_leaf_104_wb_clk_i),
    .D(\u_cpu.REG_FILE._00398_ ),
    .Q(\u_cpu.REG_FILE.rf[11][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11843_  (.CLK(clknet_leaf_102_wb_clk_i),
    .D(\u_cpu.REG_FILE._00399_ ),
    .Q(\u_cpu.REG_FILE.rf[11][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11844_  (.CLK(clknet_leaf_107_wb_clk_i),
    .D(\u_cpu.REG_FILE._00400_ ),
    .Q(\u_cpu.REG_FILE.rf[11][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11845_  (.CLK(clknet_leaf_92_wb_clk_i),
    .D(\u_cpu.REG_FILE._00401_ ),
    .Q(\u_cpu.REG_FILE.rf[11][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11846_  (.CLK(clknet_leaf_105_wb_clk_i),
    .D(\u_cpu.REG_FILE._00402_ ),
    .Q(\u_cpu.REG_FILE.rf[11][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11847_  (.CLK(clknet_leaf_109_wb_clk_i),
    .D(\u_cpu.REG_FILE._00403_ ),
    .Q(\u_cpu.REG_FILE.rf[11][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11848_  (.CLK(clknet_leaf_79_wb_clk_i),
    .D(\u_cpu.REG_FILE._00404_ ),
    .Q(\u_cpu.REG_FILE.rf[11][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11849_  (.CLK(clknet_leaf_82_wb_clk_i),
    .D(\u_cpu.REG_FILE._00405_ ),
    .Q(\u_cpu.REG_FILE.rf[11][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11850_  (.CLK(clknet_leaf_82_wb_clk_i),
    .D(\u_cpu.REG_FILE._00406_ ),
    .Q(\u_cpu.REG_FILE.rf[11][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11851_  (.CLK(clknet_leaf_79_wb_clk_i),
    .D(\u_cpu.REG_FILE._00407_ ),
    .Q(\u_cpu.REG_FILE.rf[11][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11852_  (.CLK(clknet_leaf_82_wb_clk_i),
    .D(\u_cpu.REG_FILE._00408_ ),
    .Q(\u_cpu.REG_FILE.rf[11][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11853_  (.CLK(clknet_leaf_83_wb_clk_i),
    .D(\u_cpu.REG_FILE._00409_ ),
    .Q(\u_cpu.REG_FILE.rf[11][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11854_  (.CLK(clknet_leaf_84_wb_clk_i),
    .D(\u_cpu.REG_FILE._00410_ ),
    .Q(\u_cpu.REG_FILE.rf[11][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11855_  (.CLK(clknet_leaf_80_wb_clk_i),
    .D(\u_cpu.REG_FILE._00411_ ),
    .Q(\u_cpu.REG_FILE.rf[11][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11856_  (.CLK(clknet_leaf_81_wb_clk_i),
    .D(\u_cpu.REG_FILE._00412_ ),
    .Q(\u_cpu.REG_FILE.rf[11][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11857_  (.CLK(clknet_leaf_69_wb_clk_i),
    .D(\u_cpu.REG_FILE._00413_ ),
    .Q(\u_cpu.REG_FILE.rf[11][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11858_  (.CLK(clknet_leaf_112_wb_clk_i),
    .D(\u_cpu.REG_FILE._00414_ ),
    .Q(\u_cpu.REG_FILE.rf[11][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11859_  (.CLK(clknet_leaf_75_wb_clk_i),
    .D(\u_cpu.REG_FILE._00415_ ),
    .Q(\u_cpu.REG_FILE.rf[11][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11860_  (.CLK(clknet_leaf_125_wb_clk_i),
    .D(\u_cpu.REG_FILE._00416_ ),
    .Q(\u_cpu.REG_FILE.rf[12][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11861_  (.CLK(clknet_leaf_125_wb_clk_i),
    .D(\u_cpu.REG_FILE._00417_ ),
    .Q(\u_cpu.REG_FILE.rf[12][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11862_  (.CLK(clknet_leaf_123_wb_clk_i),
    .D(\u_cpu.REG_FILE._00418_ ),
    .Q(\u_cpu.REG_FILE.rf[12][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11863_  (.CLK(clknet_leaf_116_wb_clk_i),
    .D(\u_cpu.REG_FILE._00419_ ),
    .Q(\u_cpu.REG_FILE.rf[12][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11864_  (.CLK(clknet_leaf_121_wb_clk_i),
    .D(\u_cpu.REG_FILE._00420_ ),
    .Q(\u_cpu.REG_FILE.rf[12][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11865_  (.CLK(clknet_leaf_100_wb_clk_i),
    .D(\u_cpu.REG_FILE._00421_ ),
    .Q(\u_cpu.REG_FILE.rf[12][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11866_  (.CLK(clknet_leaf_115_wb_clk_i),
    .D(\u_cpu.REG_FILE._00422_ ),
    .Q(\u_cpu.REG_FILE.rf[12][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11867_  (.CLK(clknet_leaf_108_wb_clk_i),
    .D(\u_cpu.REG_FILE._00423_ ),
    .Q(\u_cpu.REG_FILE.rf[12][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11868_  (.CLK(clknet_leaf_98_wb_clk_i),
    .D(\u_cpu.REG_FILE._00424_ ),
    .Q(\u_cpu.REG_FILE.rf[12][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11869_  (.CLK(clknet_leaf_114_wb_clk_i),
    .D(\u_cpu.REG_FILE._00425_ ),
    .Q(\u_cpu.REG_FILE.rf[12][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11870_  (.CLK(clknet_leaf_96_wb_clk_i),
    .D(\u_cpu.REG_FILE._00426_ ),
    .Q(\u_cpu.REG_FILE.rf[12][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11871_  (.CLK(clknet_leaf_108_wb_clk_i),
    .D(\u_cpu.REG_FILE._00427_ ),
    .Q(\u_cpu.REG_FILE.rf[12][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11872_  (.CLK(clknet_leaf_95_wb_clk_i),
    .D(\u_cpu.REG_FILE._00428_ ),
    .Q(\u_cpu.REG_FILE.rf[12][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11873_  (.CLK(clknet_leaf_94_wb_clk_i),
    .D(\u_cpu.REG_FILE._00429_ ),
    .Q(\u_cpu.REG_FILE.rf[12][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11874_  (.CLK(clknet_leaf_90_wb_clk_i),
    .D(\u_cpu.REG_FILE._00430_ ),
    .Q(\u_cpu.REG_FILE.rf[12][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11875_  (.CLK(clknet_leaf_102_wb_clk_i),
    .D(\u_cpu.REG_FILE._00431_ ),
    .Q(\u_cpu.REG_FILE.rf[12][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11876_  (.CLK(clknet_leaf_108_wb_clk_i),
    .D(\u_cpu.REG_FILE._00432_ ),
    .Q(\u_cpu.REG_FILE.rf[12][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11877_  (.CLK(clknet_leaf_105_wb_clk_i),
    .D(\u_cpu.REG_FILE._00433_ ),
    .Q(\u_cpu.REG_FILE.rf[12][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11878_  (.CLK(clknet_leaf_90_wb_clk_i),
    .D(\u_cpu.REG_FILE._00434_ ),
    .Q(\u_cpu.REG_FILE.rf[12][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11879_  (.CLK(clknet_leaf_107_wb_clk_i),
    .D(\u_cpu.REG_FILE._00435_ ),
    .Q(\u_cpu.REG_FILE.rf[12][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11880_  (.CLK(clknet_leaf_79_wb_clk_i),
    .D(\u_cpu.REG_FILE._00436_ ),
    .Q(\u_cpu.REG_FILE.rf[12][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11881_  (.CLK(clknet_leaf_106_wb_clk_i),
    .D(\u_cpu.REG_FILE._00437_ ),
    .Q(\u_cpu.REG_FILE.rf[12][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11882_  (.CLK(clknet_leaf_81_wb_clk_i),
    .D(\u_cpu.REG_FILE._00438_ ),
    .Q(\u_cpu.REG_FILE.rf[12][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11883_  (.CLK(clknet_leaf_79_wb_clk_i),
    .D(\u_cpu.REG_FILE._00439_ ),
    .Q(\u_cpu.REG_FILE.rf[12][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11884_  (.CLK(clknet_leaf_82_wb_clk_i),
    .D(\u_cpu.REG_FILE._00440_ ),
    .Q(\u_cpu.REG_FILE.rf[12][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11885_  (.CLK(clknet_leaf_84_wb_clk_i),
    .D(\u_cpu.REG_FILE._00441_ ),
    .Q(\u_cpu.REG_FILE.rf[12][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11886_  (.CLK(clknet_leaf_84_wb_clk_i),
    .D(\u_cpu.REG_FILE._00442_ ),
    .Q(\u_cpu.REG_FILE.rf[12][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11887_  (.CLK(clknet_leaf_86_wb_clk_i),
    .D(\u_cpu.REG_FILE._00443_ ),
    .Q(\u_cpu.REG_FILE.rf[12][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11888_  (.CLK(clknet_leaf_81_wb_clk_i),
    .D(\u_cpu.REG_FILE._00444_ ),
    .Q(\u_cpu.REG_FILE.rf[12][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11889_  (.CLK(clknet_leaf_86_wb_clk_i),
    .D(\u_cpu.REG_FILE._00445_ ),
    .Q(\u_cpu.REG_FILE.rf[12][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11890_  (.CLK(clknet_leaf_110_wb_clk_i),
    .D(\u_cpu.REG_FILE._00446_ ),
    .Q(\u_cpu.REG_FILE.rf[12][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11891_  (.CLK(clknet_leaf_80_wb_clk_i),
    .D(\u_cpu.REG_FILE._00447_ ),
    .Q(\u_cpu.REG_FILE.rf[12][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11892_  (.CLK(clknet_leaf_125_wb_clk_i),
    .D(\u_cpu.REG_FILE._00448_ ),
    .Q(\u_cpu.REG_FILE.rf[13][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11893_  (.CLK(clknet_leaf_125_wb_clk_i),
    .D(\u_cpu.REG_FILE._00449_ ),
    .Q(\u_cpu.REG_FILE.rf[13][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11894_  (.CLK(clknet_leaf_124_wb_clk_i),
    .D(\u_cpu.REG_FILE._00450_ ),
    .Q(\u_cpu.REG_FILE.rf[13][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11895_  (.CLK(clknet_leaf_116_wb_clk_i),
    .D(\u_cpu.REG_FILE._00451_ ),
    .Q(\u_cpu.REG_FILE.rf[13][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11896_  (.CLK(clknet_leaf_121_wb_clk_i),
    .D(\u_cpu.REG_FILE._00452_ ),
    .Q(\u_cpu.REG_FILE.rf[13][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11897_  (.CLK(clknet_leaf_100_wb_clk_i),
    .D(\u_cpu.REG_FILE._00453_ ),
    .Q(\u_cpu.REG_FILE.rf[13][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11898_  (.CLK(clknet_leaf_116_wb_clk_i),
    .D(\u_cpu.REG_FILE._00454_ ),
    .Q(\u_cpu.REG_FILE.rf[13][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11899_  (.CLK(clknet_leaf_108_wb_clk_i),
    .D(\u_cpu.REG_FILE._00455_ ),
    .Q(\u_cpu.REG_FILE.rf[13][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11900_  (.CLK(clknet_leaf_97_wb_clk_i),
    .D(\u_cpu.REG_FILE._00456_ ),
    .Q(\u_cpu.REG_FILE.rf[13][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11901_  (.CLK(clknet_leaf_115_wb_clk_i),
    .D(\u_cpu.REG_FILE._00457_ ),
    .Q(\u_cpu.REG_FILE.rf[13][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11902_  (.CLK(clknet_leaf_97_wb_clk_i),
    .D(\u_cpu.REG_FILE._00458_ ),
    .Q(\u_cpu.REG_FILE.rf[13][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11903_  (.CLK(clknet_leaf_101_wb_clk_i),
    .D(\u_cpu.REG_FILE._00459_ ),
    .Q(\u_cpu.REG_FILE.rf[13][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11904_  (.CLK(clknet_leaf_95_wb_clk_i),
    .D(\u_cpu.REG_FILE._00460_ ),
    .Q(\u_cpu.REG_FILE.rf[13][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11905_  (.CLK(clknet_leaf_94_wb_clk_i),
    .D(\u_cpu.REG_FILE._00461_ ),
    .Q(\u_cpu.REG_FILE.rf[13][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11906_  (.CLK(clknet_leaf_91_wb_clk_i),
    .D(\u_cpu.REG_FILE._00462_ ),
    .Q(\u_cpu.REG_FILE.rf[13][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11907_  (.CLK(clknet_leaf_101_wb_clk_i),
    .D(\u_cpu.REG_FILE._00463_ ),
    .Q(\u_cpu.REG_FILE.rf[13][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11908_  (.CLK(clknet_leaf_107_wb_clk_i),
    .D(\u_cpu.REG_FILE._00464_ ),
    .Q(\u_cpu.REG_FILE.rf[13][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11909_  (.CLK(clknet_leaf_105_wb_clk_i),
    .D(\u_cpu.REG_FILE._00465_ ),
    .Q(\u_cpu.REG_FILE.rf[13][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11910_  (.CLK(clknet_leaf_90_wb_clk_i),
    .D(\u_cpu.REG_FILE._00466_ ),
    .Q(\u_cpu.REG_FILE.rf[13][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11911_  (.CLK(clknet_leaf_106_wb_clk_i),
    .D(\u_cpu.REG_FILE._00467_ ),
    .Q(\u_cpu.REG_FILE.rf[13][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11912_  (.CLK(clknet_leaf_78_wb_clk_i),
    .D(\u_cpu.REG_FILE._00468_ ),
    .Q(\u_cpu.REG_FILE.rf[13][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11913_  (.CLK(clknet_leaf_105_wb_clk_i),
    .D(\u_cpu.REG_FILE._00469_ ),
    .Q(\u_cpu.REG_FILE.rf[13][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11914_  (.CLK(clknet_leaf_82_wb_clk_i),
    .D(\u_cpu.REG_FILE._00470_ ),
    .Q(\u_cpu.REG_FILE.rf[13][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11915_  (.CLK(clknet_leaf_79_wb_clk_i),
    .D(\u_cpu.REG_FILE._00471_ ),
    .Q(\u_cpu.REG_FILE.rf[13][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11916_  (.CLK(clknet_leaf_105_wb_clk_i),
    .D(\u_cpu.REG_FILE._00472_ ),
    .Q(\u_cpu.REG_FILE.rf[13][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11917_  (.CLK(clknet_leaf_84_wb_clk_i),
    .D(\u_cpu.REG_FILE._00473_ ),
    .Q(\u_cpu.REG_FILE.rf[13][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11918_  (.CLK(clknet_leaf_85_wb_clk_i),
    .D(\u_cpu.REG_FILE._00474_ ),
    .Q(\u_cpu.REG_FILE.rf[13][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11919_  (.CLK(clknet_leaf_85_wb_clk_i),
    .D(\u_cpu.REG_FILE._00475_ ),
    .Q(\u_cpu.REG_FILE.rf[13][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11920_  (.CLK(clknet_leaf_86_wb_clk_i),
    .D(\u_cpu.REG_FILE._00476_ ),
    .Q(\u_cpu.REG_FILE.rf[13][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11921_  (.CLK(clknet_leaf_86_wb_clk_i),
    .D(\u_cpu.REG_FILE._00477_ ),
    .Q(\u_cpu.REG_FILE.rf[13][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11922_  (.CLK(clknet_leaf_110_wb_clk_i),
    .D(\u_cpu.REG_FILE._00478_ ),
    .Q(\u_cpu.REG_FILE.rf[13][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11923_  (.CLK(clknet_leaf_80_wb_clk_i),
    .D(\u_cpu.REG_FILE._00479_ ),
    .Q(\u_cpu.REG_FILE.rf[13][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11924_  (.CLK(clknet_leaf_125_wb_clk_i),
    .D(\u_cpu.REG_FILE._00480_ ),
    .Q(\u_cpu.REG_FILE.rf[14][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11925_  (.CLK(clknet_leaf_125_wb_clk_i),
    .D(\u_cpu.REG_FILE._00481_ ),
    .Q(\u_cpu.REG_FILE.rf[14][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11926_  (.CLK(clknet_leaf_124_wb_clk_i),
    .D(\u_cpu.REG_FILE._00482_ ),
    .Q(\u_cpu.REG_FILE.rf[14][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11927_  (.CLK(clknet_leaf_121_wb_clk_i),
    .D(\u_cpu.REG_FILE._00483_ ),
    .Q(\u_cpu.REG_FILE.rf[14][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11928_  (.CLK(clknet_leaf_122_wb_clk_i),
    .D(\u_cpu.REG_FILE._00484_ ),
    .Q(\u_cpu.REG_FILE.rf[14][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11929_  (.CLK(clknet_leaf_100_wb_clk_i),
    .D(\u_cpu.REG_FILE._00485_ ),
    .Q(\u_cpu.REG_FILE.rf[14][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11930_  (.CLK(clknet_leaf_101_wb_clk_i),
    .D(\u_cpu.REG_FILE._00486_ ),
    .Q(\u_cpu.REG_FILE.rf[14][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11931_  (.CLK(clknet_leaf_108_wb_clk_i),
    .D(\u_cpu.REG_FILE._00487_ ),
    .Q(\u_cpu.REG_FILE.rf[14][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11932_  (.CLK(clknet_leaf_97_wb_clk_i),
    .D(\u_cpu.REG_FILE._00488_ ),
    .Q(\u_cpu.REG_FILE.rf[14][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11933_  (.CLK(clknet_leaf_115_wb_clk_i),
    .D(\u_cpu.REG_FILE._00489_ ),
    .Q(\u_cpu.REG_FILE.rf[14][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11934_  (.CLK(clknet_leaf_97_wb_clk_i),
    .D(\u_cpu.REG_FILE._00490_ ),
    .Q(\u_cpu.REG_FILE.rf[14][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11935_  (.CLK(clknet_leaf_101_wb_clk_i),
    .D(\u_cpu.REG_FILE._00491_ ),
    .Q(\u_cpu.REG_FILE.rf[14][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11936_  (.CLK(clknet_leaf_95_wb_clk_i),
    .D(\u_cpu.REG_FILE._00492_ ),
    .Q(\u_cpu.REG_FILE.rf[14][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11937_  (.CLK(clknet_leaf_94_wb_clk_i),
    .D(\u_cpu.REG_FILE._00493_ ),
    .Q(\u_cpu.REG_FILE.rf[14][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11938_  (.CLK(clknet_leaf_91_wb_clk_i),
    .D(\u_cpu.REG_FILE._00494_ ),
    .Q(\u_cpu.REG_FILE.rf[14][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11939_  (.CLK(clknet_leaf_102_wb_clk_i),
    .D(\u_cpu.REG_FILE._00495_ ),
    .Q(\u_cpu.REG_FILE.rf[14][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11940_  (.CLK(clknet_leaf_107_wb_clk_i),
    .D(\u_cpu.REG_FILE._00496_ ),
    .Q(\u_cpu.REG_FILE.rf[14][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11941_  (.CLK(clknet_leaf_104_wb_clk_i),
    .D(\u_cpu.REG_FILE._00497_ ),
    .Q(\u_cpu.REG_FILE.rf[14][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11942_  (.CLK(clknet_leaf_90_wb_clk_i),
    .D(\u_cpu.REG_FILE._00498_ ),
    .Q(\u_cpu.REG_FILE.rf[14][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11943_  (.CLK(clknet_leaf_106_wb_clk_i),
    .D(\u_cpu.REG_FILE._00499_ ),
    .Q(\u_cpu.REG_FILE.rf[14][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11944_  (.CLK(clknet_leaf_79_wb_clk_i),
    .D(\u_cpu.REG_FILE._00500_ ),
    .Q(\u_cpu.REG_FILE.rf[14][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11945_  (.CLK(clknet_leaf_82_wb_clk_i),
    .D(\u_cpu.REG_FILE._00501_ ),
    .Q(\u_cpu.REG_FILE.rf[14][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11946_  (.CLK(clknet_leaf_81_wb_clk_i),
    .D(\u_cpu.REG_FILE._00502_ ),
    .Q(\u_cpu.REG_FILE.rf[14][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11947_  (.CLK(clknet_leaf_79_wb_clk_i),
    .D(\u_cpu.REG_FILE._00503_ ),
    .Q(\u_cpu.REG_FILE.rf[14][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11948_  (.CLK(clknet_leaf_83_wb_clk_i),
    .D(\u_cpu.REG_FILE._00504_ ),
    .Q(\u_cpu.REG_FILE.rf[14][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11949_  (.CLK(clknet_leaf_84_wb_clk_i),
    .D(\u_cpu.REG_FILE._00505_ ),
    .Q(\u_cpu.REG_FILE.rf[14][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11950_  (.CLK(clknet_leaf_85_wb_clk_i),
    .D(\u_cpu.REG_FILE._00506_ ),
    .Q(\u_cpu.REG_FILE.rf[14][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11951_  (.CLK(clknet_leaf_86_wb_clk_i),
    .D(\u_cpu.REG_FILE._00507_ ),
    .Q(\u_cpu.REG_FILE.rf[14][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11952_  (.CLK(clknet_leaf_85_wb_clk_i),
    .D(\u_cpu.REG_FILE._00508_ ),
    .Q(\u_cpu.REG_FILE.rf[14][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11953_  (.CLK(clknet_leaf_86_wb_clk_i),
    .D(\u_cpu.REG_FILE._00509_ ),
    .Q(\u_cpu.REG_FILE.rf[14][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11954_  (.CLK(clknet_leaf_109_wb_clk_i),
    .D(\u_cpu.REG_FILE._00510_ ),
    .Q(\u_cpu.REG_FILE.rf[14][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11955_  (.CLK(clknet_leaf_80_wb_clk_i),
    .D(\u_cpu.REG_FILE._00511_ ),
    .Q(\u_cpu.REG_FILE.rf[14][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11956_  (.CLK(clknet_leaf_125_wb_clk_i),
    .D(\u_cpu.REG_FILE._00512_ ),
    .Q(\u_cpu.REG_FILE.rf[15][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11957_  (.CLK(clknet_leaf_126_wb_clk_i),
    .D(\u_cpu.REG_FILE._00513_ ),
    .Q(\u_cpu.REG_FILE.rf[15][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11958_  (.CLK(clknet_leaf_123_wb_clk_i),
    .D(\u_cpu.REG_FILE._00514_ ),
    .Q(\u_cpu.REG_FILE.rf[15][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11959_  (.CLK(clknet_leaf_121_wb_clk_i),
    .D(\u_cpu.REG_FILE._00515_ ),
    .Q(\u_cpu.REG_FILE.rf[15][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11960_  (.CLK(clknet_leaf_122_wb_clk_i),
    .D(\u_cpu.REG_FILE._00516_ ),
    .Q(\u_cpu.REG_FILE.rf[15][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11961_  (.CLK(clknet_leaf_101_wb_clk_i),
    .D(\u_cpu.REG_FILE._00517_ ),
    .Q(\u_cpu.REG_FILE.rf[15][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11962_  (.CLK(clknet_leaf_101_wb_clk_i),
    .D(\u_cpu.REG_FILE._00518_ ),
    .Q(\u_cpu.REG_FILE.rf[15][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11963_  (.CLK(clknet_leaf_108_wb_clk_i),
    .D(\u_cpu.REG_FILE._00519_ ),
    .Q(\u_cpu.REG_FILE.rf[15][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11964_  (.CLK(clknet_leaf_97_wb_clk_i),
    .D(\u_cpu.REG_FILE._00520_ ),
    .Q(\u_cpu.REG_FILE.rf[15][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11965_  (.CLK(clknet_leaf_115_wb_clk_i),
    .D(\u_cpu.REG_FILE._00521_ ),
    .Q(\u_cpu.REG_FILE.rf[15][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11966_  (.CLK(clknet_leaf_97_wb_clk_i),
    .D(\u_cpu.REG_FILE._00522_ ),
    .Q(\u_cpu.REG_FILE.rf[15][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11967_  (.CLK(clknet_leaf_101_wb_clk_i),
    .D(\u_cpu.REG_FILE._00523_ ),
    .Q(\u_cpu.REG_FILE.rf[15][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11968_  (.CLK(clknet_leaf_95_wb_clk_i),
    .D(\u_cpu.REG_FILE._00524_ ),
    .Q(\u_cpu.REG_FILE.rf[15][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11969_  (.CLK(clknet_leaf_95_wb_clk_i),
    .D(\u_cpu.REG_FILE._00525_ ),
    .Q(\u_cpu.REG_FILE.rf[15][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11970_  (.CLK(clknet_leaf_91_wb_clk_i),
    .D(\u_cpu.REG_FILE._00526_ ),
    .Q(\u_cpu.REG_FILE.rf[15][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11971_  (.CLK(clknet_leaf_102_wb_clk_i),
    .D(\u_cpu.REG_FILE._00527_ ),
    .Q(\u_cpu.REG_FILE.rf[15][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11972_  (.CLK(clknet_leaf_107_wb_clk_i),
    .D(\u_cpu.REG_FILE._00528_ ),
    .Q(\u_cpu.REG_FILE.rf[15][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11973_  (.CLK(clknet_leaf_105_wb_clk_i),
    .D(\u_cpu.REG_FILE._00529_ ),
    .Q(\u_cpu.REG_FILE.rf[15][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11974_  (.CLK(clknet_leaf_83_wb_clk_i),
    .D(\u_cpu.REG_FILE._00530_ ),
    .Q(\u_cpu.REG_FILE.rf[15][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11975_  (.CLK(clknet_leaf_106_wb_clk_i),
    .D(\u_cpu.REG_FILE._00531_ ),
    .Q(\u_cpu.REG_FILE.rf[15][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11976_  (.CLK(clknet_leaf_78_wb_clk_i),
    .D(\u_cpu.REG_FILE._00532_ ),
    .Q(\u_cpu.REG_FILE.rf[15][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11977_  (.CLK(clknet_leaf_106_wb_clk_i),
    .D(\u_cpu.REG_FILE._00533_ ),
    .Q(\u_cpu.REG_FILE.rf[15][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11978_  (.CLK(clknet_leaf_82_wb_clk_i),
    .D(\u_cpu.REG_FILE._00534_ ),
    .Q(\u_cpu.REG_FILE.rf[15][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11979_  (.CLK(clknet_leaf_79_wb_clk_i),
    .D(\u_cpu.REG_FILE._00535_ ),
    .Q(\u_cpu.REG_FILE.rf[15][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11980_  (.CLK(clknet_leaf_90_wb_clk_i),
    .D(\u_cpu.REG_FILE._00536_ ),
    .Q(\u_cpu.REG_FILE.rf[15][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11981_  (.CLK(clknet_leaf_84_wb_clk_i),
    .D(\u_cpu.REG_FILE._00537_ ),
    .Q(\u_cpu.REG_FILE.rf[15][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11982_  (.CLK(clknet_leaf_85_wb_clk_i),
    .D(\u_cpu.REG_FILE._00538_ ),
    .Q(\u_cpu.REG_FILE.rf[15][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11983_  (.CLK(clknet_leaf_85_wb_clk_i),
    .D(\u_cpu.REG_FILE._00539_ ),
    .Q(\u_cpu.REG_FILE.rf[15][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11984_  (.CLK(clknet_leaf_86_wb_clk_i),
    .D(\u_cpu.REG_FILE._00540_ ),
    .Q(\u_cpu.REG_FILE.rf[15][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11985_  (.CLK(clknet_leaf_86_wb_clk_i),
    .D(\u_cpu.REG_FILE._00541_ ),
    .Q(\u_cpu.REG_FILE.rf[15][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11986_  (.CLK(clknet_leaf_109_wb_clk_i),
    .D(\u_cpu.REG_FILE._00542_ ),
    .Q(\u_cpu.REG_FILE.rf[15][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11987_  (.CLK(clknet_leaf_80_wb_clk_i),
    .D(\u_cpu.REG_FILE._00543_ ),
    .Q(\u_cpu.REG_FILE.rf[15][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11988_  (.CLK(clknet_leaf_128_wb_clk_i),
    .D(\u_cpu.REG_FILE._00544_ ),
    .Q(\u_cpu.REG_FILE.rf[16][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11989_  (.CLK(clknet_leaf_129_wb_clk_i),
    .D(\u_cpu.REG_FILE._00545_ ),
    .Q(\u_cpu.REG_FILE.rf[16][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11990_  (.CLK(clknet_leaf_128_wb_clk_i),
    .D(\u_cpu.REG_FILE._00546_ ),
    .Q(\u_cpu.REG_FILE.rf[16][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11991_  (.CLK(clknet_leaf_117_wb_clk_i),
    .D(\u_cpu.REG_FILE._00547_ ),
    .Q(\u_cpu.REG_FILE.rf[16][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11992_  (.CLK(clknet_leaf_119_wb_clk_i),
    .D(\u_cpu.REG_FILE._00548_ ),
    .Q(\u_cpu.REG_FILE.rf[16][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11993_  (.CLK(clknet_leaf_128_wb_clk_i),
    .D(\u_cpu.REG_FILE._00549_ ),
    .Q(\u_cpu.REG_FILE.rf[16][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11994_  (.CLK(clknet_leaf_129_wb_clk_i),
    .D(\u_cpu.REG_FILE._00550_ ),
    .Q(\u_cpu.REG_FILE.rf[16][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11995_  (.CLK(clknet_leaf_118_wb_clk_i),
    .D(\u_cpu.REG_FILE._00551_ ),
    .Q(\u_cpu.REG_FILE.rf[16][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11996_  (.CLK(clknet_leaf_128_wb_clk_i),
    .D(\u_cpu.REG_FILE._00552_ ),
    .Q(\u_cpu.REG_FILE.rf[16][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11997_  (.CLK(clknet_leaf_5_wb_clk_i),
    .D(\u_cpu.REG_FILE._00553_ ),
    .Q(\u_cpu.REG_FILE.rf[16][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11998_  (.CLK(clknet_leaf_128_wb_clk_i),
    .D(\u_cpu.REG_FILE._00554_ ),
    .Q(\u_cpu.REG_FILE.rf[16][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._11999_  (.CLK(clknet_leaf_41_wb_clk_i),
    .D(\u_cpu.REG_FILE._00555_ ),
    .Q(\u_cpu.REG_FILE.rf[16][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12000_  (.CLK(clknet_leaf_119_wb_clk_i),
    .D(\u_cpu.REG_FILE._00556_ ),
    .Q(\u_cpu.REG_FILE.rf[16][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12001_  (.CLK(clknet_leaf_119_wb_clk_i),
    .D(\u_cpu.REG_FILE._00557_ ),
    .Q(\u_cpu.REG_FILE.rf[16][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12002_  (.CLK(clknet_leaf_119_wb_clk_i),
    .D(\u_cpu.REG_FILE._00558_ ),
    .Q(\u_cpu.REG_FILE.rf[16][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12003_  (.CLK(clknet_leaf_37_wb_clk_i),
    .D(\u_cpu.REG_FILE._00559_ ),
    .Q(\u_cpu.REG_FILE.rf[16][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12004_  (.CLK(clknet_leaf_41_wb_clk_i),
    .D(\u_cpu.REG_FILE._00560_ ),
    .Q(\u_cpu.REG_FILE.rf[16][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12005_  (.CLK(clknet_leaf_36_wb_clk_i),
    .D(\u_cpu.REG_FILE._00561_ ),
    .Q(\u_cpu.REG_FILE.rf[16][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12006_  (.CLK(clknet_leaf_35_wb_clk_i),
    .D(\u_cpu.REG_FILE._00562_ ),
    .Q(\u_cpu.REG_FILE.rf[16][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12007_  (.CLK(clknet_leaf_41_wb_clk_i),
    .D(\u_cpu.REG_FILE._00563_ ),
    .Q(\u_cpu.REG_FILE.rf[16][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12008_  (.CLK(clknet_leaf_44_wb_clk_i),
    .D(\u_cpu.REG_FILE._00564_ ),
    .Q(\u_cpu.REG_FILE.rf[16][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12009_  (.CLK(clknet_leaf_49_wb_clk_i),
    .D(\u_cpu.REG_FILE._00565_ ),
    .Q(\u_cpu.REG_FILE.rf[16][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12010_  (.CLK(clknet_leaf_77_wb_clk_i),
    .D(\u_cpu.REG_FILE._00566_ ),
    .Q(\u_cpu.REG_FILE.rf[16][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12011_  (.CLK(clknet_leaf_47_wb_clk_i),
    .D(\u_cpu.REG_FILE._00567_ ),
    .Q(\u_cpu.REG_FILE.rf[16][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12012_  (.CLK(clknet_leaf_50_wb_clk_i),
    .D(\u_cpu.REG_FILE._00568_ ),
    .Q(\u_cpu.REG_FILE.rf[16][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12013_  (.CLK(clknet_leaf_77_wb_clk_i),
    .D(\u_cpu.REG_FILE._00569_ ),
    .Q(\u_cpu.REG_FILE.rf[16][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12014_  (.CLK(clknet_leaf_49_wb_clk_i),
    .D(\u_cpu.REG_FILE._00570_ ),
    .Q(\u_cpu.REG_FILE.rf[16][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12015_  (.CLK(clknet_leaf_49_wb_clk_i),
    .D(\u_cpu.REG_FILE._00571_ ),
    .Q(\u_cpu.REG_FILE.rf[16][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12016_  (.CLK(clknet_leaf_59_wb_clk_i),
    .D(\u_cpu.REG_FILE._00572_ ),
    .Q(\u_cpu.REG_FILE.rf[16][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12017_  (.CLK(clknet_leaf_77_wb_clk_i),
    .D(\u_cpu.REG_FILE._00573_ ),
    .Q(\u_cpu.REG_FILE.rf[16][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12018_  (.CLK(clknet_leaf_9_wb_clk_i),
    .D(\u_cpu.REG_FILE._00574_ ),
    .Q(\u_cpu.REG_FILE.rf[16][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12019_  (.CLK(clknet_leaf_112_wb_clk_i),
    .D(\u_cpu.REG_FILE._00575_ ),
    .Q(\u_cpu.REG_FILE.rf[16][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12020_  (.CLK(clknet_leaf_2_wb_clk_i),
    .D(\u_cpu.REG_FILE._00576_ ),
    .Q(\u_cpu.REG_FILE.rf[17][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12021_  (.CLK(clknet_leaf_2_wb_clk_i),
    .D(\u_cpu.REG_FILE._00577_ ),
    .Q(\u_cpu.REG_FILE.rf[17][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12022_  (.CLK(clknet_leaf_7_wb_clk_i),
    .D(\u_cpu.REG_FILE._00578_ ),
    .Q(\u_cpu.REG_FILE.rf[17][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12023_  (.CLK(clknet_leaf_10_wb_clk_i),
    .D(\u_cpu.REG_FILE._00579_ ),
    .Q(\u_cpu.REG_FILE.rf[17][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12024_  (.CLK(clknet_leaf_5_wb_clk_i),
    .D(\u_cpu.REG_FILE._00580_ ),
    .Q(\u_cpu.REG_FILE.rf[17][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12025_  (.CLK(clknet_leaf_5_wb_clk_i),
    .D(\u_cpu.REG_FILE._00581_ ),
    .Q(\u_cpu.REG_FILE.rf[17][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12026_  (.CLK(clknet_leaf_129_wb_clk_i),
    .D(\u_cpu.REG_FILE._00582_ ),
    .Q(\u_cpu.REG_FILE.rf[17][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12027_  (.CLK(clknet_leaf_117_wb_clk_i),
    .D(\u_cpu.REG_FILE._00583_ ),
    .Q(\u_cpu.REG_FILE.rf[17][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12028_  (.CLK(clknet_leaf_129_wb_clk_i),
    .D(\u_cpu.REG_FILE._00584_ ),
    .Q(\u_cpu.REG_FILE.rf[17][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12029_  (.CLK(clknet_leaf_7_wb_clk_i),
    .D(\u_cpu.REG_FILE._00585_ ),
    .Q(\u_cpu.REG_FILE.rf[17][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12030_  (.CLK(clknet_leaf_128_wb_clk_i),
    .D(\u_cpu.REG_FILE._00586_ ),
    .Q(\u_cpu.REG_FILE.rf[17][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12031_  (.CLK(clknet_leaf_38_wb_clk_i),
    .D(\u_cpu.REG_FILE._00587_ ),
    .Q(\u_cpu.REG_FILE.rf[17][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12032_  (.CLK(clknet_leaf_119_wb_clk_i),
    .D(\u_cpu.REG_FILE._00588_ ),
    .Q(\u_cpu.REG_FILE.rf[17][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12033_  (.CLK(clknet_leaf_128_wb_clk_i),
    .D(\u_cpu.REG_FILE._00589_ ),
    .Q(\u_cpu.REG_FILE.rf[17][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12034_  (.CLK(clknet_leaf_119_wb_clk_i),
    .D(\u_cpu.REG_FILE._00590_ ),
    .Q(\u_cpu.REG_FILE.rf[17][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12035_  (.CLK(clknet_leaf_36_wb_clk_i),
    .D(\u_cpu.REG_FILE._00591_ ),
    .Q(\u_cpu.REG_FILE.rf[17][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12036_  (.CLK(clknet_leaf_39_wb_clk_i),
    .D(\u_cpu.REG_FILE._00592_ ),
    .Q(\u_cpu.REG_FILE.rf[17][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12037_  (.CLK(clknet_leaf_36_wb_clk_i),
    .D(\u_cpu.REG_FILE._00593_ ),
    .Q(\u_cpu.REG_FILE.rf[17][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12038_  (.CLK(clknet_leaf_35_wb_clk_i),
    .D(\u_cpu.REG_FILE._00594_ ),
    .Q(\u_cpu.REG_FILE.rf[17][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12039_  (.CLK(clknet_leaf_41_wb_clk_i),
    .D(\u_cpu.REG_FILE._00595_ ),
    .Q(\u_cpu.REG_FILE.rf[17][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12040_  (.CLK(clknet_leaf_47_wb_clk_i),
    .D(\u_cpu.REG_FILE._00596_ ),
    .Q(\u_cpu.REG_FILE.rf[17][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12041_  (.CLK(clknet_leaf_46_wb_clk_i),
    .D(\u_cpu.REG_FILE._00597_ ),
    .Q(\u_cpu.REG_FILE.rf[17][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12042_  (.CLK(clknet_leaf_77_wb_clk_i),
    .D(\u_cpu.REG_FILE._00598_ ),
    .Q(\u_cpu.REG_FILE.rf[17][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12043_  (.CLK(clknet_leaf_46_wb_clk_i),
    .D(\u_cpu.REG_FILE._00599_ ),
    .Q(\u_cpu.REG_FILE.rf[17][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12044_  (.CLK(clknet_leaf_51_wb_clk_i),
    .D(\u_cpu.REG_FILE._00600_ ),
    .Q(\u_cpu.REG_FILE.rf[17][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12045_  (.CLK(clknet_leaf_42_wb_clk_i),
    .D(\u_cpu.REG_FILE._00601_ ),
    .Q(\u_cpu.REG_FILE.rf[17][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12046_  (.CLK(clknet_leaf_51_wb_clk_i),
    .D(\u_cpu.REG_FILE._00602_ ),
    .Q(\u_cpu.REG_FILE.rf[17][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12047_  (.CLK(clknet_leaf_46_wb_clk_i),
    .D(\u_cpu.REG_FILE._00603_ ),
    .Q(\u_cpu.REG_FILE.rf[17][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12048_  (.CLK(clknet_leaf_51_wb_clk_i),
    .D(\u_cpu.REG_FILE._00604_ ),
    .Q(\u_cpu.REG_FILE.rf[17][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12049_  (.CLK(clknet_leaf_77_wb_clk_i),
    .D(\u_cpu.REG_FILE._00605_ ),
    .Q(\u_cpu.REG_FILE.rf[17][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12050_  (.CLK(clknet_leaf_41_wb_clk_i),
    .D(\u_cpu.REG_FILE._00606_ ),
    .Q(\u_cpu.REG_FILE.rf[17][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12051_  (.CLK(clknet_leaf_9_wb_clk_i),
    .D(\u_cpu.REG_FILE._00607_ ),
    .Q(\u_cpu.REG_FILE.rf[17][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12052_  (.CLK(clknet_leaf_128_wb_clk_i),
    .D(\u_cpu.REG_FILE._00608_ ),
    .Q(\u_cpu.REG_FILE.rf[18][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12053_  (.CLK(clknet_leaf_129_wb_clk_i),
    .D(\u_cpu.REG_FILE._00609_ ),
    .Q(\u_cpu.REG_FILE.rf[18][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12054_  (.CLK(clknet_leaf_128_wb_clk_i),
    .D(\u_cpu.REG_FILE._00610_ ),
    .Q(\u_cpu.REG_FILE.rf[18][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12055_  (.CLK(clknet_leaf_114_wb_clk_i),
    .D(\u_cpu.REG_FILE._00611_ ),
    .Q(\u_cpu.REG_FILE.rf[18][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12056_  (.CLK(clknet_leaf_119_wb_clk_i),
    .D(\u_cpu.REG_FILE._00612_ ),
    .Q(\u_cpu.REG_FILE.rf[18][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12057_  (.CLK(clknet_leaf_119_wb_clk_i),
    .D(\u_cpu.REG_FILE._00613_ ),
    .Q(\u_cpu.REG_FILE.rf[18][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12058_  (.CLK(clknet_leaf_129_wb_clk_i),
    .D(\u_cpu.REG_FILE._00614_ ),
    .Q(\u_cpu.REG_FILE.rf[18][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12059_  (.CLK(clknet_leaf_118_wb_clk_i),
    .D(\u_cpu.REG_FILE._00615_ ),
    .Q(\u_cpu.REG_FILE.rf[18][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12060_  (.CLK(clknet_leaf_128_wb_clk_i),
    .D(\u_cpu.REG_FILE._00616_ ),
    .Q(\u_cpu.REG_FILE.rf[18][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12061_  (.CLK(clknet_leaf_7_wb_clk_i),
    .D(\u_cpu.REG_FILE._00617_ ),
    .Q(\u_cpu.REG_FILE.rf[18][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12062_  (.CLK(clknet_leaf_119_wb_clk_i),
    .D(\u_cpu.REG_FILE._00618_ ),
    .Q(\u_cpu.REG_FILE.rf[18][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12063_  (.CLK(clknet_leaf_41_wb_clk_i),
    .D(\u_cpu.REG_FILE._00619_ ),
    .Q(\u_cpu.REG_FILE.rf[18][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12064_  (.CLK(clknet_leaf_119_wb_clk_i),
    .D(\u_cpu.REG_FILE._00620_ ),
    .Q(\u_cpu.REG_FILE.rf[18][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12065_  (.CLK(clknet_leaf_119_wb_clk_i),
    .D(\u_cpu.REG_FILE._00621_ ),
    .Q(\u_cpu.REG_FILE.rf[18][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12066_  (.CLK(clknet_leaf_119_wb_clk_i),
    .D(\u_cpu.REG_FILE._00622_ ),
    .Q(\u_cpu.REG_FILE.rf[18][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12067_  (.CLK(clknet_leaf_37_wb_clk_i),
    .D(\u_cpu.REG_FILE._00623_ ),
    .Q(\u_cpu.REG_FILE.rf[18][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12068_  (.CLK(clknet_leaf_39_wb_clk_i),
    .D(\u_cpu.REG_FILE._00624_ ),
    .Q(\u_cpu.REG_FILE.rf[18][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12069_  (.CLK(clknet_leaf_37_wb_clk_i),
    .D(\u_cpu.REG_FILE._00625_ ),
    .Q(\u_cpu.REG_FILE.rf[18][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12070_  (.CLK(clknet_leaf_35_wb_clk_i),
    .D(\u_cpu.REG_FILE._00626_ ),
    .Q(\u_cpu.REG_FILE.rf[18][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12071_  (.CLK(clknet_leaf_41_wb_clk_i),
    .D(\u_cpu.REG_FILE._00627_ ),
    .Q(\u_cpu.REG_FILE.rf[18][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12072_  (.CLK(clknet_leaf_44_wb_clk_i),
    .D(\u_cpu.REG_FILE._00628_ ),
    .Q(\u_cpu.REG_FILE.rf[18][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12073_  (.CLK(clknet_leaf_47_wb_clk_i),
    .D(\u_cpu.REG_FILE._00629_ ),
    .Q(\u_cpu.REG_FILE.rf[18][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12074_  (.CLK(clknet_leaf_77_wb_clk_i),
    .D(\u_cpu.REG_FILE._00630_ ),
    .Q(\u_cpu.REG_FILE.rf[18][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12075_  (.CLK(clknet_leaf_47_wb_clk_i),
    .D(\u_cpu.REG_FILE._00631_ ),
    .Q(\u_cpu.REG_FILE.rf[18][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12076_  (.CLK(clknet_leaf_49_wb_clk_i),
    .D(\u_cpu.REG_FILE._00632_ ),
    .Q(\u_cpu.REG_FILE.rf[18][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12077_  (.CLK(clknet_leaf_112_wb_clk_i),
    .D(\u_cpu.REG_FILE._00633_ ),
    .Q(\u_cpu.REG_FILE.rf[18][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12078_  (.CLK(clknet_leaf_49_wb_clk_i),
    .D(\u_cpu.REG_FILE._00634_ ),
    .Q(\u_cpu.REG_FILE.rf[18][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12079_  (.CLK(clknet_leaf_49_wb_clk_i),
    .D(\u_cpu.REG_FILE._00635_ ),
    .Q(\u_cpu.REG_FILE.rf[18][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12080_  (.CLK(clknet_leaf_49_wb_clk_i),
    .D(\u_cpu.REG_FILE._00636_ ),
    .Q(\u_cpu.REG_FILE.rf[18][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12081_  (.CLK(clknet_leaf_111_wb_clk_i),
    .D(\u_cpu.REG_FILE._00637_ ),
    .Q(\u_cpu.REG_FILE.rf[18][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12082_  (.CLK(clknet_leaf_10_wb_clk_i),
    .D(\u_cpu.REG_FILE._00638_ ),
    .Q(\u_cpu.REG_FILE.rf[18][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12083_  (.CLK(clknet_leaf_42_wb_clk_i),
    .D(\u_cpu.REG_FILE._00639_ ),
    .Q(\u_cpu.REG_FILE.rf[18][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12084_  (.CLK(clknet_leaf_127_wb_clk_i),
    .D(\u_cpu.REG_FILE._00640_ ),
    .Q(\u_cpu.REG_FILE.rf[1][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12085_  (.CLK(clknet_leaf_127_wb_clk_i),
    .D(\u_cpu.REG_FILE._00641_ ),
    .Q(\u_cpu.REG_FILE.rf[1][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12086_  (.CLK(clknet_leaf_120_wb_clk_i),
    .D(\u_cpu.REG_FILE._00642_ ),
    .Q(\u_cpu.REG_FILE.rf[1][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12087_  (.CLK(clknet_leaf_117_wb_clk_i),
    .D(\u_cpu.REG_FILE._00643_ ),
    .Q(\u_cpu.REG_FILE.rf[1][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12088_  (.CLK(clknet_leaf_119_wb_clk_i),
    .D(\u_cpu.REG_FILE._00644_ ),
    .Q(\u_cpu.REG_FILE.rf[1][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12089_  (.CLK(clknet_leaf_120_wb_clk_i),
    .D(\u_cpu.REG_FILE._00645_ ),
    .Q(\u_cpu.REG_FILE.rf[1][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12090_  (.CLK(clknet_leaf_127_wb_clk_i),
    .D(\u_cpu.REG_FILE._00646_ ),
    .Q(\u_cpu.REG_FILE.rf[1][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12091_  (.CLK(clknet_leaf_8_wb_clk_i),
    .D(\u_cpu.REG_FILE._00647_ ),
    .Q(\u_cpu.REG_FILE.rf[1][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12092_  (.CLK(clknet_leaf_127_wb_clk_i),
    .D(\u_cpu.REG_FILE._00648_ ),
    .Q(\u_cpu.REG_FILE.rf[1][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12093_  (.CLK(clknet_leaf_9_wb_clk_i),
    .D(\u_cpu.REG_FILE._00649_ ),
    .Q(\u_cpu.REG_FILE.rf[1][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12094_  (.CLK(clknet_leaf_99_wb_clk_i),
    .D(\u_cpu.REG_FILE._00650_ ),
    .Q(\u_cpu.REG_FILE.rf[1][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12095_  (.CLK(clknet_leaf_111_wb_clk_i),
    .D(\u_cpu.REG_FILE._00651_ ),
    .Q(\u_cpu.REG_FILE.rf[1][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12096_  (.CLK(clknet_leaf_93_wb_clk_i),
    .D(\u_cpu.REG_FILE._00652_ ),
    .Q(\u_cpu.REG_FILE.rf[1][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12097_  (.CLK(clknet_leaf_92_wb_clk_i),
    .D(\u_cpu.REG_FILE._00653_ ),
    .Q(\u_cpu.REG_FILE.rf[1][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12098_  (.CLK(clknet_leaf_91_wb_clk_i),
    .D(\u_cpu.REG_FILE._00654_ ),
    .Q(\u_cpu.REG_FILE.rf[1][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12099_  (.CLK(clknet_leaf_100_wb_clk_i),
    .D(\u_cpu.REG_FILE._00655_ ),
    .Q(\u_cpu.REG_FILE.rf[1][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12100_  (.CLK(clknet_leaf_110_wb_clk_i),
    .D(\u_cpu.REG_FILE._00656_ ),
    .Q(\u_cpu.REG_FILE.rf[1][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12101_  (.CLK(clknet_leaf_105_wb_clk_i),
    .D(\u_cpu.REG_FILE._00657_ ),
    .Q(\u_cpu.REG_FILE.rf[1][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12102_  (.CLK(clknet_leaf_49_wb_clk_i),
    .D(\u_cpu.REG_FILE._00658_ ),
    .Q(\u_cpu.REG_FILE.rf[1][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12103_  (.CLK(clknet_leaf_44_wb_clk_i),
    .D(\u_cpu.REG_FILE._00659_ ),
    .Q(\u_cpu.REG_FILE.rf[1][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12104_  (.CLK(clknet_leaf_49_wb_clk_i),
    .D(\u_cpu.REG_FILE._00660_ ),
    .Q(\u_cpu.REG_FILE.rf[1][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12105_  (.CLK(clknet_leaf_47_wb_clk_i),
    .D(\u_cpu.REG_FILE._00661_ ),
    .Q(\u_cpu.REG_FILE.rf[1][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12106_  (.CLK(clknet_leaf_49_wb_clk_i),
    .D(\u_cpu.REG_FILE._00662_ ),
    .Q(\u_cpu.REG_FILE.rf[1][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12107_  (.CLK(clknet_leaf_72_wb_clk_i),
    .D(\u_cpu.REG_FILE._00663_ ),
    .Q(\u_cpu.REG_FILE.rf[1][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12108_  (.CLK(clknet_leaf_59_wb_clk_i),
    .D(\u_cpu.REG_FILE._00664_ ),
    .Q(\u_cpu.REG_FILE.rf[1][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12109_  (.CLK(clknet_leaf_71_wb_clk_i),
    .D(\u_cpu.REG_FILE._00665_ ),
    .Q(\u_cpu.REG_FILE.rf[1][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12110_  (.CLK(clknet_leaf_60_wb_clk_i),
    .D(\u_cpu.REG_FILE._00666_ ),
    .Q(\u_cpu.REG_FILE.rf[1][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12111_  (.CLK(clknet_leaf_59_wb_clk_i),
    .D(\u_cpu.REG_FILE._00667_ ),
    .Q(\u_cpu.REG_FILE.rf[1][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12112_  (.CLK(clknet_leaf_59_wb_clk_i),
    .D(\u_cpu.REG_FILE._00668_ ),
    .Q(\u_cpu.REG_FILE.rf[1][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12113_  (.CLK(clknet_leaf_60_wb_clk_i),
    .D(\u_cpu.REG_FILE._00669_ ),
    .Q(\u_cpu.REG_FILE.rf[1][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12114_  (.CLK(clknet_leaf_9_wb_clk_i),
    .D(\u_cpu.REG_FILE._00670_ ),
    .Q(\u_cpu.REG_FILE.rf[1][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12115_  (.CLK(clknet_leaf_74_wb_clk_i),
    .D(\u_cpu.REG_FILE._00671_ ),
    .Q(\u_cpu.REG_FILE.rf[1][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12116_  (.CLK(clknet_leaf_0_wb_clk_i),
    .D(\u_cpu.REG_FILE._00672_ ),
    .Q(\u_cpu.REG_FILE.rf[20][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12117_  (.CLK(clknet_leaf_0_wb_clk_i),
    .D(\u_cpu.REG_FILE._00673_ ),
    .Q(\u_cpu.REG_FILE.rf[20][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12118_  (.CLK(clknet_leaf_12_wb_clk_i),
    .D(\u_cpu.REG_FILE._00674_ ),
    .Q(\u_cpu.REG_FILE.rf[20][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12119_  (.CLK(clknet_leaf_11_wb_clk_i),
    .D(\u_cpu.REG_FILE._00675_ ),
    .Q(\u_cpu.REG_FILE.rf[20][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12120_  (.CLK(clknet_leaf_12_wb_clk_i),
    .D(\u_cpu.REG_FILE._00676_ ),
    .Q(\u_cpu.REG_FILE.rf[20][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12121_  (.CLK(clknet_leaf_18_wb_clk_i),
    .D(\u_cpu.REG_FILE._00677_ ),
    .Q(\u_cpu.REG_FILE.rf[20][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12122_  (.CLK(clknet_leaf_0_wb_clk_i),
    .D(\u_cpu.REG_FILE._00678_ ),
    .Q(\u_cpu.REG_FILE.rf[20][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12123_  (.CLK(clknet_leaf_7_wb_clk_i),
    .D(\u_cpu.REG_FILE._00679_ ),
    .Q(\u_cpu.REG_FILE.rf[20][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12124_  (.CLK(clknet_leaf_18_wb_clk_i),
    .D(\u_cpu.REG_FILE._00680_ ),
    .Q(\u_cpu.REG_FILE.rf[20][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12125_  (.CLK(clknet_leaf_13_wb_clk_i),
    .D(\u_cpu.REG_FILE._00681_ ),
    .Q(\u_cpu.REG_FILE.rf[20][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12126_  (.CLK(clknet_leaf_16_wb_clk_i),
    .D(\u_cpu.REG_FILE._00682_ ),
    .Q(\u_cpu.REG_FILE.rf[20][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12127_  (.CLK(clknet_leaf_38_wb_clk_i),
    .D(\u_cpu.REG_FILE._00683_ ),
    .Q(\u_cpu.REG_FILE.rf[20][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12128_  (.CLK(clknet_leaf_29_wb_clk_i),
    .D(\u_cpu.REG_FILE._00684_ ),
    .Q(\u_cpu.REG_FILE.rf[20][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12129_  (.CLK(clknet_leaf_28_wb_clk_i),
    .D(\u_cpu.REG_FILE._00685_ ),
    .Q(\u_cpu.REG_FILE.rf[20][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12130_  (.CLK(clknet_leaf_15_wb_clk_i),
    .D(\u_cpu.REG_FILE._00686_ ),
    .Q(\u_cpu.REG_FILE.rf[20][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12131_  (.CLK(clknet_leaf_29_wb_clk_i),
    .D(\u_cpu.REG_FILE._00687_ ),
    .Q(\u_cpu.REG_FILE.rf[20][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12132_  (.CLK(clknet_leaf_39_wb_clk_i),
    .D(\u_cpu.REG_FILE._00688_ ),
    .Q(\u_cpu.REG_FILE.rf[20][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12133_  (.CLK(clknet_leaf_29_wb_clk_i),
    .D(\u_cpu.REG_FILE._00689_ ),
    .Q(\u_cpu.REG_FILE.rf[20][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12134_  (.CLK(clknet_leaf_30_wb_clk_i),
    .D(\u_cpu.REG_FILE._00690_ ),
    .Q(\u_cpu.REG_FILE.rf[20][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12135_  (.CLK(clknet_leaf_41_wb_clk_i),
    .D(\u_cpu.REG_FILE._00691_ ),
    .Q(\u_cpu.REG_FILE.rf[20][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12136_  (.CLK(clknet_leaf_57_wb_clk_i),
    .D(\u_cpu.REG_FILE._00692_ ),
    .Q(\u_cpu.REG_FILE.rf[20][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12137_  (.CLK(clknet_leaf_56_wb_clk_i),
    .D(\u_cpu.REG_FILE._00693_ ),
    .Q(\u_cpu.REG_FILE.rf[20][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12138_  (.CLK(clknet_leaf_55_wb_clk_i),
    .D(\u_cpu.REG_FILE._00694_ ),
    .Q(\u_cpu.REG_FILE.rf[20][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12139_  (.CLK(clknet_leaf_57_wb_clk_i),
    .D(\u_cpu.REG_FILE._00695_ ),
    .Q(\u_cpu.REG_FILE.rf[20][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12140_  (.CLK(clknet_leaf_55_wb_clk_i),
    .D(\u_cpu.REG_FILE._00696_ ),
    .Q(\u_cpu.REG_FILE.rf[20][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12141_  (.CLK(clknet_leaf_54_wb_clk_i),
    .D(\u_cpu.REG_FILE._00697_ ),
    .Q(\u_cpu.REG_FILE.rf[20][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12142_  (.CLK(clknet_leaf_57_wb_clk_i),
    .D(\u_cpu.REG_FILE._00698_ ),
    .Q(\u_cpu.REG_FILE.rf[20][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12143_  (.CLK(clknet_leaf_55_wb_clk_i),
    .D(\u_cpu.REG_FILE._00699_ ),
    .Q(\u_cpu.REG_FILE.rf[20][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12144_  (.CLK(clknet_leaf_55_wb_clk_i),
    .D(\u_cpu.REG_FILE._00700_ ),
    .Q(\u_cpu.REG_FILE.rf[20][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12145_  (.CLK(clknet_leaf_54_wb_clk_i),
    .D(\u_cpu.REG_FILE._00701_ ),
    .Q(\u_cpu.REG_FILE.rf[20][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12146_  (.CLK(clknet_leaf_31_wb_clk_i),
    .D(\u_cpu.REG_FILE._00702_ ),
    .Q(\u_cpu.REG_FILE.rf[20][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12147_  (.CLK(clknet_leaf_31_wb_clk_i),
    .D(\u_cpu.REG_FILE._00703_ ),
    .Q(\u_cpu.REG_FILE.rf[20][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12148_  (.CLK(clknet_leaf_0_wb_clk_i),
    .D(\u_cpu.REG_FILE._00704_ ),
    .Q(\u_cpu.REG_FILE.rf[21][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12149_  (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\u_cpu.REG_FILE._00705_ ),
    .Q(\u_cpu.REG_FILE.rf[21][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12150_  (.CLK(clknet_leaf_13_wb_clk_i),
    .D(\u_cpu.REG_FILE._00706_ ),
    .Q(\u_cpu.REG_FILE.rf[21][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12151_  (.CLK(clknet_leaf_11_wb_clk_i),
    .D(\u_cpu.REG_FILE._00707_ ),
    .Q(\u_cpu.REG_FILE.rf[21][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12152_  (.CLK(clknet_leaf_12_wb_clk_i),
    .D(\u_cpu.REG_FILE._00708_ ),
    .Q(\u_cpu.REG_FILE.rf[21][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12153_  (.CLK(clknet_leaf_18_wb_clk_i),
    .D(\u_cpu.REG_FILE._00709_ ),
    .Q(\u_cpu.REG_FILE.rf[21][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12154_  (.CLK(clknet_leaf_0_wb_clk_i),
    .D(\u_cpu.REG_FILE._00710_ ),
    .Q(\u_cpu.REG_FILE.rf[21][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12155_  (.CLK(clknet_leaf_7_wb_clk_i),
    .D(\u_cpu.REG_FILE._00711_ ),
    .Q(\u_cpu.REG_FILE.rf[21][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12156_  (.CLK(clknet_leaf_18_wb_clk_i),
    .D(\u_cpu.REG_FILE._00712_ ),
    .Q(\u_cpu.REG_FILE.rf[21][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12157_  (.CLK(clknet_leaf_14_wb_clk_i),
    .D(\u_cpu.REG_FILE._00713_ ),
    .Q(\u_cpu.REG_FILE.rf[21][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12158_  (.CLK(clknet_leaf_15_wb_clk_i),
    .D(\u_cpu.REG_FILE._00714_ ),
    .Q(\u_cpu.REG_FILE.rf[21][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12159_  (.CLK(clknet_leaf_38_wb_clk_i),
    .D(\u_cpu.REG_FILE._00715_ ),
    .Q(\u_cpu.REG_FILE.rf[21][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12160_  (.CLK(clknet_leaf_28_wb_clk_i),
    .D(\u_cpu.REG_FILE._00716_ ),
    .Q(\u_cpu.REG_FILE.rf[21][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12161_  (.CLK(clknet_leaf_28_wb_clk_i),
    .D(\u_cpu.REG_FILE._00717_ ),
    .Q(\u_cpu.REG_FILE.rf[21][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12162_  (.CLK(clknet_leaf_15_wb_clk_i),
    .D(\u_cpu.REG_FILE._00718_ ),
    .Q(\u_cpu.REG_FILE.rf[21][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12163_  (.CLK(clknet_leaf_28_wb_clk_i),
    .D(\u_cpu.REG_FILE._00719_ ),
    .Q(\u_cpu.REG_FILE.rf[21][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12164_  (.CLK(clknet_leaf_40_wb_clk_i),
    .D(\u_cpu.REG_FILE._00720_ ),
    .Q(\u_cpu.REG_FILE.rf[21][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12165_  (.CLK(clknet_leaf_29_wb_clk_i),
    .D(\u_cpu.REG_FILE._00721_ ),
    .Q(\u_cpu.REG_FILE.rf[21][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12166_  (.CLK(clknet_leaf_30_wb_clk_i),
    .D(\u_cpu.REG_FILE._00722_ ),
    .Q(\u_cpu.REG_FILE.rf[21][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12167_  (.CLK(clknet_leaf_41_wb_clk_i),
    .D(\u_cpu.REG_FILE._00723_ ),
    .Q(\u_cpu.REG_FILE.rf[21][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12168_  (.CLK(clknet_leaf_57_wb_clk_i),
    .D(\u_cpu.REG_FILE._00724_ ),
    .Q(\u_cpu.REG_FILE.rf[21][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12169_  (.CLK(clknet_leaf_55_wb_clk_i),
    .D(\u_cpu.REG_FILE._00725_ ),
    .Q(\u_cpu.REG_FILE.rf[21][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12170_  (.CLK(clknet_leaf_55_wb_clk_i),
    .D(\u_cpu.REG_FILE._00726_ ),
    .Q(\u_cpu.REG_FILE.rf[21][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12171_  (.CLK(clknet_leaf_57_wb_clk_i),
    .D(\u_cpu.REG_FILE._00727_ ),
    .Q(\u_cpu.REG_FILE.rf[21][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12172_  (.CLK(clknet_leaf_55_wb_clk_i),
    .D(\u_cpu.REG_FILE._00728_ ),
    .Q(\u_cpu.REG_FILE.rf[21][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12173_  (.CLK(clknet_leaf_31_wb_clk_i),
    .D(\u_cpu.REG_FILE._00729_ ),
    .Q(\u_cpu.REG_FILE.rf[21][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12174_  (.CLK(clknet_leaf_55_wb_clk_i),
    .D(\u_cpu.REG_FILE._00730_ ),
    .Q(\u_cpu.REG_FILE.rf[21][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12175_  (.CLK(clknet_leaf_55_wb_clk_i),
    .D(\u_cpu.REG_FILE._00731_ ),
    .Q(\u_cpu.REG_FILE.rf[21][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12176_  (.CLK(clknet_leaf_55_wb_clk_i),
    .D(\u_cpu.REG_FILE._00732_ ),
    .Q(\u_cpu.REG_FILE.rf[21][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12177_  (.CLK(clknet_leaf_55_wb_clk_i),
    .D(\u_cpu.REG_FILE._00733_ ),
    .Q(\u_cpu.REG_FILE.rf[21][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12178_  (.CLK(clknet_leaf_30_wb_clk_i),
    .D(\u_cpu.REG_FILE._00734_ ),
    .Q(\u_cpu.REG_FILE.rf[21][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12179_  (.CLK(clknet_leaf_31_wb_clk_i),
    .D(\u_cpu.REG_FILE._00735_ ),
    .Q(\u_cpu.REG_FILE.rf[21][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12180_  (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\u_cpu.REG_FILE._00736_ ),
    .Q(\u_cpu.REG_FILE.rf[22][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12181_  (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\u_cpu.REG_FILE._00737_ ),
    .Q(\u_cpu.REG_FILE.rf[22][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12182_  (.CLK(clknet_leaf_13_wb_clk_i),
    .D(\u_cpu.REG_FILE._00738_ ),
    .Q(\u_cpu.REG_FILE.rf[22][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12183_  (.CLK(clknet_leaf_11_wb_clk_i),
    .D(\u_cpu.REG_FILE._00739_ ),
    .Q(\u_cpu.REG_FILE.rf[22][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12184_  (.CLK(clknet_leaf_12_wb_clk_i),
    .D(\u_cpu.REG_FILE._00740_ ),
    .Q(\u_cpu.REG_FILE.rf[22][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12185_  (.CLK(clknet_leaf_18_wb_clk_i),
    .D(\u_cpu.REG_FILE._00741_ ),
    .Q(\u_cpu.REG_FILE.rf[22][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12186_  (.CLK(clknet_leaf_0_wb_clk_i),
    .D(\u_cpu.REG_FILE._00742_ ),
    .Q(\u_cpu.REG_FILE.rf[22][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12187_  (.CLK(clknet_leaf_7_wb_clk_i),
    .D(\u_cpu.REG_FILE._00743_ ),
    .Q(\u_cpu.REG_FILE.rf[22][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12188_  (.CLK(clknet_leaf_18_wb_clk_i),
    .D(\u_cpu.REG_FILE._00744_ ),
    .Q(\u_cpu.REG_FILE.rf[22][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12189_  (.CLK(clknet_leaf_14_wb_clk_i),
    .D(\u_cpu.REG_FILE._00745_ ),
    .Q(\u_cpu.REG_FILE.rf[22][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12190_  (.CLK(clknet_leaf_16_wb_clk_i),
    .D(\u_cpu.REG_FILE._00746_ ),
    .Q(\u_cpu.REG_FILE.rf[22][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12191_  (.CLK(clknet_leaf_38_wb_clk_i),
    .D(\u_cpu.REG_FILE._00747_ ),
    .Q(\u_cpu.REG_FILE.rf[22][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12192_  (.CLK(clknet_leaf_28_wb_clk_i),
    .D(\u_cpu.REG_FILE._00748_ ),
    .Q(\u_cpu.REG_FILE.rf[22][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12193_  (.CLK(clknet_leaf_28_wb_clk_i),
    .D(\u_cpu.REG_FILE._00749_ ),
    .Q(\u_cpu.REG_FILE.rf[22][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12194_  (.CLK(clknet_leaf_38_wb_clk_i),
    .D(\u_cpu.REG_FILE._00750_ ),
    .Q(\u_cpu.REG_FILE.rf[22][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12195_  (.CLK(clknet_leaf_29_wb_clk_i),
    .D(\u_cpu.REG_FILE._00751_ ),
    .Q(\u_cpu.REG_FILE.rf[22][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12196_  (.CLK(clknet_leaf_39_wb_clk_i),
    .D(\u_cpu.REG_FILE._00752_ ),
    .Q(\u_cpu.REG_FILE.rf[22][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12197_  (.CLK(clknet_leaf_29_wb_clk_i),
    .D(\u_cpu.REG_FILE._00753_ ),
    .Q(\u_cpu.REG_FILE.rf[22][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12198_  (.CLK(clknet_leaf_30_wb_clk_i),
    .D(\u_cpu.REG_FILE._00754_ ),
    .Q(\u_cpu.REG_FILE.rf[22][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12199_  (.CLK(clknet_leaf_40_wb_clk_i),
    .D(\u_cpu.REG_FILE._00755_ ),
    .Q(\u_cpu.REG_FILE.rf[22][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12200_  (.CLK(clknet_leaf_57_wb_clk_i),
    .D(\u_cpu.REG_FILE._00756_ ),
    .Q(\u_cpu.REG_FILE.rf[22][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12201_  (.CLK(clknet_leaf_56_wb_clk_i),
    .D(\u_cpu.REG_FILE._00757_ ),
    .Q(\u_cpu.REG_FILE.rf[22][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12202_  (.CLK(clknet_leaf_54_wb_clk_i),
    .D(\u_cpu.REG_FILE._00758_ ),
    .Q(\u_cpu.REG_FILE.rf[22][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12203_  (.CLK(clknet_leaf_57_wb_clk_i),
    .D(\u_cpu.REG_FILE._00759_ ),
    .Q(\u_cpu.REG_FILE.rf[22][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12204_  (.CLK(clknet_leaf_55_wb_clk_i),
    .D(\u_cpu.REG_FILE._00760_ ),
    .Q(\u_cpu.REG_FILE.rf[22][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12205_  (.CLK(clknet_leaf_31_wb_clk_i),
    .D(\u_cpu.REG_FILE._00761_ ),
    .Q(\u_cpu.REG_FILE.rf[22][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12206_  (.CLK(clknet_leaf_56_wb_clk_i),
    .D(\u_cpu.REG_FILE._00762_ ),
    .Q(\u_cpu.REG_FILE.rf[22][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12207_  (.CLK(clknet_leaf_55_wb_clk_i),
    .D(\u_cpu.REG_FILE._00763_ ),
    .Q(\u_cpu.REG_FILE.rf[22][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12208_  (.CLK(clknet_leaf_55_wb_clk_i),
    .D(\u_cpu.REG_FILE._00764_ ),
    .Q(\u_cpu.REG_FILE.rf[22][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12209_  (.CLK(clknet_leaf_54_wb_clk_i),
    .D(\u_cpu.REG_FILE._00765_ ),
    .Q(\u_cpu.REG_FILE.rf[22][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12210_  (.CLK(clknet_leaf_30_wb_clk_i),
    .D(\u_cpu.REG_FILE._00766_ ),
    .Q(\u_cpu.REG_FILE.rf[22][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12211_  (.CLK(clknet_leaf_31_wb_clk_i),
    .D(\u_cpu.REG_FILE._00767_ ),
    .Q(\u_cpu.REG_FILE.rf[22][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12212_  (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\u_cpu.REG_FILE._00768_ ),
    .Q(\u_cpu.REG_FILE.rf[23][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12213_  (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\u_cpu.REG_FILE._00769_ ),
    .Q(\u_cpu.REG_FILE.rf[23][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12214_  (.CLK(clknet_leaf_13_wb_clk_i),
    .D(\u_cpu.REG_FILE._00770_ ),
    .Q(\u_cpu.REG_FILE.rf[23][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12215_  (.CLK(clknet_leaf_11_wb_clk_i),
    .D(\u_cpu.REG_FILE._00771_ ),
    .Q(\u_cpu.REG_FILE.rf[23][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12216_  (.CLK(clknet_leaf_12_wb_clk_i),
    .D(\u_cpu.REG_FILE._00772_ ),
    .Q(\u_cpu.REG_FILE.rf[23][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12217_  (.CLK(clknet_leaf_18_wb_clk_i),
    .D(\u_cpu.REG_FILE._00773_ ),
    .Q(\u_cpu.REG_FILE.rf[23][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12218_  (.CLK(clknet_leaf_0_wb_clk_i),
    .D(\u_cpu.REG_FILE._00774_ ),
    .Q(\u_cpu.REG_FILE.rf[23][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12219_  (.CLK(clknet_leaf_12_wb_clk_i),
    .D(\u_cpu.REG_FILE._00775_ ),
    .Q(\u_cpu.REG_FILE.rf[23][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12220_  (.CLK(clknet_leaf_18_wb_clk_i),
    .D(\u_cpu.REG_FILE._00776_ ),
    .Q(\u_cpu.REG_FILE.rf[23][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12221_  (.CLK(clknet_leaf_14_wb_clk_i),
    .D(\u_cpu.REG_FILE._00777_ ),
    .Q(\u_cpu.REG_FILE.rf[23][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12222_  (.CLK(clknet_leaf_16_wb_clk_i),
    .D(\u_cpu.REG_FILE._00778_ ),
    .Q(\u_cpu.REG_FILE.rf[23][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12223_  (.CLK(clknet_leaf_38_wb_clk_i),
    .D(\u_cpu.REG_FILE._00779_ ),
    .Q(\u_cpu.REG_FILE.rf[23][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12224_  (.CLK(clknet_leaf_29_wb_clk_i),
    .D(\u_cpu.REG_FILE._00780_ ),
    .Q(\u_cpu.REG_FILE.rf[23][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12225_  (.CLK(clknet_leaf_28_wb_clk_i),
    .D(\u_cpu.REG_FILE._00781_ ),
    .Q(\u_cpu.REG_FILE.rf[23][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12226_  (.CLK(clknet_leaf_38_wb_clk_i),
    .D(\u_cpu.REG_FILE._00782_ ),
    .Q(\u_cpu.REG_FILE.rf[23][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12227_  (.CLK(clknet_leaf_28_wb_clk_i),
    .D(\u_cpu.REG_FILE._00783_ ),
    .Q(\u_cpu.REG_FILE.rf[23][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12228_  (.CLK(clknet_leaf_39_wb_clk_i),
    .D(\u_cpu.REG_FILE._00784_ ),
    .Q(\u_cpu.REG_FILE.rf[23][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12229_  (.CLK(clknet_leaf_29_wb_clk_i),
    .D(\u_cpu.REG_FILE._00785_ ),
    .Q(\u_cpu.REG_FILE.rf[23][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12230_  (.CLK(clknet_leaf_29_wb_clk_i),
    .D(\u_cpu.REG_FILE._00786_ ),
    .Q(\u_cpu.REG_FILE.rf[23][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12231_  (.CLK(clknet_leaf_40_wb_clk_i),
    .D(\u_cpu.REG_FILE._00787_ ),
    .Q(\u_cpu.REG_FILE.rf[23][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12232_  (.CLK(clknet_leaf_57_wb_clk_i),
    .D(\u_cpu.REG_FILE._00788_ ),
    .Q(\u_cpu.REG_FILE.rf[23][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12233_  (.CLK(clknet_leaf_53_wb_clk_i),
    .D(\u_cpu.REG_FILE._00789_ ),
    .Q(\u_cpu.REG_FILE.rf[23][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12234_  (.CLK(clknet_leaf_54_wb_clk_i),
    .D(\u_cpu.REG_FILE._00790_ ),
    .Q(\u_cpu.REG_FILE.rf[23][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12235_  (.CLK(clknet_leaf_57_wb_clk_i),
    .D(\u_cpu.REG_FILE._00791_ ),
    .Q(\u_cpu.REG_FILE.rf[23][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12236_  (.CLK(clknet_leaf_55_wb_clk_i),
    .D(\u_cpu.REG_FILE._00792_ ),
    .Q(\u_cpu.REG_FILE.rf[23][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12237_  (.CLK(clknet_leaf_54_wb_clk_i),
    .D(\u_cpu.REG_FILE._00793_ ),
    .Q(\u_cpu.REG_FILE.rf[23][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12238_  (.CLK(clknet_leaf_55_wb_clk_i),
    .D(\u_cpu.REG_FILE._00794_ ),
    .Q(\u_cpu.REG_FILE.rf[23][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12239_  (.CLK(clknet_leaf_55_wb_clk_i),
    .D(\u_cpu.REG_FILE._00795_ ),
    .Q(\u_cpu.REG_FILE.rf[23][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12240_  (.CLK(clknet_leaf_55_wb_clk_i),
    .D(\u_cpu.REG_FILE._00796_ ),
    .Q(\u_cpu.REG_FILE.rf[23][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12241_  (.CLK(clknet_leaf_55_wb_clk_i),
    .D(\u_cpu.REG_FILE._00797_ ),
    .Q(\u_cpu.REG_FILE.rf[23][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12242_  (.CLK(clknet_leaf_32_wb_clk_i),
    .D(\u_cpu.REG_FILE._00798_ ),
    .Q(\u_cpu.REG_FILE.rf[23][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12243_  (.CLK(clknet_leaf_31_wb_clk_i),
    .D(\u_cpu.REG_FILE._00799_ ),
    .Q(\u_cpu.REG_FILE.rf[23][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12244_  (.CLK(clknet_leaf_13_wb_clk_i),
    .D(\u_cpu.REG_FILE._00800_ ),
    .Q(\u_cpu.REG_FILE.rf[24][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12245_  (.CLK(clknet_leaf_18_wb_clk_i),
    .D(\u_cpu.REG_FILE._00801_ ),
    .Q(\u_cpu.REG_FILE.rf[24][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12246_  (.CLK(clknet_leaf_18_wb_clk_i),
    .D(\u_cpu.REG_FILE._00802_ ),
    .Q(\u_cpu.REG_FILE.rf[24][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12247_  (.CLK(clknet_leaf_41_wb_clk_i),
    .D(\u_cpu.REG_FILE._00803_ ),
    .Q(\u_cpu.REG_FILE.rf[24][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12248_  (.CLK(clknet_leaf_14_wb_clk_i),
    .D(\u_cpu.REG_FILE._00804_ ),
    .Q(\u_cpu.REG_FILE.rf[24][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12249_  (.CLK(clknet_leaf_17_wb_clk_i),
    .D(\u_cpu.REG_FILE._00805_ ),
    .Q(\u_cpu.REG_FILE.rf[24][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12250_  (.CLK(clknet_leaf_18_wb_clk_i),
    .D(\u_cpu.REG_FILE._00806_ ),
    .Q(\u_cpu.REG_FILE.rf[24][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12251_  (.CLK(clknet_leaf_11_wb_clk_i),
    .D(\u_cpu.REG_FILE._00807_ ),
    .Q(\u_cpu.REG_FILE.rf[24][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12252_  (.CLK(clknet_leaf_13_wb_clk_i),
    .D(\u_cpu.REG_FILE._00808_ ),
    .Q(\u_cpu.REG_FILE.rf[24][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12253_  (.CLK(clknet_leaf_17_wb_clk_i),
    .D(\u_cpu.REG_FILE._00809_ ),
    .Q(\u_cpu.REG_FILE.rf[24][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12254_  (.CLK(clknet_leaf_16_wb_clk_i),
    .D(\u_cpu.REG_FILE._00810_ ),
    .Q(\u_cpu.REG_FILE.rf[24][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12255_  (.CLK(clknet_leaf_32_wb_clk_i),
    .D(\u_cpu.REG_FILE._00811_ ),
    .Q(\u_cpu.REG_FILE.rf[24][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12256_  (.CLK(clknet_leaf_37_wb_clk_i),
    .D(\u_cpu.REG_FILE._00812_ ),
    .Q(\u_cpu.REG_FILE.rf[24][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12257_  (.CLK(clknet_leaf_37_wb_clk_i),
    .D(\u_cpu.REG_FILE._00813_ ),
    .Q(\u_cpu.REG_FILE.rf[24][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12258_  (.CLK(clknet_leaf_38_wb_clk_i),
    .D(\u_cpu.REG_FILE._00814_ ),
    .Q(\u_cpu.REG_FILE.rf[24][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12259_  (.CLK(clknet_leaf_27_wb_clk_i),
    .D(\u_cpu.REG_FILE._00815_ ),
    .Q(\u_cpu.REG_FILE.rf[24][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12260_  (.CLK(clknet_leaf_32_wb_clk_i),
    .D(\u_cpu.REG_FILE._00816_ ),
    .Q(\u_cpu.REG_FILE.rf[24][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12261_  (.CLK(clknet_leaf_36_wb_clk_i),
    .D(\u_cpu.REG_FILE._00817_ ),
    .Q(\u_cpu.REG_FILE.rf[24][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12262_  (.CLK(clknet_leaf_32_wb_clk_i),
    .D(\u_cpu.REG_FILE._00818_ ),
    .Q(\u_cpu.REG_FILE.rf[24][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12263_  (.CLK(clknet_leaf_32_wb_clk_i),
    .D(\u_cpu.REG_FILE._00819_ ),
    .Q(\u_cpu.REG_FILE.rf[24][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12264_  (.CLK(clknet_leaf_58_wb_clk_i),
    .D(\u_cpu.REG_FILE._00820_ ),
    .Q(\u_cpu.REG_FILE.rf[24][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12265_  (.CLK(clknet_leaf_56_wb_clk_i),
    .D(\u_cpu.REG_FILE._00821_ ),
    .Q(\u_cpu.REG_FILE.rf[24][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12266_  (.CLK(clknet_leaf_53_wb_clk_i),
    .D(\u_cpu.REG_FILE._00822_ ),
    .Q(\u_cpu.REG_FILE.rf[24][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12267_  (.CLK(clknet_leaf_57_wb_clk_i),
    .D(\u_cpu.REG_FILE._00823_ ),
    .Q(\u_cpu.REG_FILE.rf[24][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12268_  (.CLK(clknet_leaf_53_wb_clk_i),
    .D(\u_cpu.REG_FILE._00824_ ),
    .Q(\u_cpu.REG_FILE.rf[24][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12269_  (.CLK(clknet_leaf_54_wb_clk_i),
    .D(\u_cpu.REG_FILE._00825_ ),
    .Q(\u_cpu.REG_FILE.rf[24][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12270_  (.CLK(clknet_leaf_56_wb_clk_i),
    .D(\u_cpu.REG_FILE._00826_ ),
    .Q(\u_cpu.REG_FILE.rf[24][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12271_  (.CLK(clknet_leaf_54_wb_clk_i),
    .D(\u_cpu.REG_FILE._00827_ ),
    .Q(\u_cpu.REG_FILE.rf[24][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12272_  (.CLK(clknet_leaf_53_wb_clk_i),
    .D(\u_cpu.REG_FILE._00828_ ),
    .Q(\u_cpu.REG_FILE.rf[24][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12273_  (.CLK(clknet_leaf_53_wb_clk_i),
    .D(\u_cpu.REG_FILE._00829_ ),
    .Q(\u_cpu.REG_FILE.rf[24][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12274_  (.CLK(clknet_leaf_31_wb_clk_i),
    .D(\u_cpu.REG_FILE._00830_ ),
    .Q(\u_cpu.REG_FILE.rf[24][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12275_  (.CLK(clknet_leaf_40_wb_clk_i),
    .D(\u_cpu.REG_FILE._00831_ ),
    .Q(\u_cpu.REG_FILE.rf[24][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12276_  (.CLK(clknet_leaf_18_wb_clk_i),
    .D(\u_cpu.REG_FILE._00832_ ),
    .Q(\u_cpu.REG_FILE.rf[25][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12277_  (.CLK(clknet_leaf_0_wb_clk_i),
    .D(\u_cpu.REG_FILE._00833_ ),
    .Q(\u_cpu.REG_FILE.rf[25][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12278_  (.CLK(clknet_leaf_18_wb_clk_i),
    .D(\u_cpu.REG_FILE._00834_ ),
    .Q(\u_cpu.REG_FILE.rf[25][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12279_  (.CLK(clknet_leaf_11_wb_clk_i),
    .D(\u_cpu.REG_FILE._00835_ ),
    .Q(\u_cpu.REG_FILE.rf[25][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12280_  (.CLK(clknet_leaf_14_wb_clk_i),
    .D(\u_cpu.REG_FILE._00836_ ),
    .Q(\u_cpu.REG_FILE.rf[25][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12281_  (.CLK(clknet_leaf_17_wb_clk_i),
    .D(\u_cpu.REG_FILE._00837_ ),
    .Q(\u_cpu.REG_FILE.rf[25][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12282_  (.CLK(clknet_leaf_0_wb_clk_i),
    .D(\u_cpu.REG_FILE._00838_ ),
    .Q(\u_cpu.REG_FILE.rf[25][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12283_  (.CLK(clknet_leaf_12_wb_clk_i),
    .D(\u_cpu.REG_FILE._00839_ ),
    .Q(\u_cpu.REG_FILE.rf[25][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12284_  (.CLK(clknet_leaf_6_wb_clk_i),
    .D(\u_cpu.REG_FILE._00840_ ),
    .Q(\u_cpu.REG_FILE.rf[25][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12285_  (.CLK(clknet_leaf_17_wb_clk_i),
    .D(\u_cpu.REG_FILE._00841_ ),
    .Q(\u_cpu.REG_FILE.rf[25][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12286_  (.CLK(clknet_leaf_16_wb_clk_i),
    .D(\u_cpu.REG_FILE._00842_ ),
    .Q(\u_cpu.REG_FILE.rf[25][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12287_  (.CLK(clknet_leaf_35_wb_clk_i),
    .D(\u_cpu.REG_FILE._00843_ ),
    .Q(\u_cpu.REG_FILE.rf[25][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12288_  (.CLK(clknet_leaf_38_wb_clk_i),
    .D(\u_cpu.REG_FILE._00844_ ),
    .Q(\u_cpu.REG_FILE.rf[25][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12289_  (.CLK(clknet_leaf_37_wb_clk_i),
    .D(\u_cpu.REG_FILE._00845_ ),
    .Q(\u_cpu.REG_FILE.rf[25][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12290_  (.CLK(clknet_leaf_38_wb_clk_i),
    .D(\u_cpu.REG_FILE._00846_ ),
    .Q(\u_cpu.REG_FILE.rf[25][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12291_  (.CLK(clknet_leaf_27_wb_clk_i),
    .D(\u_cpu.REG_FILE._00847_ ),
    .Q(\u_cpu.REG_FILE.rf[25][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12292_  (.CLK(clknet_leaf_32_wb_clk_i),
    .D(\u_cpu.REG_FILE._00848_ ),
    .Q(\u_cpu.REG_FILE.rf[25][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12293_  (.CLK(clknet_leaf_36_wb_clk_i),
    .D(\u_cpu.REG_FILE._00849_ ),
    .Q(\u_cpu.REG_FILE.rf[25][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12294_  (.CLK(clknet_leaf_32_wb_clk_i),
    .D(\u_cpu.REG_FILE._00850_ ),
    .Q(\u_cpu.REG_FILE.rf[25][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12295_  (.CLK(clknet_leaf_33_wb_clk_i),
    .D(\u_cpu.REG_FILE._00851_ ),
    .Q(\u_cpu.REG_FILE.rf[25][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12296_  (.CLK(clknet_leaf_58_wb_clk_i),
    .D(\u_cpu.REG_FILE._00852_ ),
    .Q(\u_cpu.REG_FILE.rf[25][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12297_  (.CLK(clknet_leaf_58_wb_clk_i),
    .D(\u_cpu.REG_FILE._00853_ ),
    .Q(\u_cpu.REG_FILE.rf[25][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12298_  (.CLK(clknet_leaf_53_wb_clk_i),
    .D(\u_cpu.REG_FILE._00854_ ),
    .Q(\u_cpu.REG_FILE.rf[25][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12299_  (.CLK(clknet_leaf_58_wb_clk_i),
    .D(\u_cpu.REG_FILE._00855_ ),
    .Q(\u_cpu.REG_FILE.rf[25][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12300_  (.CLK(clknet_leaf_53_wb_clk_i),
    .D(\u_cpu.REG_FILE._00856_ ),
    .Q(\u_cpu.REG_FILE.rf[25][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12301_  (.CLK(clknet_leaf_40_wb_clk_i),
    .D(\u_cpu.REG_FILE._00857_ ),
    .Q(\u_cpu.REG_FILE.rf[25][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12302_  (.CLK(clknet_leaf_53_wb_clk_i),
    .D(\u_cpu.REG_FILE._00858_ ),
    .Q(\u_cpu.REG_FILE.rf[25][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12303_  (.CLK(clknet_leaf_53_wb_clk_i),
    .D(\u_cpu.REG_FILE._00859_ ),
    .Q(\u_cpu.REG_FILE.rf[25][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12304_  (.CLK(clknet_leaf_53_wb_clk_i),
    .D(\u_cpu.REG_FILE._00860_ ),
    .Q(\u_cpu.REG_FILE.rf[25][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12305_  (.CLK(clknet_leaf_46_wb_clk_i),
    .D(\u_cpu.REG_FILE._00861_ ),
    .Q(\u_cpu.REG_FILE.rf[25][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12306_  (.CLK(clknet_leaf_33_wb_clk_i),
    .D(\u_cpu.REG_FILE._00862_ ),
    .Q(\u_cpu.REG_FILE.rf[25][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12307_  (.CLK(clknet_leaf_39_wb_clk_i),
    .D(\u_cpu.REG_FILE._00863_ ),
    .Q(\u_cpu.REG_FILE.rf[25][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12308_  (.CLK(clknet_leaf_0_wb_clk_i),
    .D(\u_cpu.REG_FILE._00864_ ),
    .Q(\u_cpu.REG_FILE.rf[26][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12309_  (.CLK(clknet_leaf_0_wb_clk_i),
    .D(\u_cpu.REG_FILE._00865_ ),
    .Q(\u_cpu.REG_FILE.rf[26][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12310_  (.CLK(clknet_leaf_18_wb_clk_i),
    .D(\u_cpu.REG_FILE._00866_ ),
    .Q(\u_cpu.REG_FILE.rf[26][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12311_  (.CLK(clknet_leaf_11_wb_clk_i),
    .D(\u_cpu.REG_FILE._00867_ ),
    .Q(\u_cpu.REG_FILE.rf[26][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12312_  (.CLK(clknet_leaf_14_wb_clk_i),
    .D(\u_cpu.REG_FILE._00868_ ),
    .Q(\u_cpu.REG_FILE.rf[26][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12313_  (.CLK(clknet_leaf_18_wb_clk_i),
    .D(\u_cpu.REG_FILE._00869_ ),
    .Q(\u_cpu.REG_FILE.rf[26][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12314_  (.CLK(clknet_leaf_0_wb_clk_i),
    .D(\u_cpu.REG_FILE._00870_ ),
    .Q(\u_cpu.REG_FILE.rf[26][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12315_  (.CLK(clknet_leaf_8_wb_clk_i),
    .D(\u_cpu.REG_FILE._00871_ ),
    .Q(\u_cpu.REG_FILE.rf[26][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12316_  (.CLK(clknet_leaf_6_wb_clk_i),
    .D(\u_cpu.REG_FILE._00872_ ),
    .Q(\u_cpu.REG_FILE.rf[26][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12317_  (.CLK(clknet_leaf_17_wb_clk_i),
    .D(\u_cpu.REG_FILE._00873_ ),
    .Q(\u_cpu.REG_FILE.rf[26][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12318_  (.CLK(clknet_leaf_16_wb_clk_i),
    .D(\u_cpu.REG_FILE._00874_ ),
    .Q(\u_cpu.REG_FILE.rf[26][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12319_  (.CLK(clknet_leaf_32_wb_clk_i),
    .D(\u_cpu.REG_FILE._00875_ ),
    .Q(\u_cpu.REG_FILE.rf[26][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12320_  (.CLK(clknet_leaf_15_wb_clk_i),
    .D(\u_cpu.REG_FILE._00876_ ),
    .Q(\u_cpu.REG_FILE.rf[26][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12321_  (.CLK(clknet_leaf_15_wb_clk_i),
    .D(\u_cpu.REG_FILE._00877_ ),
    .Q(\u_cpu.REG_FILE.rf[26][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12322_  (.CLK(clknet_leaf_38_wb_clk_i),
    .D(\u_cpu.REG_FILE._00878_ ),
    .Q(\u_cpu.REG_FILE.rf[26][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12323_  (.CLK(clknet_leaf_27_wb_clk_i),
    .D(\u_cpu.REG_FILE._00879_ ),
    .Q(\u_cpu.REG_FILE.rf[26][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12324_  (.CLK(clknet_leaf_32_wb_clk_i),
    .D(\u_cpu.REG_FILE._00880_ ),
    .Q(\u_cpu.REG_FILE.rf[26][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12325_  (.CLK(clknet_leaf_36_wb_clk_i),
    .D(\u_cpu.REG_FILE._00881_ ),
    .Q(\u_cpu.REG_FILE.rf[26][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12326_  (.CLK(clknet_leaf_32_wb_clk_i),
    .D(\u_cpu.REG_FILE._00882_ ),
    .Q(\u_cpu.REG_FILE.rf[26][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12327_  (.CLK(clknet_leaf_31_wb_clk_i),
    .D(\u_cpu.REG_FILE._00883_ ),
    .Q(\u_cpu.REG_FILE.rf[26][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12328_  (.CLK(clknet_leaf_58_wb_clk_i),
    .D(\u_cpu.REG_FILE._00884_ ),
    .Q(\u_cpu.REG_FILE.rf[26][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12329_  (.CLK(clknet_leaf_58_wb_clk_i),
    .D(\u_cpu.REG_FILE._00885_ ),
    .Q(\u_cpu.REG_FILE.rf[26][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12330_  (.CLK(clknet_leaf_53_wb_clk_i),
    .D(\u_cpu.REG_FILE._00886_ ),
    .Q(\u_cpu.REG_FILE.rf[26][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12331_  (.CLK(clknet_leaf_58_wb_clk_i),
    .D(\u_cpu.REG_FILE._00887_ ),
    .Q(\u_cpu.REG_FILE.rf[26][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12332_  (.CLK(clknet_leaf_53_wb_clk_i),
    .D(\u_cpu.REG_FILE._00888_ ),
    .Q(\u_cpu.REG_FILE.rf[26][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12333_  (.CLK(clknet_leaf_33_wb_clk_i),
    .D(\u_cpu.REG_FILE._00889_ ),
    .Q(\u_cpu.REG_FILE.rf[26][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12334_  (.CLK(clknet_leaf_53_wb_clk_i),
    .D(\u_cpu.REG_FILE._00890_ ),
    .Q(\u_cpu.REG_FILE.rf[26][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12335_  (.CLK(clknet_leaf_53_wb_clk_i),
    .D(\u_cpu.REG_FILE._00891_ ),
    .Q(\u_cpu.REG_FILE.rf[26][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12336_  (.CLK(clknet_leaf_53_wb_clk_i),
    .D(\u_cpu.REG_FILE._00892_ ),
    .Q(\u_cpu.REG_FILE.rf[26][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12337_  (.CLK(clknet_leaf_53_wb_clk_i),
    .D(\u_cpu.REG_FILE._00893_ ),
    .Q(\u_cpu.REG_FILE.rf[26][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12338_  (.CLK(clknet_leaf_33_wb_clk_i),
    .D(\u_cpu.REG_FILE._00894_ ),
    .Q(\u_cpu.REG_FILE.rf[26][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12339_  (.CLK(clknet_leaf_34_wb_clk_i),
    .D(\u_cpu.REG_FILE._00895_ ),
    .Q(\u_cpu.REG_FILE.rf[26][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12340_  (.CLK(clknet_leaf_0_wb_clk_i),
    .D(\u_cpu.REG_FILE._00896_ ),
    .Q(\u_cpu.REG_FILE.rf[27][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12341_  (.CLK(clknet_leaf_0_wb_clk_i),
    .D(\u_cpu.REG_FILE._00897_ ),
    .Q(\u_cpu.REG_FILE.rf[27][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12342_  (.CLK(clknet_leaf_18_wb_clk_i),
    .D(\u_cpu.REG_FILE._00898_ ),
    .Q(\u_cpu.REG_FILE.rf[27][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12343_  (.CLK(clknet_leaf_11_wb_clk_i),
    .D(\u_cpu.REG_FILE._00899_ ),
    .Q(\u_cpu.REG_FILE.rf[27][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12344_  (.CLK(clknet_leaf_14_wb_clk_i),
    .D(\u_cpu.REG_FILE._00900_ ),
    .Q(\u_cpu.REG_FILE.rf[27][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12345_  (.CLK(clknet_leaf_17_wb_clk_i),
    .D(\u_cpu.REG_FILE._00901_ ),
    .Q(\u_cpu.REG_FILE.rf[27][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12346_  (.CLK(clknet_leaf_0_wb_clk_i),
    .D(\u_cpu.REG_FILE._00902_ ),
    .Q(\u_cpu.REG_FILE.rf[27][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12347_  (.CLK(clknet_leaf_7_wb_clk_i),
    .D(\u_cpu.REG_FILE._00903_ ),
    .Q(\u_cpu.REG_FILE.rf[27][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12348_  (.CLK(clknet_leaf_0_wb_clk_i),
    .D(\u_cpu.REG_FILE._00904_ ),
    .Q(\u_cpu.REG_FILE.rf[27][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12349_  (.CLK(clknet_leaf_17_wb_clk_i),
    .D(\u_cpu.REG_FILE._00905_ ),
    .Q(\u_cpu.REG_FILE.rf[27][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12350_  (.CLK(clknet_leaf_15_wb_clk_i),
    .D(\u_cpu.REG_FILE._00906_ ),
    .Q(\u_cpu.REG_FILE.rf[27][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12351_  (.CLK(clknet_leaf_32_wb_clk_i),
    .D(\u_cpu.REG_FILE._00907_ ),
    .Q(\u_cpu.REG_FILE.rf[27][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12352_  (.CLK(clknet_leaf_38_wb_clk_i),
    .D(\u_cpu.REG_FILE._00908_ ),
    .Q(\u_cpu.REG_FILE.rf[27][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12353_  (.CLK(clknet_leaf_15_wb_clk_i),
    .D(\u_cpu.REG_FILE._00909_ ),
    .Q(\u_cpu.REG_FILE.rf[27][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12354_  (.CLK(clknet_leaf_38_wb_clk_i),
    .D(\u_cpu.REG_FILE._00910_ ),
    .Q(\u_cpu.REG_FILE.rf[27][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12355_  (.CLK(clknet_leaf_27_wb_clk_i),
    .D(\u_cpu.REG_FILE._00911_ ),
    .Q(\u_cpu.REG_FILE.rf[27][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12356_  (.CLK(clknet_leaf_32_wb_clk_i),
    .D(\u_cpu.REG_FILE._00912_ ),
    .Q(\u_cpu.REG_FILE.rf[27][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12357_  (.CLK(clknet_leaf_28_wb_clk_i),
    .D(\u_cpu.REG_FILE._00913_ ),
    .Q(\u_cpu.REG_FILE.rf[27][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12358_  (.CLK(clknet_leaf_29_wb_clk_i),
    .D(\u_cpu.REG_FILE._00914_ ),
    .Q(\u_cpu.REG_FILE.rf[27][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12359_  (.CLK(clknet_leaf_32_wb_clk_i),
    .D(\u_cpu.REG_FILE._00915_ ),
    .Q(\u_cpu.REG_FILE.rf[27][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12360_  (.CLK(clknet_leaf_58_wb_clk_i),
    .D(\u_cpu.REG_FILE._00916_ ),
    .Q(\u_cpu.REG_FILE.rf[27][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12361_  (.CLK(clknet_leaf_56_wb_clk_i),
    .D(\u_cpu.REG_FILE._00917_ ),
    .Q(\u_cpu.REG_FILE.rf[27][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12362_  (.CLK(clknet_leaf_53_wb_clk_i),
    .D(\u_cpu.REG_FILE._00918_ ),
    .Q(\u_cpu.REG_FILE.rf[27][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12363_  (.CLK(clknet_leaf_58_wb_clk_i),
    .D(\u_cpu.REG_FILE._00919_ ),
    .Q(\u_cpu.REG_FILE.rf[27][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12364_  (.CLK(clknet_leaf_53_wb_clk_i),
    .D(\u_cpu.REG_FILE._00920_ ),
    .Q(\u_cpu.REG_FILE.rf[27][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12365_  (.CLK(clknet_leaf_31_wb_clk_i),
    .D(\u_cpu.REG_FILE._00921_ ),
    .Q(\u_cpu.REG_FILE.rf[27][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12366_  (.CLK(clknet_leaf_56_wb_clk_i),
    .D(\u_cpu.REG_FILE._00922_ ),
    .Q(\u_cpu.REG_FILE.rf[27][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12367_  (.CLK(clknet_leaf_33_wb_clk_i),
    .D(\u_cpu.REG_FILE._00923_ ),
    .Q(\u_cpu.REG_FILE.rf[27][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12368_  (.CLK(clknet_leaf_53_wb_clk_i),
    .D(\u_cpu.REG_FILE._00924_ ),
    .Q(\u_cpu.REG_FILE.rf[27][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12369_  (.CLK(clknet_leaf_53_wb_clk_i),
    .D(\u_cpu.REG_FILE._00925_ ),
    .Q(\u_cpu.REG_FILE.rf[27][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12370_  (.CLK(clknet_leaf_33_wb_clk_i),
    .D(\u_cpu.REG_FILE._00926_ ),
    .Q(\u_cpu.REG_FILE.rf[27][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12371_  (.CLK(clknet_leaf_34_wb_clk_i),
    .D(\u_cpu.REG_FILE._00927_ ),
    .Q(\u_cpu.REG_FILE.rf[27][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12372_  (.CLK(clknet_leaf_2_wb_clk_i),
    .D(\u_cpu.REG_FILE._00928_ ),
    .Q(\u_cpu.REG_FILE.rf[28][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12373_  (.CLK(clknet_leaf_2_wb_clk_i),
    .D(\u_cpu.REG_FILE._00929_ ),
    .Q(\u_cpu.REG_FILE.rf[28][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12374_  (.CLK(clknet_leaf_4_wb_clk_i),
    .D(\u_cpu.REG_FILE._00930_ ),
    .Q(\u_cpu.REG_FILE.rf[28][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12375_  (.CLK(clknet_leaf_10_wb_clk_i),
    .D(\u_cpu.REG_FILE._00931_ ),
    .Q(\u_cpu.REG_FILE.rf[28][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12376_  (.CLK(clknet_leaf_4_wb_clk_i),
    .D(\u_cpu.REG_FILE._00932_ ),
    .Q(\u_cpu.REG_FILE.rf[28][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12377_  (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\u_cpu.REG_FILE._00933_ ),
    .Q(\u_cpu.REG_FILE.rf[28][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12378_  (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\u_cpu.REG_FILE._00934_ ),
    .Q(\u_cpu.REG_FILE.rf[28][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12379_  (.CLK(clknet_leaf_114_wb_clk_i),
    .D(\u_cpu.REG_FILE._00935_ ),
    .Q(\u_cpu.REG_FILE.rf[28][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12380_  (.CLK(clknet_leaf_117_wb_clk_i),
    .D(\u_cpu.REG_FILE._00936_ ),
    .Q(\u_cpu.REG_FILE.rf[28][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12381_  (.CLK(clknet_leaf_5_wb_clk_i),
    .D(\u_cpu.REG_FILE._00937_ ),
    .Q(\u_cpu.REG_FILE.rf[28][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12382_  (.CLK(clknet_leaf_3_wb_clk_i),
    .D(\u_cpu.REG_FILE._00938_ ),
    .Q(\u_cpu.REG_FILE.rf[28][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12383_  (.CLK(clknet_leaf_39_wb_clk_i),
    .D(\u_cpu.REG_FILE._00939_ ),
    .Q(\u_cpu.REG_FILE.rf[28][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12384_  (.CLK(clknet_leaf_118_wb_clk_i),
    .D(\u_cpu.REG_FILE._00940_ ),
    .Q(\u_cpu.REG_FILE.rf[28][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12385_  (.CLK(clknet_leaf_118_wb_clk_i),
    .D(\u_cpu.REG_FILE._00941_ ),
    .Q(\u_cpu.REG_FILE.rf[28][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12386_  (.CLK(clknet_leaf_117_wb_clk_i),
    .D(\u_cpu.REG_FILE._00942_ ),
    .Q(\u_cpu.REG_FILE.rf[28][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12387_  (.CLK(clknet_leaf_37_wb_clk_i),
    .D(\u_cpu.REG_FILE._00943_ ),
    .Q(\u_cpu.REG_FILE.rf[28][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12388_  (.CLK(clknet_leaf_34_wb_clk_i),
    .D(\u_cpu.REG_FILE._00944_ ),
    .Q(\u_cpu.REG_FILE.rf[28][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12389_  (.CLK(clknet_leaf_27_wb_clk_i),
    .D(\u_cpu.REG_FILE._00945_ ),
    .Q(\u_cpu.REG_FILE.rf[28][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12390_  (.CLK(clknet_leaf_35_wb_clk_i),
    .D(\u_cpu.REG_FILE._00946_ ),
    .Q(\u_cpu.REG_FILE.rf[28][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12391_  (.CLK(clknet_leaf_33_wb_clk_i),
    .D(\u_cpu.REG_FILE._00947_ ),
    .Q(\u_cpu.REG_FILE.rf[28][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12392_  (.CLK(clknet_leaf_50_wb_clk_i),
    .D(\u_cpu.REG_FILE._00948_ ),
    .Q(\u_cpu.REG_FILE.rf[28][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12393_  (.CLK(clknet_leaf_76_wb_clk_i),
    .D(\u_cpu.REG_FILE._00949_ ),
    .Q(\u_cpu.REG_FILE.rf[28][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12394_  (.CLK(clknet_leaf_45_wb_clk_i),
    .D(\u_cpu.REG_FILE._00950_ ),
    .Q(\u_cpu.REG_FILE.rf[28][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12395_  (.CLK(clknet_leaf_48_wb_clk_i),
    .D(\u_cpu.REG_FILE._00951_ ),
    .Q(\u_cpu.REG_FILE.rf[28][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12396_  (.CLK(clknet_leaf_52_wb_clk_i),
    .D(\u_cpu.REG_FILE._00952_ ),
    .Q(\u_cpu.REG_FILE.rf[28][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12397_  (.CLK(clknet_leaf_45_wb_clk_i),
    .D(\u_cpu.REG_FILE._00953_ ),
    .Q(\u_cpu.REG_FILE.rf[28][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12398_  (.CLK(clknet_leaf_50_wb_clk_i),
    .D(\u_cpu.REG_FILE._00954_ ),
    .Q(\u_cpu.REG_FILE.rf[28][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12399_  (.CLK(clknet_leaf_34_wb_clk_i),
    .D(\u_cpu.REG_FILE._00955_ ),
    .Q(\u_cpu.REG_FILE.rf[28][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12400_  (.CLK(clknet_leaf_52_wb_clk_i),
    .D(\u_cpu.REG_FILE._00956_ ),
    .Q(\u_cpu.REG_FILE.rf[28][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12401_  (.CLK(clknet_leaf_43_wb_clk_i),
    .D(\u_cpu.REG_FILE._00957_ ),
    .Q(\u_cpu.REG_FILE.rf[28][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12402_  (.CLK(clknet_leaf_42_wb_clk_i),
    .D(\u_cpu.REG_FILE._00958_ ),
    .Q(\u_cpu.REG_FILE.rf[28][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12403_  (.CLK(clknet_leaf_42_wb_clk_i),
    .D(\u_cpu.REG_FILE._00959_ ),
    .Q(\u_cpu.REG_FILE.rf[28][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12404_  (.CLK(clknet_leaf_127_wb_clk_i),
    .D(\u_cpu.REG_FILE._00960_ ),
    .Q(\u_cpu.REG_FILE.rf[2][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12405_  (.CLK(clknet_leaf_127_wb_clk_i),
    .D(\u_cpu.REG_FILE._00961_ ),
    .Q(\u_cpu.REG_FILE.rf[2][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12406_  (.CLK(clknet_leaf_127_wb_clk_i),
    .D(\u_cpu.REG_FILE._00962_ ),
    .Q(\u_cpu.REG_FILE.rf[2][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12407_  (.CLK(clknet_leaf_117_wb_clk_i),
    .D(\u_cpu.REG_FILE._00963_ ),
    .Q(\u_cpu.REG_FILE.rf[2][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12408_  (.CLK(clknet_leaf_120_wb_clk_i),
    .D(\u_cpu.REG_FILE._00964_ ),
    .Q(\u_cpu.REG_FILE.rf[2][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12409_  (.CLK(clknet_leaf_119_wb_clk_i),
    .D(\u_cpu.REG_FILE._00965_ ),
    .Q(\u_cpu.REG_FILE.rf[2][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12410_  (.CLK(clknet_leaf_127_wb_clk_i),
    .D(\u_cpu.REG_FILE._00966_ ),
    .Q(\u_cpu.REG_FILE.rf[2][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12411_  (.CLK(clknet_leaf_8_wb_clk_i),
    .D(\u_cpu.REG_FILE._00967_ ),
    .Q(\u_cpu.REG_FILE.rf[2][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12412_  (.CLK(clknet_leaf_127_wb_clk_i),
    .D(\u_cpu.REG_FILE._00968_ ),
    .Q(\u_cpu.REG_FILE.rf[2][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12413_  (.CLK(clknet_leaf_8_wb_clk_i),
    .D(\u_cpu.REG_FILE._00969_ ),
    .Q(\u_cpu.REG_FILE.rf[2][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12414_  (.CLK(clknet_leaf_99_wb_clk_i),
    .D(\u_cpu.REG_FILE._00970_ ),
    .Q(\u_cpu.REG_FILE.rf[2][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12415_  (.CLK(clknet_leaf_77_wb_clk_i),
    .D(\u_cpu.REG_FILE._00971_ ),
    .Q(\u_cpu.REG_FILE.rf[2][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12416_  (.CLK(clknet_leaf_93_wb_clk_i),
    .D(\u_cpu.REG_FILE._00972_ ),
    .Q(\u_cpu.REG_FILE.rf[2][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12417_  (.CLK(clknet_leaf_92_wb_clk_i),
    .D(\u_cpu.REG_FILE._00973_ ),
    .Q(\u_cpu.REG_FILE.rf[2][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12418_  (.CLK(clknet_leaf_91_wb_clk_i),
    .D(\u_cpu.REG_FILE._00974_ ),
    .Q(\u_cpu.REG_FILE.rf[2][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12419_  (.CLK(clknet_leaf_100_wb_clk_i),
    .D(\u_cpu.REG_FILE._00975_ ),
    .Q(\u_cpu.REG_FILE.rf[2][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12420_  (.CLK(clknet_leaf_109_wb_clk_i),
    .D(\u_cpu.REG_FILE._00976_ ),
    .Q(\u_cpu.REG_FILE.rf[2][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12421_  (.CLK(clknet_leaf_105_wb_clk_i),
    .D(\u_cpu.REG_FILE._00977_ ),
    .Q(\u_cpu.REG_FILE.rf[2][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12422_  (.CLK(clknet_leaf_49_wb_clk_i),
    .D(\u_cpu.REG_FILE._00978_ ),
    .Q(\u_cpu.REG_FILE.rf[2][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12423_  (.CLK(clknet_leaf_44_wb_clk_i),
    .D(\u_cpu.REG_FILE._00979_ ),
    .Q(\u_cpu.REG_FILE.rf[2][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12424_  (.CLK(clknet_leaf_50_wb_clk_i),
    .D(\u_cpu.REG_FILE._00980_ ),
    .Q(\u_cpu.REG_FILE.rf[2][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12425_  (.CLK(clknet_leaf_47_wb_clk_i),
    .D(\u_cpu.REG_FILE._00981_ ),
    .Q(\u_cpu.REG_FILE.rf[2][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12426_  (.CLK(clknet_leaf_48_wb_clk_i),
    .D(\u_cpu.REG_FILE._00982_ ),
    .Q(\u_cpu.REG_FILE.rf[2][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12427_  (.CLK(clknet_leaf_73_wb_clk_i),
    .D(\u_cpu.REG_FILE._00983_ ),
    .Q(\u_cpu.REG_FILE.rf[2][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12428_  (.CLK(clknet_leaf_59_wb_clk_i),
    .D(\u_cpu.REG_FILE._00984_ ),
    .Q(\u_cpu.REG_FILE.rf[2][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12429_  (.CLK(clknet_leaf_49_wb_clk_i),
    .D(\u_cpu.REG_FILE._00985_ ),
    .Q(\u_cpu.REG_FILE.rf[2][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12430_  (.CLK(clknet_leaf_59_wb_clk_i),
    .D(\u_cpu.REG_FILE._00986_ ),
    .Q(\u_cpu.REG_FILE.rf[2][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12431_  (.CLK(clknet_leaf_59_wb_clk_i),
    .D(\u_cpu.REG_FILE._00987_ ),
    .Q(\u_cpu.REG_FILE.rf[2][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12432_  (.CLK(clknet_leaf_59_wb_clk_i),
    .D(\u_cpu.REG_FILE._00988_ ),
    .Q(\u_cpu.REG_FILE.rf[2][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12433_  (.CLK(clknet_leaf_63_wb_clk_i),
    .D(\u_cpu.REG_FILE._00989_ ),
    .Q(\u_cpu.REG_FILE.rf[2][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12434_  (.CLK(clknet_leaf_9_wb_clk_i),
    .D(\u_cpu.REG_FILE._00990_ ),
    .Q(\u_cpu.REG_FILE.rf[2][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12435_  (.CLK(clknet_leaf_74_wb_clk_i),
    .D(\u_cpu.REG_FILE._00991_ ),
    .Q(\u_cpu.REG_FILE.rf[2][31] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12436_  (.CLK(clknet_leaf_128_wb_clk_i),
    .D(\u_cpu.REG_FILE._00992_ ),
    .Q(\u_cpu.REG_FILE.rf[30][0] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12437_  (.CLK(clknet_leaf_129_wb_clk_i),
    .D(\u_cpu.REG_FILE._00993_ ),
    .Q(\u_cpu.REG_FILE.rf[30][1] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12438_  (.CLK(clknet_leaf_128_wb_clk_i),
    .D(\u_cpu.REG_FILE._00994_ ),
    .Q(\u_cpu.REG_FILE.rf[30][2] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12439_  (.CLK(clknet_leaf_114_wb_clk_i),
    .D(\u_cpu.REG_FILE._00995_ ),
    .Q(\u_cpu.REG_FILE.rf[30][3] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12440_  (.CLK(clknet_leaf_119_wb_clk_i),
    .D(\u_cpu.REG_FILE._00996_ ),
    .Q(\u_cpu.REG_FILE.rf[30][4] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12441_  (.CLK(clknet_leaf_128_wb_clk_i),
    .D(\u_cpu.REG_FILE._00997_ ),
    .Q(\u_cpu.REG_FILE.rf[30][5] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12442_  (.CLK(clknet_leaf_129_wb_clk_i),
    .D(\u_cpu.REG_FILE._00998_ ),
    .Q(\u_cpu.REG_FILE.rf[30][6] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12443_  (.CLK(clknet_leaf_5_wb_clk_i),
    .D(\u_cpu.REG_FILE._00999_ ),
    .Q(\u_cpu.REG_FILE.rf[30][7] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12444_  (.CLK(clknet_leaf_128_wb_clk_i),
    .D(\u_cpu.REG_FILE._01000_ ),
    .Q(\u_cpu.REG_FILE.rf[30][8] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12445_  (.CLK(clknet_leaf_6_wb_clk_i),
    .D(\u_cpu.REG_FILE._01001_ ),
    .Q(\u_cpu.REG_FILE.rf[30][9] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12446_  (.CLK(clknet_leaf_118_wb_clk_i),
    .D(\u_cpu.REG_FILE._01002_ ),
    .Q(\u_cpu.REG_FILE.rf[30][10] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12447_  (.CLK(clknet_leaf_38_wb_clk_i),
    .D(\u_cpu.REG_FILE._01003_ ),
    .Q(\u_cpu.REG_FILE.rf[30][11] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12448_  (.CLK(clknet_leaf_118_wb_clk_i),
    .D(\u_cpu.REG_FILE._01004_ ),
    .Q(\u_cpu.REG_FILE.rf[30][12] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12449_  (.CLK(clknet_leaf_119_wb_clk_i),
    .D(\u_cpu.REG_FILE._01005_ ),
    .Q(\u_cpu.REG_FILE.rf[30][13] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12450_  (.CLK(clknet_leaf_121_wb_clk_i),
    .D(\u_cpu.REG_FILE._01006_ ),
    .Q(\u_cpu.REG_FILE.rf[30][14] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12451_  (.CLK(clknet_leaf_37_wb_clk_i),
    .D(\u_cpu.REG_FILE._01007_ ),
    .Q(\u_cpu.REG_FILE.rf[30][15] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12452_  (.CLK(clknet_leaf_39_wb_clk_i),
    .D(\u_cpu.REG_FILE._01008_ ),
    .Q(\u_cpu.REG_FILE.rf[30][16] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12453_  (.CLK(clknet_leaf_36_wb_clk_i),
    .D(\u_cpu.REG_FILE._01009_ ),
    .Q(\u_cpu.REG_FILE.rf[30][17] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12454_  (.CLK(clknet_leaf_35_wb_clk_i),
    .D(\u_cpu.REG_FILE._01010_ ),
    .Q(\u_cpu.REG_FILE.rf[30][18] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12455_  (.CLK(clknet_leaf_34_wb_clk_i),
    .D(\u_cpu.REG_FILE._01011_ ),
    .Q(\u_cpu.REG_FILE.rf[30][19] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12456_  (.CLK(clknet_leaf_50_wb_clk_i),
    .D(\u_cpu.REG_FILE._01012_ ),
    .Q(\u_cpu.REG_FILE.rf[30][20] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12457_  (.CLK(clknet_leaf_72_wb_clk_i),
    .D(\u_cpu.REG_FILE._01013_ ),
    .Q(\u_cpu.REG_FILE.rf[30][21] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12458_  (.CLK(clknet_leaf_46_wb_clk_i),
    .D(\u_cpu.REG_FILE._01014_ ),
    .Q(\u_cpu.REG_FILE.rf[30][22] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12459_  (.CLK(clknet_leaf_48_wb_clk_i),
    .D(\u_cpu.REG_FILE._01015_ ),
    .Q(\u_cpu.REG_FILE.rf[30][23] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12460_  (.CLK(clknet_leaf_50_wb_clk_i),
    .D(\u_cpu.REG_FILE._01016_ ),
    .Q(\u_cpu.REG_FILE.rf[30][24] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12461_  (.CLK(clknet_leaf_45_wb_clk_i),
    .D(\u_cpu.REG_FILE._01017_ ),
    .Q(\u_cpu.REG_FILE.rf[30][25] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12462_  (.CLK(clknet_leaf_58_wb_clk_i),
    .D(\u_cpu.REG_FILE._01018_ ),
    .Q(\u_cpu.REG_FILE.rf[30][26] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12463_  (.CLK(clknet_leaf_49_wb_clk_i),
    .D(\u_cpu.REG_FILE._01019_ ),
    .Q(\u_cpu.REG_FILE.rf[30][27] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12464_  (.CLK(clknet_leaf_59_wb_clk_i),
    .D(\u_cpu.REG_FILE._01020_ ),
    .Q(\u_cpu.REG_FILE.rf[30][28] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12465_  (.CLK(clknet_leaf_45_wb_clk_i),
    .D(\u_cpu.REG_FILE._01021_ ),
    .Q(\u_cpu.REG_FILE.rf[30][29] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12466_  (.CLK(clknet_leaf_10_wb_clk_i),
    .D(\u_cpu.REG_FILE._01022_ ),
    .Q(\u_cpu.REG_FILE.rf[30][30] ));
 sky130_fd_sc_hd__dfxtp_2 \u_cpu.REG_FILE._12467_  (.CLK(clknet_leaf_43_wb_clk_i),
    .D(\u_cpu.REG_FILE._01023_ ),
    .Q(\u_cpu.REG_FILE.rf[30][31] ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0696_  (.A(\u_cpu.ALUResult_W_Reg[29] ),
    .B(\u_cpu.ALUResult_W_Reg[28] ),
    .Y(\u_cpu._0169_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0697_  (.A(\u_cpu.ALUResult_W_Reg[29] ),
    .B(\u_cpu.ALUResult_W_Reg[28] ),
    .X(\u_cpu._0170_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0698_  (.A(\u_cpu.ALUResult_W_Reg[25] ),
    .B(\u_cpu.ALUResult_W_Reg[24] ),
    .Y(\u_cpu._0171_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0699_  (.A(\u_cpu.ALUResult_W_Reg[25] ),
    .B(\u_cpu.ALUResult_W_Reg[24] ),
    .X(\u_cpu._0172_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu._0700_  (.A1(\u_cpu._0169_ ),
    .A2(\u_cpu._0170_ ),
    .B1(\u_cpu._0171_ ),
    .B2(\u_cpu._0172_ ),
    .Y(\u_cpu._0173_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu._0701_  (.A(\u_cpu._0169_ ),
    .B(\u_cpu._0170_ ),
    .C(\u_cpu._0171_ ),
    .D(\u_cpu._0172_ ),
    .X(\u_cpu._0174_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0702_  (.A(\u_cpu.ALUResult_W_Reg[19] ),
    .B(\u_cpu.ALUResult_W_Reg[18] ),
    .Y(\u_cpu._0175_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0703_  (.A(\u_cpu.ALUResult_W_Reg[19] ),
    .B(\u_cpu.ALUResult_W_Reg[18] ),
    .X(\u_cpu._0176_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0704_  (.A(\u_cpu.ALUResult_W_Reg[23] ),
    .B(\u_cpu.ALUResult_W_Reg[22] ),
    .Y(\u_cpu._0177_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0705_  (.A(\u_cpu.ALUResult_W_Reg[23] ),
    .B(\u_cpu.ALUResult_W_Reg[22] ),
    .X(\u_cpu._0178_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._0706_  (.A(\u_cpu._0175_ ),
    .B(\u_cpu._0176_ ),
    .C(\u_cpu._0177_ ),
    .D(\u_cpu._0178_ ),
    .Y(\u_cpu._0179_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0707_  (.A(\u_cpu.ALUResult_W_Reg[23] ),
    .B(\u_cpu.ALUResult_W_Reg[22] ),
    .X(\u_cpu._0180_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0708_  (.A(\u_cpu.ALUResult_W_Reg[23] ),
    .B(\u_cpu.ALUResult_W_Reg[22] ),
    .Y(\u_cpu._0181_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu._0709_  (.A1_N(\u_cpu._0175_ ),
    .A2_N(\u_cpu._0176_ ),
    .B1(\u_cpu._0180_ ),
    .B2(\u_cpu._0181_ ),
    .Y(\u_cpu._0182_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0710_  (.A(\u_cpu.ALUResult_W_Reg[21] ),
    .B(\u_cpu.ALUResult_W_Reg[20] ),
    .Y(\u_cpu._0183_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0711_  (.A(\u_cpu.ALUResult_W_Reg[21] ),
    .B(\u_cpu.ALUResult_W_Reg[20] ),
    .X(\u_cpu._0184_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0712_  (.A(\u_cpu.ALUResult_W_Reg[16] ),
    .B_N(\u_cpu.ALUResult_W_Reg[17] ),
    .X(\u_cpu._0185_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0713_  (.A(\u_cpu.ALUResult_W_Reg[17] ),
    .B_N(\u_cpu.ALUResult_W_Reg[16] ),
    .X(\u_cpu._0186_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu._0714_  (.A1_N(\u_cpu._0183_ ),
    .A2_N(\u_cpu._0184_ ),
    .B1(\u_cpu._0185_ ),
    .B2(\u_cpu._0186_ ),
    .Y(\u_cpu._0187_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0715_  (.A(\u_cpu.ALUResult_W_Reg[21] ),
    .B_N(\u_cpu.ALUResult_W_Reg[20] ),
    .X(\u_cpu._0188_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0716_  (.A(\u_cpu.ALUResult_W_Reg[20] ),
    .B_N(\u_cpu.ALUResult_W_Reg[21] ),
    .X(\u_cpu._0189_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0717_  (.A(\u_cpu.ALUResult_W_Reg[17] ),
    .B(\u_cpu.ALUResult_W_Reg[16] ),
    .Y(\u_cpu._0190_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0718_  (.A(\u_cpu.ALUResult_W_Reg[17] ),
    .B(\u_cpu.ALUResult_W_Reg[16] ),
    .X(\u_cpu._0191_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu._0719_  (.A1(\u_cpu._0188_ ),
    .A2(\u_cpu._0189_ ),
    .B1(\u_cpu._0190_ ),
    .B2(\u_cpu._0191_ ),
    .Y(\u_cpu._0192_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu._0720_  (.A1_N(\u_cpu._0179_ ),
    .A2_N(\u_cpu._0182_ ),
    .B1(\u_cpu._0187_ ),
    .B2(\u_cpu._0192_ ),
    .Y(\u_cpu._0193_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu._0721_  (.A1(\u_cpu._0183_ ),
    .A2(\u_cpu._0184_ ),
    .B1(\u_cpu._0190_ ),
    .C1(\u_cpu._0191_ ),
    .Y(\u_cpu._0194_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0722_  (.A(\u_cpu.ALUResult_W_Reg[21] ),
    .B(\u_cpu.ALUResult_W_Reg[20] ),
    .Y(\u_cpu._0195_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu._0723_  (.A_N(\u_cpu._0183_ ),
    .B(\u_cpu._0195_ ),
    .C(\u_cpu._0185_ ),
    .D(\u_cpu._0186_ ),
    .Y(\u_cpu._0196_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._0724_  (.A(\u_cpu._0179_ ),
    .B(\u_cpu._0182_ ),
    .C(\u_cpu._0194_ ),
    .D(\u_cpu._0196_ ),
    .Y(\u_cpu._0197_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu._0725_  (.A1(\u_cpu._0173_ ),
    .A2(\u_cpu._0174_ ),
    .B1(\u_cpu._0193_ ),
    .C1(\u_cpu._0197_ ),
    .X(\u_cpu._0198_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu._0726_  (.A1(\u_cpu._0169_ ),
    .A2(\u_cpu._0170_ ),
    .B1(\u_cpu._0171_ ),
    .B2(\u_cpu._0172_ ),
    .X(\u_cpu._0199_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._0727_  (.A(\u_cpu._0169_ ),
    .B(\u_cpu._0170_ ),
    .C(\u_cpu._0171_ ),
    .D(\u_cpu._0172_ ),
    .Y(\u_cpu._0200_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0728_  (.A(\u_cpu._0199_ ),
    .B(\u_cpu._0200_ ),
    .Y(\u_cpu._0201_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu._0729_  (.A1(\u_cpu._0193_ ),
    .A2(\u_cpu._0197_ ),
    .B1(\u_cpu._0201_ ),
    .X(\u_cpu._0202_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu._0730_  (.A(\u_cpu.ALUResult_W_Reg[31] ),
    .B(\u_cpu.ALUResult_W_Reg[30] ),
    .Y(\u_cpu._0203_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu._0731_  (.A(\u_cpu.ALUResult_W_Reg[27] ),
    .B(\u_cpu.ALUResult_W_Reg[26] ),
    .Y(\u_cpu._0204_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu._0732_  (.A(\u_cpu._0203_ ),
    .B(\u_cpu._0204_ ),
    .Y(\u_cpu._0205_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0733_  (.A(\u_cpu._0202_ ),
    .B(\u_cpu._0205_ ),
    .Y(\u_cpu._0206_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu._0734_  (.A1(\u_cpu._0193_ ),
    .A2(\u_cpu._0197_ ),
    .B1(\u_cpu._0201_ ),
    .Y(\u_cpu._0207_ ));
 sky130_fd_sc_hd__o21bai_2 \u_cpu._0735_  (.A1(\u_cpu._0207_ ),
    .A2(\u_cpu._0198_ ),
    .B1_N(\u_cpu._0205_ ),
    .Y(\u_cpu._0208_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu._0736_  (.A1(\u_cpu._0198_ ),
    .A2(\u_cpu._0206_ ),
    .B1(\u_cpu._0208_ ),
    .Y(\u_cpu._0209_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0737_  (.A(\u_cpu.ALUResult_W_Reg[13] ),
    .B(\u_cpu.ALUResult_W_Reg[12] ),
    .Y(\u_cpu._0210_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0738_  (.A(\u_cpu.ALUResult_W_Reg[13] ),
    .B(\u_cpu.ALUResult_W_Reg[12] ),
    .X(\u_cpu._0211_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0739_  (.A(\u_cpu.led[9] ),
    .B(\u_cpu.led[8] ),
    .Y(\u_cpu._0212_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0740_  (.A(\u_cpu.led[9] ),
    .B(\u_cpu.led[8] ),
    .X(\u_cpu._0213_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu._0741_  (.A1(\u_cpu._0210_ ),
    .A2(\u_cpu._0211_ ),
    .B1(\u_cpu._0212_ ),
    .B2(\u_cpu._0213_ ),
    .Y(\u_cpu._0214_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu._0742_  (.A(\u_cpu._0210_ ),
    .B(\u_cpu._0211_ ),
    .C(\u_cpu._0212_ ),
    .D(\u_cpu._0213_ ),
    .X(\u_cpu._0215_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu._0743_  (.A_N(\u_cpu.ALUResult_W_Reg[0] ),
    .B(\u_cpu.led[1] ),
    .X(\u_cpu._0216_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu._0744_  (.A(\u_cpu.ALUResult_W_Reg[0] ),
    .Y(\u_cpu._0217_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0745_  (.A(\u_cpu.led[5] ),
    .B(\u_cpu.led[4] ),
    .Y(\u_cpu._0218_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0746_  (.A(\u_cpu.led[5] ),
    .B(\u_cpu.led[4] ),
    .X(\u_cpu._0219_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu._0747_  (.A1(\u_cpu._0217_ ),
    .A2(\u_cpu.led[1] ),
    .B1(\u_cpu._0218_ ),
    .B2(\u_cpu._0219_ ),
    .Y(\u_cpu._0220_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0748_  (.A(\u_cpu.led[2] ),
    .B_N(\u_cpu.led[3] ),
    .X(\u_cpu._0221_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0749_  (.A(\u_cpu.led[3] ),
    .B_N(\u_cpu.led[2] ),
    .X(\u_cpu._0222_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu._0750_  (.A_N(\u_cpu.led[6] ),
    .B(\u_cpu.led[7] ),
    .X(\u_cpu._0223_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu._0751_  (.A_N(\u_cpu.led[7] ),
    .B(\u_cpu.led[6] ),
    .X(\u_cpu._0224_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu._0752_  (.A1_N(\u_cpu._0221_ ),
    .A2_N(\u_cpu._0222_ ),
    .B1(\u_cpu._0223_ ),
    .B2(\u_cpu._0224_ ),
    .Y(\u_cpu._0225_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0753_  (.A(\u_cpu.led[6] ),
    .B_N(\u_cpu.led[7] ),
    .X(\u_cpu._0226_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0754_  (.A(\u_cpu.led[7] ),
    .B_N(\u_cpu.led[6] ),
    .X(\u_cpu._0227_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._0755_  (.A(\u_cpu._0221_ ),
    .B(\u_cpu._0222_ ),
    .C(\u_cpu._0226_ ),
    .D(\u_cpu._0227_ ),
    .Y(\u_cpu._0228_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0756_  (.A(\u_cpu.led[1] ),
    .B(\u_cpu.ALUResult_W_Reg[0] ),
    .Y(\u_cpu._0229_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0757_  (.A(\u_cpu.led[1] ),
    .B(\u_cpu.ALUResult_W_Reg[0] ),
    .Y(\u_cpu._0230_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0758_  (.A(\u_cpu.led[5] ),
    .B(\u_cpu.led[4] ),
    .Y(\u_cpu._0231_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0759_  (.A(\u_cpu.led[5] ),
    .B(\u_cpu.led[4] ),
    .X(\u_cpu._0232_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu._0760_  (.A_N(\u_cpu._0229_ ),
    .B(\u_cpu._0230_ ),
    .C(\u_cpu._0231_ ),
    .D(\u_cpu._0232_ ),
    .Y(\u_cpu._0233_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu._0761_  (.A1(\u_cpu._0216_ ),
    .A2(\u_cpu._0220_ ),
    .B1(\u_cpu._0225_ ),
    .C1(\u_cpu._0228_ ),
    .D1(\u_cpu._0233_ ),
    .Y(\u_cpu._0234_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0762_  (.A(\u_cpu.led[1] ),
    .B(\u_cpu.ALUResult_W_Reg[0] ),
    .X(\u_cpu._0235_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu._0763_  (.A1(\u_cpu._0229_ ),
    .A2(\u_cpu._0235_ ),
    .B1(\u_cpu._0219_ ),
    .B2(\u_cpu._0218_ ),
    .Y(\u_cpu._0236_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu._0764_  (.A1(\u_cpu._0233_ ),
    .A2(\u_cpu._0236_ ),
    .B1(\u_cpu._0225_ ),
    .B2(\u_cpu._0228_ ),
    .X(\u_cpu._0237_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu._0765_  (.A1(\u_cpu._0214_ ),
    .A2(\u_cpu._0215_ ),
    .B1(\u_cpu._0234_ ),
    .C1(\u_cpu._0237_ ),
    .Y(\u_cpu._0238_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu._0766_  (.A1(\u_cpu._0216_ ),
    .A2(\u_cpu._0220_ ),
    .B1(\u_cpu._0225_ ),
    .C1(\u_cpu._0228_ ),
    .D1(\u_cpu._0233_ ),
    .X(\u_cpu._0239_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu._0767_  (.A1(\u_cpu._0233_ ),
    .A2(\u_cpu._0236_ ),
    .B1(\u_cpu._0225_ ),
    .B2(\u_cpu._0228_ ),
    .Y(\u_cpu._0240_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0768_  (.A(\u_cpu._0214_ ),
    .B(\u_cpu._0215_ ),
    .Y(\u_cpu._0241_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu._0769_  (.A1(\u_cpu._0239_ ),
    .A2(\u_cpu._0240_ ),
    .B1(\u_cpu._0241_ ),
    .Y(\u_cpu._0242_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0770_  (.A(\u_cpu.ALUResult_W_Reg[15] ),
    .B(\u_cpu.ALUResult_W_Reg[14] ),
    .X(\u_cpu._0243_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0771_  (.A(\u_cpu.ALUResult_W_Reg[15] ),
    .B(\u_cpu.ALUResult_W_Reg[14] ),
    .Y(\u_cpu._0244_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0772_  (.A(\u_cpu.ALUResult_W_Reg[11] ),
    .B(\u_cpu.ALUResult_W_Reg[10] ),
    .Y(\u_cpu._0245_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0773_  (.A(\u_cpu.ALUResult_W_Reg[11] ),
    .B(\u_cpu.ALUResult_W_Reg[10] ),
    .X(\u_cpu._0246_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu._0774_  (.A1(\u_cpu._0243_ ),
    .A2(\u_cpu._0244_ ),
    .B1(\u_cpu._0245_ ),
    .C1(\u_cpu._0246_ ),
    .X(\u_cpu._0247_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu._0775_  (.A(\u_cpu._0247_ ),
    .Y(\u_cpu._0248_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu._0776_  (.A1(\u_cpu._0245_ ),
    .A2(\u_cpu._0246_ ),
    .B1(\u_cpu._0243_ ),
    .C1(\u_cpu._0244_ ),
    .Y(\u_cpu._0249_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu._0777_  (.A(\u_cpu._0249_ ),
    .Y(\u_cpu._0250_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu._0778_  (.A1(\u_cpu._0238_ ),
    .A2(\u_cpu._0242_ ),
    .B1(\u_cpu._0248_ ),
    .C1(\u_cpu._0250_ ),
    .X(\u_cpu._0251_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu._0779_  (.A1(\u_cpu._0248_ ),
    .A2(\u_cpu._0250_ ),
    .B1(\u_cpu._0238_ ),
    .C1(\u_cpu._0242_ ),
    .Y(\u_cpu._0252_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu._0780_  (.A(\u_cpu._0209_ ),
    .B(\u_cpu._0251_ ),
    .C(\u_cpu._0252_ ),
    .Y(\u_cpu._0253_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu._0781_  (.A1(\u_cpu._0248_ ),
    .A2(\u_cpu._0250_ ),
    .B1(\u_cpu._0238_ ),
    .C1(\u_cpu._0242_ ),
    .X(\u_cpu._0254_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0782_  (.A(\u_cpu._0247_ ),
    .B(\u_cpu._0249_ ),
    .Y(\u_cpu._0255_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu._0783_  (.A1(\u_cpu._0238_ ),
    .A2(\u_cpu._0242_ ),
    .B1(\u_cpu._0255_ ),
    .Y(\u_cpu._0256_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu._0784_  (.A1(\u_cpu._0206_ ),
    .A2(\u_cpu._0198_ ),
    .B1(\u_cpu._0254_ ),
    .B2(\u_cpu._0256_ ),
    .C1(\u_cpu._0208_ ),
    .Y(\u_cpu._0257_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu._0785_  (.A(\u_cpu.M_AXI_WDATA[14] ),
    .Y(\u_cpu._0258_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0786_  (.A(\u_cpu._0258_ ),
    .B(\u_cpu.M_AXI_WDATA[15] ),
    .X(\u_cpu._0259_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0787_  (.A(\u_cpu.M_AXI_WDATA[13] ),
    .B(\u_cpu.M_AXI_WDATA[12] ),
    .Y(\u_cpu._0260_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0788_  (.A(\u_cpu.M_AXI_WDATA[13] ),
    .B(\u_cpu.M_AXI_WDATA[12] ),
    .X(\u_cpu._0261_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu._0789_  (.A1(\u_cpu.M_AXI_WDATA[15] ),
    .A2(\u_cpu._0258_ ),
    .B1(\u_cpu._0260_ ),
    .B2(\u_cpu._0261_ ),
    .Y(\u_cpu._0262_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0790_  (.A(\u_cpu.M_AXI_WDATA[9] ),
    .B(\u_cpu.M_AXI_WDATA[8] ),
    .Y(\u_cpu._0263_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0791_  (.A(\u_cpu.M_AXI_WDATA[9] ),
    .B(\u_cpu.M_AXI_WDATA[8] ),
    .X(\u_cpu._0264_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0792_  (.A(\u_cpu.M_AXI_WDATA[11] ),
    .B(\u_cpu.M_AXI_WDATA[10] ),
    .Y(\u_cpu._0265_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0793_  (.A(\u_cpu.M_AXI_WDATA[11] ),
    .B(\u_cpu.M_AXI_WDATA[10] ),
    .X(\u_cpu._0266_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu._0794_  (.A1(\u_cpu._0263_ ),
    .A2(\u_cpu._0264_ ),
    .B1(\u_cpu._0265_ ),
    .B2(\u_cpu._0266_ ),
    .X(\u_cpu._0267_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0795_  (.A(\u_cpu.M_AXI_WDATA[9] ),
    .B_N(\u_cpu.M_AXI_WDATA[8] ),
    .X(\u_cpu._0268_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0796_  (.A(\u_cpu.M_AXI_WDATA[8] ),
    .B_N(\u_cpu.M_AXI_WDATA[9] ),
    .X(\u_cpu._0269_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0797_  (.A(\u_cpu.M_AXI_WDATA[11] ),
    .B_N(\u_cpu.M_AXI_WDATA[10] ),
    .X(\u_cpu._0270_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0798_  (.A(\u_cpu.M_AXI_WDATA[10] ),
    .B_N(\u_cpu.M_AXI_WDATA[11] ),
    .X(\u_cpu._0271_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu._0799_  (.A1(\u_cpu._0268_ ),
    .A2(\u_cpu._0269_ ),
    .B1(\u_cpu._0270_ ),
    .B2(\u_cpu._0271_ ),
    .Y(\u_cpu._0272_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0800_  (.A(\u_cpu.M_AXI_WDATA[13] ),
    .B(\u_cpu.M_AXI_WDATA[12] ),
    .Y(\u_cpu._0273_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0801_  (.A(\u_cpu.M_AXI_WDATA[15] ),
    .B(\u_cpu.M_AXI_WDATA[14] ),
    .X(\u_cpu._0274_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0802_  (.A(\u_cpu.M_AXI_WDATA[15] ),
    .B(\u_cpu.M_AXI_WDATA[14] ),
    .Y(\u_cpu._0275_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu._0803_  (.A_N(\u_cpu._0260_ ),
    .B(\u_cpu._0273_ ),
    .C(\u_cpu._0274_ ),
    .D(\u_cpu._0275_ ),
    .Y(\u_cpu._0276_ ));
 sky130_fd_sc_hd__o221ai_2 \u_cpu._0804_  (.A1(\u_cpu._0259_ ),
    .A2(\u_cpu._0262_ ),
    .B1(\u_cpu._0267_ ),
    .B2(\u_cpu._0272_ ),
    .C1(\u_cpu._0276_ ),
    .Y(\u_cpu._0277_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu._0805_  (.A1(\u_cpu._0259_ ),
    .A2(\u_cpu._0262_ ),
    .B1(\u_cpu._0276_ ),
    .Y(\u_cpu._0278_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._0806_  (.A(\u_cpu._0268_ ),
    .B(\u_cpu._0269_ ),
    .C(\u_cpu._0270_ ),
    .D(\u_cpu._0271_ ),
    .Y(\u_cpu._0279_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu._0807_  (.A1(\u_cpu._0268_ ),
    .A2(\u_cpu._0269_ ),
    .B1(\u_cpu._0270_ ),
    .B2(\u_cpu._0271_ ),
    .X(\u_cpu._0280_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu._0808_  (.A(\u_cpu._0278_ ),
    .B(\u_cpu._0279_ ),
    .C(\u_cpu._0280_ ),
    .Y(\u_cpu._0281_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0809_  (.A(\u_cpu.M_AXI_WDATA[3] ),
    .B(\u_cpu.M_AXI_WDATA[2] ),
    .Y(\u_cpu._0282_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0810_  (.A(\u_cpu.M_AXI_WDATA[3] ),
    .B(\u_cpu.M_AXI_WDATA[2] ),
    .X(\u_cpu._0283_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0811_  (.A(\u_cpu.M_AXI_WDATA[1] ),
    .B(\u_cpu.M_AXI_WDATA[0] ),
    .Y(\u_cpu._0284_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0812_  (.A(\u_cpu.M_AXI_WDATA[1] ),
    .B(\u_cpu.M_AXI_WDATA[0] ),
    .X(\u_cpu._0285_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu._0813_  (.A1(\u_cpu._0282_ ),
    .A2(\u_cpu._0283_ ),
    .B1(\u_cpu._0284_ ),
    .B2(\u_cpu._0285_ ),
    .Y(\u_cpu._0286_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0814_  (.A(\u_cpu.M_AXI_WDATA[3] ),
    .B(\u_cpu.M_AXI_WDATA[2] ),
    .Y(\u_cpu._0287_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0815_  (.A(\u_cpu.M_AXI_WDATA[1] ),
    .B(\u_cpu.M_AXI_WDATA[0] ),
    .X(\u_cpu._0288_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0816_  (.A(\u_cpu.M_AXI_WDATA[1] ),
    .B(\u_cpu.M_AXI_WDATA[0] ),
    .Y(\u_cpu._0289_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu._0817_  (.A_N(\u_cpu._0282_ ),
    .B(\u_cpu._0287_ ),
    .C(\u_cpu._0288_ ),
    .D(\u_cpu._0289_ ),
    .Y(\u_cpu._0290_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0818_  (.A(\u_cpu.M_AXI_WDATA[7] ),
    .B(\u_cpu.M_AXI_WDATA[6] ),
    .X(\u_cpu._0291_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0819_  (.A(\u_cpu.M_AXI_WDATA[7] ),
    .B(\u_cpu.M_AXI_WDATA[6] ),
    .X(\u_cpu._0292_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0820_  (.A(\u_cpu.M_AXI_WDATA[5] ),
    .B(\u_cpu.M_AXI_WDATA[4] ),
    .Y(\u_cpu._0293_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0821_  (.A(\u_cpu.M_AXI_WDATA[5] ),
    .B(\u_cpu.M_AXI_WDATA[4] ),
    .X(\u_cpu._0294_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu._0822_  (.A_N(\u_cpu._0291_ ),
    .B(\u_cpu._0292_ ),
    .C(\u_cpu._0293_ ),
    .D(\u_cpu._0294_ ),
    .Y(\u_cpu._0295_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0823_  (.A(\u_cpu.M_AXI_WDATA[7] ),
    .B(\u_cpu.M_AXI_WDATA[6] ),
    .Y(\u_cpu._0296_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0824_  (.A(\u_cpu.M_AXI_WDATA[5] ),
    .B(\u_cpu.M_AXI_WDATA[4] ),
    .X(\u_cpu._0297_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0825_  (.A(\u_cpu.M_AXI_WDATA[5] ),
    .B(\u_cpu.M_AXI_WDATA[4] ),
    .Y(\u_cpu._0298_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu._0826_  (.A1(\u_cpu._0291_ ),
    .A2(\u_cpu._0296_ ),
    .B1(\u_cpu._0297_ ),
    .B2(\u_cpu._0298_ ),
    .Y(\u_cpu._0299_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu._0827_  (.A1(\u_cpu._0286_ ),
    .A2(\u_cpu._0290_ ),
    .B1(\u_cpu._0295_ ),
    .B2(\u_cpu._0299_ ),
    .X(\u_cpu._0300_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._0828_  (.A(\u_cpu._0286_ ),
    .B(\u_cpu._0290_ ),
    .C(\u_cpu._0295_ ),
    .D(\u_cpu._0299_ ),
    .Y(\u_cpu._0301_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._0829_  (.A(\u_cpu._0277_ ),
    .B(\u_cpu._0281_ ),
    .C(\u_cpu._0300_ ),
    .D(\u_cpu._0301_ ),
    .Y(\u_cpu._0302_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu._0830_  (.A1(\u_cpu._0286_ ),
    .A2(\u_cpu._0290_ ),
    .B1(\u_cpu._0295_ ),
    .B2(\u_cpu._0299_ ),
    .Y(\u_cpu._0303_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu._0831_  (.A(\u_cpu._0286_ ),
    .B(\u_cpu._0290_ ),
    .C(\u_cpu._0295_ ),
    .D(\u_cpu._0299_ ),
    .X(\u_cpu._0304_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu._0832_  (.A1_N(\u_cpu._0277_ ),
    .A2_N(\u_cpu._0281_ ),
    .B1(\u_cpu._0303_ ),
    .B2(\u_cpu._0304_ ),
    .Y(\u_cpu._0305_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0833_  (.A(\u_cpu._0302_ ),
    .B(\u_cpu._0305_ ),
    .Y(\u_cpu._0306_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0834_  (.A(\u_cpu.M_AXI_WDATA[25] ),
    .B_N(\u_cpu.M_AXI_WDATA[24] ),
    .X(\u_cpu._0307_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0835_  (.A(\u_cpu.M_AXI_WDATA[24] ),
    .B_N(\u_cpu.M_AXI_WDATA[25] ),
    .X(\u_cpu._0308_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0836_  (.A(\u_cpu.M_AXI_WDATA[27] ),
    .B_N(\u_cpu.M_AXI_WDATA[26] ),
    .X(\u_cpu._0309_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0837_  (.A(\u_cpu.M_AXI_WDATA[26] ),
    .B_N(\u_cpu.M_AXI_WDATA[27] ),
    .X(\u_cpu._0310_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._0838_  (.A(\u_cpu._0307_ ),
    .B(\u_cpu._0308_ ),
    .C(\u_cpu._0309_ ),
    .D(\u_cpu._0310_ ),
    .Y(\u_cpu._0311_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu._0839_  (.A_N(\u_cpu.M_AXI_WDATA[27] ),
    .B(\u_cpu.M_AXI_WDATA[26] ),
    .X(\u_cpu._0312_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu._0840_  (.A_N(\u_cpu.M_AXI_WDATA[26] ),
    .B(\u_cpu.M_AXI_WDATA[27] ),
    .X(\u_cpu._0313_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu._0841_  (.A1_N(\u_cpu._0307_ ),
    .A2_N(\u_cpu._0308_ ),
    .B1(\u_cpu._0312_ ),
    .B2(\u_cpu._0313_ ),
    .Y(\u_cpu._0314_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0842_  (.A(\u_cpu.M_AXI_WDATA[29] ),
    .B_N(\u_cpu.M_AXI_WDATA[28] ),
    .X(\u_cpu._0315_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0843_  (.A(\u_cpu.M_AXI_WDATA[28] ),
    .B_N(\u_cpu.M_AXI_WDATA[29] ),
    .X(\u_cpu._0316_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu._0844_  (.A_N(\u_cpu.M_AXI_WDATA[31] ),
    .B(\u_cpu.M_AXI_WDATA[30] ),
    .X(\u_cpu._0317_ ));
 sky130_fd_sc_hd__and2b_2 \u_cpu._0845_  (.A_N(\u_cpu.M_AXI_WDATA[30] ),
    .B(\u_cpu.M_AXI_WDATA[31] ),
    .X(\u_cpu._0318_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu._0846_  (.A1_N(\u_cpu._0315_ ),
    .A2_N(\u_cpu._0316_ ),
    .B1(\u_cpu._0317_ ),
    .B2(\u_cpu._0318_ ),
    .Y(\u_cpu._0319_ ));
 sky130_fd_sc_hd__a21boi_2 \u_cpu._0847_  (.A1(\u_cpu._0311_ ),
    .A2(\u_cpu._0314_ ),
    .B1_N(\u_cpu._0319_ ),
    .Y(\u_cpu._0320_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0848_  (.A(\u_cpu.M_AXI_WDATA[31] ),
    .B(\u_cpu.M_AXI_WDATA[30] ),
    .Y(\u_cpu._0321_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0849_  (.A(\u_cpu.M_AXI_WDATA[31] ),
    .B(\u_cpu.M_AXI_WDATA[30] ),
    .X(\u_cpu._0322_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu._0850_  (.A1(\u_cpu._0321_ ),
    .A2(\u_cpu._0322_ ),
    .B1(\u_cpu._0315_ ),
    .C1(\u_cpu._0316_ ),
    .Y(\u_cpu._0323_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0851_  (.A(\u_cpu.M_AXI_WDATA[17] ),
    .B(\u_cpu.M_AXI_WDATA[16] ),
    .Y(\u_cpu._0324_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0852_  (.A(\u_cpu.M_AXI_WDATA[17] ),
    .B(\u_cpu.M_AXI_WDATA[16] ),
    .X(\u_cpu._0325_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0853_  (.A(\u_cpu.M_AXI_WDATA[19] ),
    .B(\u_cpu.M_AXI_WDATA[18] ),
    .X(\u_cpu._0326_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0854_  (.A(\u_cpu.M_AXI_WDATA[19] ),
    .B(\u_cpu.M_AXI_WDATA[18] ),
    .Y(\u_cpu._0327_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu._0855_  (.A1(\u_cpu._0324_ ),
    .A2(\u_cpu._0325_ ),
    .B1(\u_cpu._0326_ ),
    .C1(\u_cpu._0327_ ),
    .Y(\u_cpu._0328_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0856_  (.A(\u_cpu.M_AXI_WDATA[17] ),
    .B(\u_cpu.M_AXI_WDATA[16] ),
    .Y(\u_cpu._0329_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0857_  (.A(\u_cpu.M_AXI_WDATA[18] ),
    .B_N(\u_cpu.M_AXI_WDATA[19] ),
    .X(\u_cpu._0330_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0858_  (.A(\u_cpu.M_AXI_WDATA[19] ),
    .B_N(\u_cpu.M_AXI_WDATA[18] ),
    .X(\u_cpu._0331_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu._0859_  (.A_N(\u_cpu._0324_ ),
    .B(\u_cpu._0329_ ),
    .C(\u_cpu._0330_ ),
    .D(\u_cpu._0331_ ),
    .Y(\u_cpu._0332_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0860_  (.A(\u_cpu.M_AXI_WDATA[21] ),
    .B(\u_cpu.M_AXI_WDATA[20] ),
    .X(\u_cpu._0333_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0861_  (.A(\u_cpu.M_AXI_WDATA[21] ),
    .B(\u_cpu.M_AXI_WDATA[20] ),
    .Y(\u_cpu._0334_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0862_  (.A(\u_cpu.M_AXI_WDATA[23] ),
    .B(\u_cpu.M_AXI_WDATA[22] ),
    .X(\u_cpu._0335_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0863_  (.A(\u_cpu.M_AXI_WDATA[23] ),
    .B(\u_cpu.M_AXI_WDATA[22] ),
    .Y(\u_cpu._0336_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \u_cpu._0864_  (.A1_N(\u_cpu._0333_ ),
    .A2_N(\u_cpu._0334_ ),
    .B1(\u_cpu._0335_ ),
    .B2(\u_cpu._0336_ ),
    .Y(\u_cpu._0337_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0865_  (.A(\u_cpu.M_AXI_WDATA[20] ),
    .B_N(\u_cpu.M_AXI_WDATA[21] ),
    .X(\u_cpu._0338_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0866_  (.A(\u_cpu.M_AXI_WDATA[21] ),
    .B_N(\u_cpu.M_AXI_WDATA[20] ),
    .X(\u_cpu._0339_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0867_  (.A(\u_cpu.M_AXI_WDATA[22] ),
    .B_N(\u_cpu.M_AXI_WDATA[23] ),
    .X(\u_cpu._0340_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0868_  (.A(\u_cpu.M_AXI_WDATA[23] ),
    .B_N(\u_cpu.M_AXI_WDATA[22] ),
    .X(\u_cpu._0341_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu._0869_  (.A1(\u_cpu._0338_ ),
    .A2(\u_cpu._0339_ ),
    .B1(\u_cpu._0340_ ),
    .B2(\u_cpu._0341_ ),
    .Y(\u_cpu._0342_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu._0870_  (.A1_N(\u_cpu._0328_ ),
    .A2_N(\u_cpu._0332_ ),
    .B1(\u_cpu._0337_ ),
    .B2(\u_cpu._0342_ ),
    .Y(\u_cpu._0343_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._0871_  (.A(\u_cpu._0338_ ),
    .B(\u_cpu._0339_ ),
    .C(\u_cpu._0340_ ),
    .D(\u_cpu._0341_ ),
    .Y(\u_cpu._0344_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0872_  (.A(\u_cpu.M_AXI_WDATA[21] ),
    .B(\u_cpu.M_AXI_WDATA[20] ),
    .X(\u_cpu._0345_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu._0873_  (.A_N(\u_cpu._0333_ ),
    .B(\u_cpu._0345_ ),
    .C(\u_cpu._0335_ ),
    .D(\u_cpu._0336_ ),
    .Y(\u_cpu._0346_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._0874_  (.A(\u_cpu._0328_ ),
    .B(\u_cpu._0332_ ),
    .C(\u_cpu._0344_ ),
    .D(\u_cpu._0346_ ),
    .Y(\u_cpu._0347_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0875_  (.A(\u_cpu.M_AXI_WDATA[25] ),
    .B(\u_cpu.M_AXI_WDATA[24] ),
    .Y(\u_cpu._0348_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0876_  (.A(\u_cpu.M_AXI_WDATA[25] ),
    .B(\u_cpu.M_AXI_WDATA[24] ),
    .X(\u_cpu._0349_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0877_  (.A(\u_cpu.M_AXI_WDATA[27] ),
    .B(\u_cpu.M_AXI_WDATA[26] ),
    .Y(\u_cpu._0350_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0878_  (.A(\u_cpu.M_AXI_WDATA[27] ),
    .B(\u_cpu.M_AXI_WDATA[26] ),
    .X(\u_cpu._0351_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu._0879_  (.A1(\u_cpu._0348_ ),
    .A2(\u_cpu._0349_ ),
    .B1(\u_cpu._0350_ ),
    .B2(\u_cpu._0351_ ),
    .X(\u_cpu._0352_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu._0880_  (.A1(\u_cpu._0307_ ),
    .A2(\u_cpu._0308_ ),
    .B1(\u_cpu._0309_ ),
    .B2(\u_cpu._0310_ ),
    .Y(\u_cpu._0353_ ));
 sky130_fd_sc_hd__a211oi_2 \u_cpu._0881_  (.A1(\u_cpu._0323_ ),
    .A2(\u_cpu._0319_ ),
    .B1(\u_cpu._0352_ ),
    .C1(\u_cpu._0353_ ),
    .Y(\u_cpu._0354_ ));
 sky130_fd_sc_hd__a221o_2 \u_cpu._0882_  (.A1(\u_cpu._0320_ ),
    .A2(\u_cpu._0323_ ),
    .B1(\u_cpu._0343_ ),
    .B2(\u_cpu._0347_ ),
    .C1(\u_cpu._0354_ ),
    .X(\u_cpu._0355_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0883_  (.A(\u_cpu._0320_ ),
    .B(\u_cpu._0323_ ),
    .Y(\u_cpu._0356_ ));
 sky130_fd_sc_hd__a211o_2 \u_cpu._0884_  (.A1(\u_cpu._0323_ ),
    .A2(\u_cpu._0319_ ),
    .B1(\u_cpu._0352_ ),
    .C1(\u_cpu._0353_ ),
    .X(\u_cpu._0357_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu._0885_  (.A(\u_cpu._0328_ ),
    .B(\u_cpu._0332_ ),
    .C(\u_cpu._0346_ ),
    .Y(\u_cpu._0358_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu._0886_  (.A1(\u_cpu._0337_ ),
    .A2(\u_cpu._0358_ ),
    .B1(\u_cpu._0343_ ),
    .Y(\u_cpu._0359_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu._0887_  (.A1(\u_cpu._0356_ ),
    .A2(\u_cpu._0357_ ),
    .B1(\u_cpu._0359_ ),
    .X(\u_cpu._0360_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu._0888_  (.A(\u_cpu._0306_ ),
    .B(\u_cpu._0355_ ),
    .C(\u_cpu._0360_ ),
    .Y(\u_cpu._0361_ ));
 sky130_fd_sc_hd__a221oi_2 \u_cpu._0889_  (.A1(\u_cpu._0320_ ),
    .A2(\u_cpu._0323_ ),
    .B1(\u_cpu._0343_ ),
    .B2(\u_cpu._0347_ ),
    .C1(\u_cpu._0354_ ),
    .Y(\u_cpu._0362_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu._0890_  (.A1(\u_cpu._0356_ ),
    .A2(\u_cpu._0357_ ),
    .B1(\u_cpu._0359_ ),
    .Y(\u_cpu._0363_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu._0891_  (.A1(\u_cpu._0362_ ),
    .A2(\u_cpu._0363_ ),
    .B1(\u_cpu._0302_ ),
    .C1(\u_cpu._0305_ ),
    .Y(\u_cpu._0364_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0892_  (.A(\u_cpu.IMEM.a[3] ),
    .B(\u_cpu.IMEM.a[2] ),
    .Y(\u_cpu._0365_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0893_  (.A(\u_cpu.IMEM.a[3] ),
    .B(\u_cpu.IMEM.a[2] ),
    .X(\u_cpu._0366_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0894_  (.A(\u_cpu.IMEM.a[5] ),
    .B(\u_cpu.IMEM.a[4] ),
    .Y(\u_cpu._0367_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0895_  (.A(\u_cpu.IMEM.a[5] ),
    .B(\u_cpu.IMEM.a[4] ),
    .X(\u_cpu._0368_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu._0896_  (.A1(\u_cpu._0365_ ),
    .A2(\u_cpu._0366_ ),
    .B1(\u_cpu._0367_ ),
    .C1(\u_cpu._0368_ ),
    .Y(\u_cpu._0369_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0897_  (.A(\u_cpu.IMEM.a[5] ),
    .B(\u_cpu.IMEM.a[4] ),
    .X(\u_cpu._0370_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0898_  (.A(\u_cpu.IMEM.a[5] ),
    .B(\u_cpu.IMEM.a[4] ),
    .Y(\u_cpu._0371_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0899_  (.A(\u_cpu.IMEM.a[3] ),
    .B(\u_cpu.IMEM.a[2] ),
    .X(\u_cpu._0372_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0900_  (.A(\u_cpu.IMEM.a[3] ),
    .B(\u_cpu.IMEM.a[2] ),
    .Y(\u_cpu._0373_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu._0901_  (.A1(\u_cpu._0370_ ),
    .A2(\u_cpu._0371_ ),
    .B1(\u_cpu._0372_ ),
    .C1(\u_cpu._0373_ ),
    .Y(\u_cpu._0374_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0902_  (.A(\u_cpu.IMEM.a[7] ),
    .B(\u_cpu.IMEM.a[6] ),
    .X(\u_cpu._0375_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0903_  (.A(\u_cpu.IMEM.a[7] ),
    .B(\u_cpu.IMEM.a[6] ),
    .Y(\u_cpu._0376_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0904_  (.A(\u_cpu._0375_ ),
    .B(\u_cpu._0376_ ),
    .Y(\u_cpu._0377_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu._0905_  (.A1(\u_cpu._0369_ ),
    .A2(\u_cpu._0374_ ),
    .B1(\u_cpu._0377_ ),
    .X(\u_cpu._0378_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu._0906_  (.A1(\u_cpu._0365_ ),
    .A2(\u_cpu._0366_ ),
    .B1(\u_cpu._0368_ ),
    .Y(\u_cpu._0379_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu._0907_  (.A1(\u_cpu._0370_ ),
    .A2(\u_cpu._0379_ ),
    .B1(\u_cpu._0374_ ),
    .C1(\u_cpu._0377_ ),
    .Y(\u_cpu._0380_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0908_  (.A(\u_cpu.IMEM.a[15] ),
    .B(\u_cpu.IMEM.a[14] ),
    .Y(\u_cpu._0381_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0909_  (.A(\u_cpu.IMEM.a[15] ),
    .B(\u_cpu.IMEM.a[14] ),
    .X(\u_cpu._0382_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0910_  (.A(\u_cpu.IMEM.a[9] ),
    .B(\u_cpu.IMEM.a[8] ),
    .Y(\u_cpu._0383_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0911_  (.A(\u_cpu.IMEM.a[9] ),
    .B(\u_cpu.IMEM.a[8] ),
    .X(\u_cpu._0384_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu._0912_  (.A1(\u_cpu._0381_ ),
    .A2(\u_cpu._0382_ ),
    .B1(\u_cpu._0383_ ),
    .C1(\u_cpu._0384_ ),
    .Y(\u_cpu._0385_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0913_  (.A(\u_cpu.IMEM.a[9] ),
    .B(\u_cpu.IMEM.a[8] ),
    .X(\u_cpu._0386_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0914_  (.A(\u_cpu.IMEM.a[9] ),
    .B(\u_cpu.IMEM.a[8] ),
    .Y(\u_cpu._0387_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0915_  (.A(\u_cpu.IMEM.a[15] ),
    .B(\u_cpu.IMEM.a[14] ),
    .X(\u_cpu._0388_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0916_  (.A(\u_cpu.IMEM.a[15] ),
    .B(\u_cpu.IMEM.a[14] ),
    .Y(\u_cpu._0389_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu._0917_  (.A1(\u_cpu._0386_ ),
    .A2(\u_cpu._0387_ ),
    .B1(\u_cpu._0388_ ),
    .C1(\u_cpu._0389_ ),
    .Y(\u_cpu._0390_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0918_  (.A(\u_cpu.IMEM.a[13] ),
    .B(\u_cpu.IMEM.a[12] ),
    .Y(\u_cpu._0391_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0919_  (.A(\u_cpu.IMEM.a[13] ),
    .B(\u_cpu.IMEM.a[12] ),
    .X(\u_cpu._0392_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0920_  (.A(\u_cpu.IMEM.a[11] ),
    .B(\u_cpu.IMEM.a[10] ),
    .Y(\u_cpu._0393_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0921_  (.A(\u_cpu.IMEM.a[11] ),
    .B(\u_cpu.IMEM.a[10] ),
    .X(\u_cpu._0394_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu._0922_  (.A1(\u_cpu._0391_ ),
    .A2(\u_cpu._0392_ ),
    .B1(\u_cpu._0393_ ),
    .B2(\u_cpu._0394_ ),
    .Y(\u_cpu._0395_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0923_  (.A(\u_cpu.IMEM.a[13] ),
    .B(\u_cpu.IMEM.a[12] ),
    .Y(\u_cpu._0396_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0924_  (.A(\u_cpu.IMEM.a[11] ),
    .B(\u_cpu.IMEM.a[10] ),
    .X(\u_cpu._0397_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0925_  (.A(\u_cpu.IMEM.a[11] ),
    .B(\u_cpu.IMEM.a[10] ),
    .Y(\u_cpu._0398_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu._0926_  (.A_N(\u_cpu._0391_ ),
    .B(\u_cpu._0396_ ),
    .C(\u_cpu._0397_ ),
    .D(\u_cpu._0398_ ),
    .Y(\u_cpu._0399_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._0927_  (.A(\u_cpu._0385_ ),
    .B(\u_cpu._0390_ ),
    .C(\u_cpu._0395_ ),
    .D(\u_cpu._0399_ ),
    .Y(\u_cpu._0400_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu._0928_  (.A(\u_cpu._0378_ ),
    .B(\u_cpu._0380_ ),
    .C(\u_cpu._0400_ ),
    .Y(\u_cpu._0401_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu._0929_  (.A1(\u_cpu._0385_ ),
    .A2(\u_cpu._0390_ ),
    .B1(\u_cpu._0395_ ),
    .B2(\u_cpu._0399_ ),
    .Y(\u_cpu._0402_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu._0930_  (.A1(\u_cpu._0369_ ),
    .A2(\u_cpu._0374_ ),
    .B1(\u_cpu._0377_ ),
    .Y(\u_cpu._0403_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu._0931_  (.A1(\u_cpu._0370_ ),
    .A2(\u_cpu._0379_ ),
    .B1(\u_cpu._0374_ ),
    .C1(\u_cpu._0377_ ),
    .X(\u_cpu._0404_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu._0932_  (.A(\u_cpu._0385_ ),
    .B(\u_cpu._0390_ ),
    .C(\u_cpu._0395_ ),
    .D(\u_cpu._0399_ ),
    .X(\u_cpu._0405_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu._0933_  (.A1(\u_cpu._0403_ ),
    .A2(\u_cpu._0404_ ),
    .B1(\u_cpu._0402_ ),
    .B2(\u_cpu._0405_ ),
    .Y(\u_cpu._0406_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0934_  (.A(\u_cpu.IMEM.a[17] ),
    .B(\u_cpu.IMEM.a[16] ),
    .X(\u_cpu._0407_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0935_  (.A(\u_cpu.IMEM.a[23] ),
    .B(\u_cpu.IMEM.a[22] ),
    .Y(\u_cpu._0408_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0936_  (.A(\u_cpu.IMEM.a[23] ),
    .B(\u_cpu.IMEM.a[22] ),
    .X(\u_cpu._0409_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0937_  (.A(\u_cpu.IMEM.a[17] ),
    .B(\u_cpu.IMEM.a[16] ),
    .X(\u_cpu._0410_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu._0938_  (.A1(\u_cpu._0408_ ),
    .A2(\u_cpu._0409_ ),
    .B1(\u_cpu._0410_ ),
    .Y(\u_cpu._0411_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0939_  (.A(\u_cpu.IMEM.a[17] ),
    .B(\u_cpu.IMEM.a[16] ),
    .Y(\u_cpu._0412_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0940_  (.A(\u_cpu._0408_ ),
    .B(\u_cpu._0409_ ),
    .Y(\u_cpu._0413_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu._0941_  (.A1(\u_cpu._0407_ ),
    .A2(\u_cpu._0412_ ),
    .B1(\u_cpu._0413_ ),
    .Y(\u_cpu._0414_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0942_  (.A(\u_cpu.IMEM.a[21] ),
    .B(\u_cpu.IMEM.a[20] ),
    .Y(\u_cpu._0415_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0943_  (.A(\u_cpu.IMEM.a[21] ),
    .B(\u_cpu.IMEM.a[20] ),
    .X(\u_cpu._0416_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0944_  (.A(\u_cpu.IMEM.a[19] ),
    .B(\u_cpu.IMEM.a[18] ),
    .X(\u_cpu._0417_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0945_  (.A(\u_cpu.IMEM.a[19] ),
    .B(\u_cpu.IMEM.a[18] ),
    .Y(\u_cpu._0418_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu._0946_  (.A1(\u_cpu._0415_ ),
    .A2(\u_cpu._0416_ ),
    .B1(\u_cpu._0417_ ),
    .B2(\u_cpu._0418_ ),
    .Y(\u_cpu._0419_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0947_  (.A(\u_cpu._0415_ ),
    .B(\u_cpu._0416_ ),
    .Y(\u_cpu._0420_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0948_  (.A(\u_cpu._0417_ ),
    .B(\u_cpu._0418_ ),
    .Y(\u_cpu._0421_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0949_  (.A(\u_cpu._0420_ ),
    .B(\u_cpu._0421_ ),
    .Y(\u_cpu._0422_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu._0950_  (.A1(\u_cpu._0407_ ),
    .A2(\u_cpu._0411_ ),
    .B1(\u_cpu._0414_ ),
    .C1(\u_cpu._0419_ ),
    .D1(\u_cpu._0422_ ),
    .Y(\u_cpu._0423_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu._0951_  (.A1(\u_cpu._0415_ ),
    .A2(\u_cpu._0416_ ),
    .B1(\u_cpu._0421_ ),
    .Y(\u_cpu._0424_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu._0952_  (.A1(\u_cpu._0417_ ),
    .A2(\u_cpu._0418_ ),
    .B1(\u_cpu._0420_ ),
    .Y(\u_cpu._0425_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu._0953_  (.A1(\u_cpu._0408_ ),
    .A2(\u_cpu._0409_ ),
    .B1(\u_cpu._0407_ ),
    .B2(\u_cpu._0412_ ),
    .Y(\u_cpu._0426_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0954_  (.A(\u_cpu.IMEM.a[23] ),
    .B(\u_cpu.IMEM.a[22] ),
    .Y(\u_cpu._0427_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0955_  (.A(\u_cpu.IMEM.a[17] ),
    .B(\u_cpu.IMEM.a[16] ),
    .Y(\u_cpu._0428_ ));
 sky130_fd_sc_hd__nand4b_2 \u_cpu._0956_  (.A_N(\u_cpu._0408_ ),
    .B(\u_cpu._0427_ ),
    .C(\u_cpu._0428_ ),
    .D(\u_cpu._0410_ ),
    .Y(\u_cpu._0429_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._0957_  (.A(\u_cpu._0424_ ),
    .B(\u_cpu._0425_ ),
    .C(\u_cpu._0426_ ),
    .D(\u_cpu._0429_ ),
    .Y(\u_cpu._0430_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0958_  (.A(\u_cpu._0423_ ),
    .B(\u_cpu._0430_ ),
    .Y(\u_cpu._0431_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0959_  (.A(\u_cpu.IMEM.a[25] ),
    .B(\u_cpu.IMEM.a[24] ),
    .X(\u_cpu._0432_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0960_  (.A(\u_cpu.IMEM.a[25] ),
    .B(\u_cpu.IMEM.a[24] ),
    .Y(\u_cpu._0433_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu._0961_  (.A(\u_cpu.IMEM.a[27] ),
    .B(\u_cpu.IMEM.a[26] ),
    .Y(\u_cpu._0434_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu._0962_  (.A1(\u_cpu._0432_ ),
    .A2(\u_cpu._0433_ ),
    .B1(\u_cpu._0434_ ),
    .Y(\u_cpu._0435_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0963_  (.A(\u_cpu.IMEM.a[27] ),
    .B_N(\u_cpu.IMEM.a[26] ),
    .X(\u_cpu._0436_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0964_  (.A(\u_cpu.IMEM.a[26] ),
    .B_N(\u_cpu.IMEM.a[27] ),
    .X(\u_cpu._0437_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0965_  (.A(\u_cpu.IMEM.a[25] ),
    .B_N(\u_cpu.IMEM.a[24] ),
    .X(\u_cpu._0438_ ));
 sky130_fd_sc_hd__or2b_2 \u_cpu._0966_  (.A(\u_cpu.IMEM.a[24] ),
    .B_N(\u_cpu.IMEM.a[25] ),
    .X(\u_cpu._0439_ ));
 sky130_fd_sc_hd__a22o_2 \u_cpu._0967_  (.A1(\u_cpu._0436_ ),
    .A2(\u_cpu._0437_ ),
    .B1(\u_cpu._0438_ ),
    .B2(\u_cpu._0439_ ),
    .X(\u_cpu._0440_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0968_  (.A(\u_cpu.IMEM.a[29] ),
    .B(\u_cpu.IMEM.a[28] ),
    .Y(\u_cpu._0441_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0969_  (.A(\u_cpu.IMEM.a[29] ),
    .B(\u_cpu.IMEM.a[28] ),
    .X(\u_cpu._0442_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._0970_  (.A(\u_cpu.IMEM.a[31] ),
    .B(\u_cpu.IMEM.a[30] ),
    .Y(\u_cpu._0443_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._0971_  (.A(\u_cpu.IMEM.a[31] ),
    .B(\u_cpu.IMEM.a[30] ),
    .X(\u_cpu._0444_ ));
 sky130_fd_sc_hd__o22ai_2 \u_cpu._0972_  (.A1(\u_cpu._0441_ ),
    .A2(\u_cpu._0442_ ),
    .B1(\u_cpu._0443_ ),
    .B2(\u_cpu._0444_ ),
    .Y(\u_cpu._0445_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0973_  (.A(\u_cpu.IMEM.a[29] ),
    .B(\u_cpu.IMEM.a[28] ),
    .X(\u_cpu._0446_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0974_  (.A(\u_cpu.IMEM.a[29] ),
    .B(\u_cpu.IMEM.a[28] ),
    .Y(\u_cpu._0447_ ));
 sky130_fd_sc_hd__or2_2 \u_cpu._0975_  (.A(\u_cpu.IMEM.a[31] ),
    .B(\u_cpu.IMEM.a[30] ),
    .X(\u_cpu._0448_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0976_  (.A(\u_cpu.IMEM.a[31] ),
    .B(\u_cpu.IMEM.a[30] ),
    .Y(\u_cpu._0449_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._0977_  (.A(\u_cpu._0446_ ),
    .B(\u_cpu._0447_ ),
    .C(\u_cpu._0448_ ),
    .D(\u_cpu._0449_ ),
    .Y(\u_cpu._0450_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._0978_  (.A(\u_cpu._0435_ ),
    .B(\u_cpu._0440_ ),
    .C(\u_cpu._0445_ ),
    .D(\u_cpu._0450_ ),
    .Y(\u_cpu._0451_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0979_  (.A(\u_cpu._0438_ ),
    .B(\u_cpu._0439_ ),
    .Y(\u_cpu._0452_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0980_  (.A(\u_cpu._0434_ ),
    .B(\u_cpu._0452_ ),
    .Y(\u_cpu._0453_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0981_  (.A(\u_cpu._0436_ ),
    .B(\u_cpu._0437_ ),
    .Y(\u_cpu._0454_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu._0982_  (.A1(\u_cpu._0432_ ),
    .A2(\u_cpu._0433_ ),
    .B1(\u_cpu._0454_ ),
    .Y(\u_cpu._0455_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu._0983_  (.A1(\u_cpu._0443_ ),
    .A2(\u_cpu._0444_ ),
    .B1(\u_cpu._0446_ ),
    .C1(\u_cpu._0447_ ),
    .Y(\u_cpu._0456_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu._0984_  (.A1(\u_cpu._0441_ ),
    .A2(\u_cpu._0442_ ),
    .B1(\u_cpu._0448_ ),
    .C1(\u_cpu._0449_ ),
    .Y(\u_cpu._0457_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._0985_  (.A(\u_cpu._0453_ ),
    .B(\u_cpu._0455_ ),
    .C(\u_cpu._0456_ ),
    .D(\u_cpu._0457_ ),
    .Y(\u_cpu._0458_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu._0986_  (.A(\u_cpu._0431_ ),
    .B(\u_cpu._0451_ ),
    .C(\u_cpu._0458_ ),
    .Y(\u_cpu._0459_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._0987_  (.A(\u_cpu._0451_ ),
    .B(\u_cpu._0458_ ),
    .Y(\u_cpu._0460_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu._0988_  (.A(\u_cpu._0423_ ),
    .B(\u_cpu._0430_ ),
    .C(\u_cpu._0460_ ),
    .Y(\u_cpu._0461_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu._0989_  (.A1(\u_cpu._0401_ ),
    .A2(\u_cpu._0402_ ),
    .B1(\u_cpu._0406_ ),
    .C1(\u_cpu._0459_ ),
    .D1(\u_cpu._0461_ ),
    .X(\u_cpu._0462_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu._0990_  (.A1(\u_cpu._0423_ ),
    .A2(\u_cpu._0430_ ),
    .B1(\u_cpu._0460_ ),
    .Y(\u_cpu._0463_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu._0991_  (.A1(\u_cpu._0451_ ),
    .A2(\u_cpu._0458_ ),
    .B1(\u_cpu._0431_ ),
    .Y(\u_cpu._0464_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu._0992_  (.A1(\u_cpu._0402_ ),
    .A2(\u_cpu._0401_ ),
    .B1(\u_cpu._0406_ ),
    .Y(\u_cpu._0465_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu._0993_  (.A1(\u_cpu._0463_ ),
    .A2(\u_cpu._0464_ ),
    .B1(\u_cpu._0465_ ),
    .X(\u_cpu._0466_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \u_cpu._0994_  (.A1_N(\u_cpu._0361_ ),
    .A2_N(\u_cpu._0364_ ),
    .B1(\u_cpu._0462_ ),
    .B2(\u_cpu._0466_ ),
    .Y(\u_cpu._0467_ ));
 sky130_fd_sc_hd__o2111ai_2 \u_cpu._0995_  (.A1(\u_cpu._0401_ ),
    .A2(\u_cpu._0402_ ),
    .B1(\u_cpu._0406_ ),
    .C1(\u_cpu._0459_ ),
    .D1(\u_cpu._0461_ ),
    .Y(\u_cpu._0468_ ));
 sky130_fd_sc_hd__o21ai_2 \u_cpu._0996_  (.A1(\u_cpu._0463_ ),
    .A2(\u_cpu._0464_ ),
    .B1(\u_cpu._0465_ ),
    .Y(\u_cpu._0469_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._0997_  (.A(\u_cpu._0361_ ),
    .B(\u_cpu._0364_ ),
    .C(\u_cpu._0468_ ),
    .D(\u_cpu._0469_ ),
    .Y(\u_cpu._0470_ ));
 sky130_fd_sc_hd__a22oi_2 \u_cpu._0998_  (.A1(\u_cpu._0253_ ),
    .A2(\u_cpu._0257_ ),
    .B1(\u_cpu._0467_ ),
    .B2(\u_cpu._0470_ ),
    .Y(\u_cpu._0471_ ));
 sky130_fd_sc_hd__o211ai_2 \u_cpu._0999_  (.A1(\u_cpu._0173_ ),
    .A2(\u_cpu._0174_ ),
    .B1(\u_cpu._0193_ ),
    .C1(\u_cpu._0197_ ),
    .Y(\u_cpu._0472_ ));
 sky130_fd_sc_hd__nand3_2 \u_cpu._1000_  (.A(\u_cpu._0202_ ),
    .B(\u_cpu._0472_ ),
    .C(\u_cpu._0205_ ),
    .Y(\u_cpu._0473_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu._1001_  (.A1(\u_cpu._0208_ ),
    .A2(\u_cpu._0473_ ),
    .B1(\u_cpu._0254_ ),
    .X(\u_cpu._0474_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu._1002_  (.A1(\u_cpu._0256_ ),
    .A2(\u_cpu._0474_ ),
    .B1(\u_cpu._0257_ ),
    .C1(\u_cpu._0467_ ),
    .D1(\u_cpu._0470_ ),
    .X(\u_cpu._0475_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._1003_  (.A(\u_cpu._0471_ ),
    .B(\u_cpu._0475_ ),
    .Y(\u_cpu.led[0] ));
 sky130_fd_sc_hd__xor2_2 \u_cpu._1004_  (.A(\u_cpu.counter[1] ),
    .B(\u_cpu.counter[0] ),
    .X(\u_cpu._0011_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1005_  (.A(\u_cpu.counter[1] ),
    .B(\u_cpu.counter[0] ),
    .C(\u_cpu.counter[2] ),
    .X(\u_cpu._0476_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu._1006_  (.A1(\u_cpu.counter[1] ),
    .A2(\u_cpu.counter[0] ),
    .B1(\u_cpu.counter[2] ),
    .Y(\u_cpu._0477_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._1007_  (.A(\u_cpu._0476_ ),
    .B(\u_cpu._0477_ ),
    .Y(\u_cpu._0018_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._1008_  (.A(\u_cpu.counter[1] ),
    .B(\u_cpu.counter[0] ),
    .C(\u_cpu.counter[3] ),
    .D(\u_cpu.counter[2] ),
    .Y(\u_cpu._0478_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu._1009_  (.A1(\u_cpu.counter[1] ),
    .A2(\u_cpu.counter[0] ),
    .A3(\u_cpu.counter[2] ),
    .B1(\u_cpu.counter[3] ),
    .X(\u_cpu._0479_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._1010_  (.A(\u_cpu._0478_ ),
    .B(\u_cpu._0479_ ),
    .X(\u_cpu._0480_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1011_  (.A(\u_cpu._0480_ ),
    .X(\u_cpu._0019_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu._1012_  (.A(\u_cpu.counter[4] ),
    .B(\u_cpu._0478_ ),
    .Y(\u_cpu._0020_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu._1013_  (.A(\u_cpu.counter[5] ),
    .Y(\u_cpu._0481_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu._1014_  (.A(\u_cpu.counter[4] ),
    .Y(\u_cpu._0482_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu._1015_  (.A(\u_cpu._0481_ ),
    .B(\u_cpu._0482_ ),
    .C(\u_cpu._0478_ ),
    .Y(\u_cpu._0483_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu._1016_  (.A1(\u_cpu._0482_ ),
    .A2(\u_cpu._0478_ ),
    .B1(\u_cpu._0481_ ),
    .X(\u_cpu._0484_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._1017_  (.A(\u_cpu._0483_ ),
    .B(\u_cpu._0484_ ),
    .Y(\u_cpu._0021_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu._1018_  (.A(\u_cpu.counter[6] ),
    .B(\u_cpu._0483_ ),
    .X(\u_cpu._0022_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1019_  (.A(\u_cpu.counter[7] ),
    .B(\u_cpu.counter[6] ),
    .C(\u_cpu._0483_ ),
    .X(\u_cpu._0485_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu._1020_  (.A1(\u_cpu.counter[6] ),
    .A2(\u_cpu._0483_ ),
    .B1(\u_cpu.counter[7] ),
    .Y(\u_cpu._0486_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._1021_  (.A(\u_cpu._0485_ ),
    .B(\u_cpu._0486_ ),
    .Y(\u_cpu._0023_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu._1022_  (.A(\u_cpu.counter[7] ),
    .B(\u_cpu.counter[6] ),
    .C(\u_cpu.counter[8] ),
    .D(\u_cpu._0483_ ),
    .X(\u_cpu._0487_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._1023_  (.A(\u_cpu.counter[8] ),
    .B(\u_cpu._0485_ ),
    .Y(\u_cpu._0488_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._1024_  (.A(\u_cpu._0487_ ),
    .B(\u_cpu._0488_ ),
    .Y(\u_cpu._0024_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1025_  (.A(\u_cpu.counter[9] ),
    .B(\u_cpu.counter[8] ),
    .C(\u_cpu._0485_ ),
    .X(\u_cpu._0489_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu._1026_  (.A1(\u_cpu.counter[9] ),
    .A2(\u_cpu._0487_ ),
    .B1_N(\u_cpu._0489_ ),
    .X(\u_cpu._0025_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu._1027_  (.A(\u_cpu.counter[10] ),
    .B(\u_cpu._0489_ ),
    .X(\u_cpu._0001_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu._1028_  (.A(\u_cpu.counter[9] ),
    .B(\u_cpu.counter[8] ),
    .C(\u_cpu.counter[11] ),
    .D(\u_cpu.counter[10] ),
    .X(\u_cpu._0490_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu._1029_  (.A1(\u_cpu.counter[10] ),
    .A2(\u_cpu._0489_ ),
    .B1(\u_cpu.counter[11] ),
    .Y(\u_cpu._0491_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu._1030_  (.A1(\u_cpu._0485_ ),
    .A2(\u_cpu._0490_ ),
    .B1(\u_cpu._0491_ ),
    .Y(\u_cpu._0002_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1031_  (.A(\u_cpu.counter[12] ),
    .B(\u_cpu._0485_ ),
    .C(\u_cpu._0490_ ),
    .X(\u_cpu._0492_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu._1032_  (.A1(\u_cpu._0485_ ),
    .A2(\u_cpu._0490_ ),
    .B1(\u_cpu.counter[12] ),
    .Y(\u_cpu._0493_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._1033_  (.A(\u_cpu._0492_ ),
    .B(\u_cpu._0493_ ),
    .Y(\u_cpu._0003_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._1034_  (.A(\u_cpu.counter[7] ),
    .B(\u_cpu.counter[6] ),
    .C(\u_cpu._0483_ ),
    .D(\u_cpu._0490_ ),
    .Y(\u_cpu._0494_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._1035_  (.A(\u_cpu.counter[13] ),
    .B(\u_cpu.counter[12] ),
    .Y(\u_cpu._0495_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu._1036_  (.A1(\u_cpu._0494_ ),
    .A2(\u_cpu._0495_ ),
    .B1(\u_cpu._0492_ ),
    .B2(\u_cpu.counter[13] ),
    .X(\u_cpu._0004_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1037_  (.A(\u_cpu.counter[11] ),
    .B(\u_cpu.counter[10] ),
    .C(\u_cpu._0489_ ),
    .X(\u_cpu._0496_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu._1038_  (.A(\u_cpu.counter[13] ),
    .B(\u_cpu.counter[12] ),
    .C(\u_cpu.counter[14] ),
    .D(\u_cpu._0496_ ),
    .X(\u_cpu._0497_ ));
 sky130_fd_sc_hd__a31oi_2 \u_cpu._1039_  (.A1(\u_cpu.counter[13] ),
    .A2(\u_cpu.counter[12] ),
    .A3(\u_cpu._0496_ ),
    .B1(\u_cpu.counter[14] ),
    .Y(\u_cpu._0498_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._1040_  (.A(\u_cpu._0497_ ),
    .B(\u_cpu._0498_ ),
    .Y(\u_cpu._0005_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._1041_  (.A(\u_cpu.counter[15] ),
    .B(\u_cpu.counter[14] ),
    .Y(\u_cpu._0499_ ));
 sky130_fd_sc_hd__o32a_2 \u_cpu._1042_  (.A1(\u_cpu._0494_ ),
    .A2(\u_cpu._0495_ ),
    .A3(\u_cpu._0499_ ),
    .B1(\u_cpu._0497_ ),
    .B2(\u_cpu.counter[15] ),
    .X(\u_cpu._0006_ ));
 sky130_fd_sc_hd__nor3_2 \u_cpu._1043_  (.A(\u_cpu._0494_ ),
    .B(\u_cpu._0495_ ),
    .C(\u_cpu._0499_ ),
    .Y(\u_cpu._0500_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu._1044_  (.A(\u_cpu.counter[16] ),
    .B(\u_cpu._0500_ ),
    .X(\u_cpu._0007_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._1045_  (.A(\u_cpu.counter[17] ),
    .B(\u_cpu.counter[16] ),
    .X(\u_cpu._0501_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu._1046_  (.A1(\u_cpu.counter[16] ),
    .A2(\u_cpu._0500_ ),
    .B1(\u_cpu.counter[17] ),
    .Y(\u_cpu._0502_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu._1047_  (.A1(\u_cpu._0500_ ),
    .A2(\u_cpu._0501_ ),
    .B1(\u_cpu._0502_ ),
    .Y(\u_cpu._0008_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1048_  (.A(\u_cpu.counter[18] ),
    .B(\u_cpu._0500_ ),
    .C(\u_cpu._0501_ ),
    .X(\u_cpu._0503_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu._1049_  (.A1(\u_cpu._0500_ ),
    .A2(\u_cpu._0501_ ),
    .B1(\u_cpu.counter[18] ),
    .Y(\u_cpu._0504_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._1050_  (.A(\u_cpu._0503_ ),
    .B(\u_cpu._0504_ ),
    .Y(\u_cpu._0009_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1051_  (.A(\u_cpu.counter[17] ),
    .B(\u_cpu.counter[16] ),
    .C(\u_cpu._0500_ ),
    .X(\u_cpu._0505_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._1052_  (.A(\u_cpu.counter[19] ),
    .B(\u_cpu.counter[18] ),
    .X(\u_cpu._0506_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1053_  (.A(\u_cpu._0506_ ),
    .X(\u_cpu._0507_ ));
 sky130_fd_sc_hd__o2bb2a_2 \u_cpu._1054_  (.A1_N(\u_cpu._0505_ ),
    .A2_N(\u_cpu._0507_ ),
    .B1(\u_cpu._0503_ ),
    .B2(\u_cpu.counter[19] ),
    .X(\u_cpu._0010_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1055_  (.A(\u_cpu.counter[20] ),
    .B(\u_cpu._0505_ ),
    .C(\u_cpu._0507_ ),
    .X(\u_cpu._0508_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu._1056_  (.A1(\u_cpu._0505_ ),
    .A2(\u_cpu._0507_ ),
    .B1(\u_cpu.counter[20] ),
    .Y(\u_cpu._0509_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._1057_  (.A(\u_cpu._0508_ ),
    .B(\u_cpu._0509_ ),
    .Y(\u_cpu._0012_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu._1058_  (.A(\u_cpu.counter[19] ),
    .B(\u_cpu.counter[18] ),
    .C(\u_cpu._0500_ ),
    .D(\u_cpu._0501_ ),
    .X(\u_cpu._0510_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1059_  (.A(\u_cpu.counter[21] ),
    .B(\u_cpu.counter[20] ),
    .C(\u_cpu._0510_ ),
    .X(\u_cpu._0511_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu._1060_  (.A1(\u_cpu.counter[21] ),
    .A2(\u_cpu._0508_ ),
    .B1_N(\u_cpu._0511_ ),
    .X(\u_cpu._0013_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu._1061_  (.A(\u_cpu.counter[22] ),
    .B(\u_cpu._0511_ ),
    .X(\u_cpu._0014_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu._1062_  (.A(\u_cpu.counter[21] ),
    .B(\u_cpu.counter[20] ),
    .C(\u_cpu.counter[23] ),
    .D(\u_cpu.counter[22] ),
    .X(\u_cpu._0512_ ));
 sky130_fd_sc_hd__a41oi_2 \u_cpu._1063_  (.A1(\u_cpu.counter[21] ),
    .A2(\u_cpu.counter[20] ),
    .A3(\u_cpu.counter[22] ),
    .A4(\u_cpu._0510_ ),
    .B1(\u_cpu.counter[23] ),
    .Y(\u_cpu._0513_ ));
 sky130_fd_sc_hd__a21oi_2 \u_cpu._1064_  (.A1(\u_cpu._0510_ ),
    .A2(\u_cpu._0512_ ),
    .B1(\u_cpu._0513_ ),
    .Y(\u_cpu._0015_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._1065_  (.A(\u_cpu.counter[24] ),
    .B(\u_cpu._0505_ ),
    .C(\u_cpu._0507_ ),
    .D(\u_cpu._0512_ ),
    .Y(\u_cpu._0514_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu._1066_  (.A1(\u_cpu._0505_ ),
    .A2(\u_cpu._0507_ ),
    .A3(\u_cpu._0512_ ),
    .B1(\u_cpu.counter[24] ),
    .X(\u_cpu._0515_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._1067_  (.A(\u_cpu._0514_ ),
    .B(\u_cpu._0515_ ),
    .X(\u_cpu._0516_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1068_  (.A(\u_cpu._0516_ ),
    .X(\u_cpu._0016_ ));
 sky130_fd_sc_hd__a31o_2 \u_cpu._1069_  (.A1(\u_cpu.counter[24] ),
    .A2(\u_cpu._0510_ ),
    .A3(\u_cpu._0512_ ),
    .B1(\u_cpu.counter[25] ),
    .X(\u_cpu._0517_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1070_  (.A(\u_cpu.counter[24] ),
    .B(\u_cpu.counter[25] ),
    .C(\u_cpu._0512_ ),
    .X(\u_cpu._0518_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._1071_  (.A(\u_cpu._0500_ ),
    .B(\u_cpu._0501_ ),
    .C(\u_cpu._0507_ ),
    .D(\u_cpu._0518_ ),
    .Y(\u_cpu._0519_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1072_  (.A(\u_cpu._0519_ ),
    .X(\u_cpu._0520_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1073_  (.A(\u_cpu._0520_ ),
    .X(\u_cpu._0521_ ));
 sky130_fd_sc_hd__and2_2 \u_cpu._1074_  (.A(\u_cpu._0517_ ),
    .B(\u_cpu._0521_ ),
    .X(\u_cpu._0522_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1075_  (.A(\u_cpu._0522_ ),
    .X(\u_cpu._0017_ ));
 sky130_fd_sc_hd__inv_2 \u_cpu._1076_  (.A(\u_cpu.counter[0] ),
    .Y(\u_cpu._0000_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1077_  (.A0(\u_cpu.IMEM.rd[0] ),
    .A1(\u_cpu.M_AXI_WDATA[0] ),
    .S(\u_cpu._0521_ ),
    .X(\u_cpu._0523_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1078_  (.A(\u_cpu._0523_ ),
    .X(\u_cpu._0026_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1079_  (.A0(\u_cpu.IMEM.rd[1] ),
    .A1(\u_cpu.M_AXI_WDATA[1] ),
    .S(\u_cpu._0521_ ),
    .X(\u_cpu._0524_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1080_  (.A(\u_cpu._0524_ ),
    .X(\u_cpu._0027_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1081_  (.A0(\u_cpu.IMEM.rd[2] ),
    .A1(\u_cpu.M_AXI_WDATA[2] ),
    .S(\u_cpu._0521_ ),
    .X(\u_cpu._0525_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1082_  (.A(\u_cpu._0525_ ),
    .X(\u_cpu._0028_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1083_  (.A0(\u_cpu.IMEM.rd[3] ),
    .A1(\u_cpu.M_AXI_WDATA[3] ),
    .S(\u_cpu._0521_ ),
    .X(\u_cpu._0526_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1084_  (.A(\u_cpu._0526_ ),
    .X(\u_cpu._0029_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1085_  (.A0(\u_cpu.IMEM.rd[4] ),
    .A1(\u_cpu.M_AXI_WDATA[4] ),
    .S(\u_cpu._0521_ ),
    .X(\u_cpu._0527_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1086_  (.A(\u_cpu._0527_ ),
    .X(\u_cpu._0030_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1087_  (.A0(\u_cpu.IMEM.rd[5] ),
    .A1(\u_cpu.M_AXI_WDATA[5] ),
    .S(\u_cpu._0521_ ),
    .X(\u_cpu._0528_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1088_  (.A(\u_cpu._0528_ ),
    .X(\u_cpu._0031_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1089_  (.A0(\u_cpu.IMEM.rd[6] ),
    .A1(\u_cpu.M_AXI_WDATA[6] ),
    .S(\u_cpu._0521_ ),
    .X(\u_cpu._0529_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1090_  (.A(\u_cpu._0529_ ),
    .X(\u_cpu._0032_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1091_  (.A0(\u_cpu.IMEM.rd[7] ),
    .A1(\u_cpu.M_AXI_WDATA[7] ),
    .S(\u_cpu._0521_ ),
    .X(\u_cpu._0530_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1092_  (.A(\u_cpu._0530_ ),
    .X(\u_cpu._0033_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1093_  (.A(\u_cpu._0520_ ),
    .X(\u_cpu._0531_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1094_  (.A0(\u_cpu.IMEM.rd[8] ),
    .A1(\u_cpu.M_AXI_WDATA[8] ),
    .S(\u_cpu._0531_ ),
    .X(\u_cpu._0532_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1095_  (.A(\u_cpu._0532_ ),
    .X(\u_cpu._0034_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1096_  (.A0(\u_cpu.IMEM.rd[9] ),
    .A1(\u_cpu.M_AXI_WDATA[9] ),
    .S(\u_cpu._0531_ ),
    .X(\u_cpu._0533_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1097_  (.A(\u_cpu._0533_ ),
    .X(\u_cpu._0035_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1098_  (.A0(\u_cpu.IMEM.rd[10] ),
    .A1(\u_cpu.M_AXI_WDATA[10] ),
    .S(\u_cpu._0531_ ),
    .X(\u_cpu._0534_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1099_  (.A(\u_cpu._0534_ ),
    .X(\u_cpu._0036_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1100_  (.A0(\u_cpu.IMEM.rd[11] ),
    .A1(\u_cpu.M_AXI_WDATA[11] ),
    .S(\u_cpu._0531_ ),
    .X(\u_cpu._0535_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1101_  (.A(\u_cpu._0535_ ),
    .X(\u_cpu._0037_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1102_  (.A0(\u_cpu.IMEM.rd[12] ),
    .A1(\u_cpu.M_AXI_WDATA[12] ),
    .S(\u_cpu._0531_ ),
    .X(\u_cpu._0536_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1103_  (.A(\u_cpu._0536_ ),
    .X(\u_cpu._0038_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1104_  (.A0(\u_cpu.IMEM.rd[13] ),
    .A1(\u_cpu.M_AXI_WDATA[13] ),
    .S(\u_cpu._0531_ ),
    .X(\u_cpu._0537_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1105_  (.A(\u_cpu._0537_ ),
    .X(\u_cpu._0039_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1106_  (.A0(\u_cpu.IMEM.rd[14] ),
    .A1(\u_cpu.M_AXI_WDATA[14] ),
    .S(\u_cpu._0531_ ),
    .X(\u_cpu._0538_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1107_  (.A(\u_cpu._0538_ ),
    .X(\u_cpu._0040_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1108_  (.A0(\u_cpu.IMEM.rd[15] ),
    .A1(\u_cpu.M_AXI_WDATA[15] ),
    .S(\u_cpu._0531_ ),
    .X(\u_cpu._0539_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1109_  (.A(\u_cpu._0539_ ),
    .X(\u_cpu._0041_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1110_  (.A0(\u_cpu.IMEM.rd[16] ),
    .A1(\u_cpu.M_AXI_WDATA[16] ),
    .S(\u_cpu._0531_ ),
    .X(\u_cpu._0540_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1111_  (.A(\u_cpu._0540_ ),
    .X(\u_cpu._0042_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1112_  (.A0(\u_cpu.IMEM.rd[17] ),
    .A1(\u_cpu.M_AXI_WDATA[17] ),
    .S(\u_cpu._0531_ ),
    .X(\u_cpu._0541_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1113_  (.A(\u_cpu._0541_ ),
    .X(\u_cpu._0043_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1114_  (.A(\u_cpu._0520_ ),
    .X(\u_cpu._0542_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1115_  (.A0(\u_cpu.IMEM.rd[18] ),
    .A1(\u_cpu.M_AXI_WDATA[18] ),
    .S(\u_cpu._0542_ ),
    .X(\u_cpu._0543_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1116_  (.A(\u_cpu._0543_ ),
    .X(\u_cpu._0044_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1117_  (.A0(\u_cpu.IMEM.rd[19] ),
    .A1(\u_cpu.M_AXI_WDATA[19] ),
    .S(\u_cpu._0542_ ),
    .X(\u_cpu._0544_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1118_  (.A(\u_cpu._0544_ ),
    .X(\u_cpu._0045_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1119_  (.A0(\u_cpu.IMEM.rd[20] ),
    .A1(\u_cpu.M_AXI_WDATA[20] ),
    .S(\u_cpu._0542_ ),
    .X(\u_cpu._0545_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1120_  (.A(\u_cpu._0545_ ),
    .X(\u_cpu._0046_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1121_  (.A0(\u_cpu.IMEM.rd[21] ),
    .A1(\u_cpu.M_AXI_WDATA[21] ),
    .S(\u_cpu._0542_ ),
    .X(\u_cpu._0546_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1122_  (.A(\u_cpu._0546_ ),
    .X(\u_cpu._0047_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1123_  (.A0(\u_cpu.IMEM.rd[22] ),
    .A1(\u_cpu.M_AXI_WDATA[22] ),
    .S(\u_cpu._0542_ ),
    .X(\u_cpu._0547_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1124_  (.A(\u_cpu._0547_ ),
    .X(\u_cpu._0048_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1125_  (.A0(\u_cpu.IMEM.rd[23] ),
    .A1(\u_cpu.M_AXI_WDATA[23] ),
    .S(\u_cpu._0542_ ),
    .X(\u_cpu._0548_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1126_  (.A(\u_cpu._0548_ ),
    .X(\u_cpu._0049_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1127_  (.A0(\u_cpu.IMEM.rd[24] ),
    .A1(\u_cpu.M_AXI_WDATA[24] ),
    .S(\u_cpu._0542_ ),
    .X(\u_cpu._0549_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1128_  (.A(\u_cpu._0549_ ),
    .X(\u_cpu._0050_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1129_  (.A0(\u_cpu.IMEM.rd[25] ),
    .A1(\u_cpu.M_AXI_WDATA[25] ),
    .S(\u_cpu._0542_ ),
    .X(\u_cpu._0550_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1130_  (.A(\u_cpu._0550_ ),
    .X(\u_cpu._0051_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1131_  (.A0(\u_cpu.IMEM.rd[26] ),
    .A1(\u_cpu.M_AXI_WDATA[26] ),
    .S(\u_cpu._0542_ ),
    .X(\u_cpu._0551_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1132_  (.A(\u_cpu._0551_ ),
    .X(\u_cpu._0052_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1133_  (.A0(\u_cpu.IMEM.rd[27] ),
    .A1(\u_cpu.M_AXI_WDATA[27] ),
    .S(\u_cpu._0542_ ),
    .X(\u_cpu._0552_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1134_  (.A(\u_cpu._0552_ ),
    .X(\u_cpu._0053_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1135_  (.A(\u_cpu._0520_ ),
    .X(\u_cpu._0553_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1136_  (.A0(\u_cpu.IMEM.rd[28] ),
    .A1(\u_cpu.M_AXI_WDATA[28] ),
    .S(\u_cpu._0553_ ),
    .X(\u_cpu._0554_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1137_  (.A(\u_cpu._0554_ ),
    .X(\u_cpu._0054_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1138_  (.A0(\u_cpu.IMEM.rd[29] ),
    .A1(\u_cpu.M_AXI_WDATA[29] ),
    .S(\u_cpu._0553_ ),
    .X(\u_cpu._0555_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1139_  (.A(\u_cpu._0555_ ),
    .X(\u_cpu._0055_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1140_  (.A0(\u_cpu.IMEM.rd[30] ),
    .A1(\u_cpu.M_AXI_WDATA[30] ),
    .S(\u_cpu._0553_ ),
    .X(\u_cpu._0556_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1141_  (.A(\u_cpu._0556_ ),
    .X(\u_cpu._0056_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1142_  (.A0(\u_cpu.IMEM.rd[31] ),
    .A1(\u_cpu.M_AXI_WDATA[31] ),
    .S(\u_cpu._0553_ ),
    .X(\u_cpu._0557_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1143_  (.A(\u_cpu._0557_ ),
    .X(\u_cpu._0057_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1144_  (.A0(\u_cpu.M_AXI_AWADDR[0] ),
    .A1(\u_cpu.ALUResult_W_Reg[0] ),
    .S(\u_cpu._0553_ ),
    .X(\u_cpu._0558_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1145_  (.A(\u_cpu._0558_ ),
    .X(\u_cpu._0058_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1146_  (.A0(\u_cpu.M_AXI_AWADDR[1] ),
    .A1(\u_cpu.led[1] ),
    .S(\u_cpu._0553_ ),
    .X(\u_cpu._0559_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1147_  (.A(\u_cpu._0559_ ),
    .X(\u_cpu._0059_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1148_  (.A0(\u_cpu.M_AXI_AWADDR[2] ),
    .A1(\u_cpu.led[2] ),
    .S(\u_cpu._0553_ ),
    .X(\u_cpu._0560_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1149_  (.A(\u_cpu._0560_ ),
    .X(\u_cpu._0060_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1150_  (.A0(\u_cpu.M_AXI_AWADDR[3] ),
    .A1(\u_cpu.led[3] ),
    .S(\u_cpu._0553_ ),
    .X(\u_cpu._0561_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1151_  (.A(\u_cpu._0561_ ),
    .X(\u_cpu._0061_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1152_  (.A0(\u_cpu.M_AXI_AWADDR[4] ),
    .A1(\u_cpu.led[4] ),
    .S(\u_cpu._0553_ ),
    .X(\u_cpu._0562_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1153_  (.A(\u_cpu._0562_ ),
    .X(\u_cpu._0062_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1154_  (.A0(\u_cpu.M_AXI_AWADDR[5] ),
    .A1(\u_cpu.led[5] ),
    .S(\u_cpu._0553_ ),
    .X(\u_cpu._0563_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1155_  (.A(\u_cpu._0563_ ),
    .X(\u_cpu._0063_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1156_  (.A(\u_cpu._0520_ ),
    .X(\u_cpu._0564_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1157_  (.A0(\u_cpu.M_AXI_AWADDR[6] ),
    .A1(\u_cpu.led[6] ),
    .S(\u_cpu._0564_ ),
    .X(\u_cpu._0565_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1158_  (.A(\u_cpu._0565_ ),
    .X(\u_cpu._0064_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1159_  (.A0(\u_cpu.M_AXI_AWADDR[7] ),
    .A1(\u_cpu.led[7] ),
    .S(\u_cpu._0564_ ),
    .X(\u_cpu._0566_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1160_  (.A(\u_cpu._0566_ ),
    .X(\u_cpu._0065_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1161_  (.A0(\u_cpu.M_AXI_AWADDR[8] ),
    .A1(\u_cpu.led[8] ),
    .S(\u_cpu._0564_ ),
    .X(\u_cpu._0567_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1162_  (.A(\u_cpu._0567_ ),
    .X(\u_cpu._0066_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1163_  (.A0(\u_cpu.M_AXI_AWADDR[9] ),
    .A1(\u_cpu.led[9] ),
    .S(\u_cpu._0564_ ),
    .X(\u_cpu._0568_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1164_  (.A(\u_cpu._0568_ ),
    .X(\u_cpu._0067_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1165_  (.A0(\u_cpu.M_AXI_AWADDR[10] ),
    .A1(\u_cpu.ALUResult_W_Reg[10] ),
    .S(\u_cpu._0564_ ),
    .X(\u_cpu._0569_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1166_  (.A(\u_cpu._0569_ ),
    .X(\u_cpu._0068_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1167_  (.A0(\u_cpu.M_AXI_AWADDR[11] ),
    .A1(\u_cpu.ALUResult_W_Reg[11] ),
    .S(\u_cpu._0564_ ),
    .X(\u_cpu._0570_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1168_  (.A(\u_cpu._0570_ ),
    .X(\u_cpu._0069_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1169_  (.A0(\u_cpu.M_AXI_AWADDR[12] ),
    .A1(\u_cpu.ALUResult_W_Reg[12] ),
    .S(\u_cpu._0564_ ),
    .X(\u_cpu._0571_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1170_  (.A(\u_cpu._0571_ ),
    .X(\u_cpu._0070_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1171_  (.A0(\u_cpu.M_AXI_AWADDR[13] ),
    .A1(\u_cpu.ALUResult_W_Reg[13] ),
    .S(\u_cpu._0564_ ),
    .X(\u_cpu._0572_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1172_  (.A(\u_cpu._0572_ ),
    .X(\u_cpu._0071_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1173_  (.A0(\u_cpu.M_AXI_AWADDR[14] ),
    .A1(\u_cpu.ALUResult_W_Reg[14] ),
    .S(\u_cpu._0564_ ),
    .X(\u_cpu._0573_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1174_  (.A(\u_cpu._0573_ ),
    .X(\u_cpu._0072_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1175_  (.A0(\u_cpu.M_AXI_AWADDR[15] ),
    .A1(\u_cpu.ALUResult_W_Reg[15] ),
    .S(\u_cpu._0564_ ),
    .X(\u_cpu._0574_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1176_  (.A(\u_cpu._0574_ ),
    .X(\u_cpu._0073_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1177_  (.A(\u_cpu._0520_ ),
    .X(\u_cpu._0575_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1178_  (.A0(\u_cpu.M_AXI_AWADDR[16] ),
    .A1(\u_cpu.ALUResult_W_Reg[16] ),
    .S(\u_cpu._0575_ ),
    .X(\u_cpu._0576_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1179_  (.A(\u_cpu._0576_ ),
    .X(\u_cpu._0074_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1180_  (.A0(\u_cpu.M_AXI_AWADDR[17] ),
    .A1(\u_cpu.ALUResult_W_Reg[17] ),
    .S(\u_cpu._0575_ ),
    .X(\u_cpu._0577_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1181_  (.A(\u_cpu._0577_ ),
    .X(\u_cpu._0075_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1182_  (.A0(\u_cpu.M_AXI_AWADDR[18] ),
    .A1(\u_cpu.ALUResult_W_Reg[18] ),
    .S(\u_cpu._0575_ ),
    .X(\u_cpu._0578_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1183_  (.A(\u_cpu._0578_ ),
    .X(\u_cpu._0076_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1184_  (.A0(\u_cpu.M_AXI_AWADDR[19] ),
    .A1(\u_cpu.ALUResult_W_Reg[19] ),
    .S(\u_cpu._0575_ ),
    .X(\u_cpu._0579_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1185_  (.A(\u_cpu._0579_ ),
    .X(\u_cpu._0077_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1186_  (.A0(\u_cpu.M_AXI_AWADDR[20] ),
    .A1(\u_cpu.ALUResult_W_Reg[20] ),
    .S(\u_cpu._0575_ ),
    .X(\u_cpu._0580_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1187_  (.A(\u_cpu._0580_ ),
    .X(\u_cpu._0078_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1188_  (.A0(\u_cpu.M_AXI_AWADDR[21] ),
    .A1(\u_cpu.ALUResult_W_Reg[21] ),
    .S(\u_cpu._0575_ ),
    .X(\u_cpu._0581_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1189_  (.A(\u_cpu._0581_ ),
    .X(\u_cpu._0079_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1190_  (.A0(\u_cpu.M_AXI_AWADDR[22] ),
    .A1(\u_cpu.ALUResult_W_Reg[22] ),
    .S(\u_cpu._0575_ ),
    .X(\u_cpu._0582_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1191_  (.A(\u_cpu._0582_ ),
    .X(\u_cpu._0080_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1192_  (.A0(\u_cpu.M_AXI_AWADDR[23] ),
    .A1(\u_cpu.ALUResult_W_Reg[23] ),
    .S(\u_cpu._0575_ ),
    .X(\u_cpu._0583_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1193_  (.A(\u_cpu._0583_ ),
    .X(\u_cpu._0081_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1194_  (.A0(\u_cpu.M_AXI_AWADDR[24] ),
    .A1(\u_cpu.ALUResult_W_Reg[24] ),
    .S(\u_cpu._0575_ ),
    .X(\u_cpu._0584_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1195_  (.A(\u_cpu._0584_ ),
    .X(\u_cpu._0082_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1196_  (.A0(\u_cpu.M_AXI_AWADDR[25] ),
    .A1(\u_cpu.ALUResult_W_Reg[25] ),
    .S(\u_cpu._0575_ ),
    .X(\u_cpu._0585_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1197_  (.A(\u_cpu._0585_ ),
    .X(\u_cpu._0083_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1198_  (.A(\u_cpu._0520_ ),
    .X(\u_cpu._0586_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1199_  (.A0(\u_cpu.M_AXI_AWADDR[26] ),
    .A1(\u_cpu.ALUResult_W_Reg[26] ),
    .S(\u_cpu._0586_ ),
    .X(\u_cpu._0587_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1200_  (.A(\u_cpu._0587_ ),
    .X(\u_cpu._0084_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1201_  (.A0(\u_cpu.M_AXI_AWADDR[27] ),
    .A1(\u_cpu.ALUResult_W_Reg[27] ),
    .S(\u_cpu._0586_ ),
    .X(\u_cpu._0588_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1202_  (.A(\u_cpu._0588_ ),
    .X(\u_cpu._0085_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1203_  (.A0(\u_cpu.M_AXI_AWADDR[28] ),
    .A1(\u_cpu.ALUResult_W_Reg[28] ),
    .S(\u_cpu._0586_ ),
    .X(\u_cpu._0589_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1204_  (.A(\u_cpu._0589_ ),
    .X(\u_cpu._0086_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1205_  (.A0(\u_cpu.M_AXI_AWADDR[29] ),
    .A1(\u_cpu.ALUResult_W_Reg[29] ),
    .S(\u_cpu._0586_ ),
    .X(\u_cpu._0590_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1206_  (.A(\u_cpu._0590_ ),
    .X(\u_cpu._0087_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1207_  (.A0(\u_cpu.M_AXI_AWADDR[30] ),
    .A1(\u_cpu.ALUResult_W_Reg[30] ),
    .S(\u_cpu._0586_ ),
    .X(\u_cpu._0591_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1208_  (.A(\u_cpu._0591_ ),
    .X(\u_cpu._0088_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1209_  (.A0(\u_cpu.M_AXI_AWADDR[31] ),
    .A1(\u_cpu.ALUResult_W_Reg[31] ),
    .S(\u_cpu._0586_ ),
    .X(\u_cpu._0592_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1210_  (.A(\u_cpu._0592_ ),
    .X(\u_cpu._0089_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1211_  (.A0(\u_cpu.ALU.ALUResult[0] ),
    .A1(\u_cpu.M_AXI_AWADDR[0] ),
    .S(\u_cpu._0586_ ),
    .X(\u_cpu._0593_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1212_  (.A(\u_cpu._0593_ ),
    .X(\u_cpu._0090_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1213_  (.A0(\u_cpu.ALU.ALUResult[1] ),
    .A1(\u_cpu.M_AXI_AWADDR[1] ),
    .S(\u_cpu._0586_ ),
    .X(\u_cpu._0594_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1214_  (.A(\u_cpu._0594_ ),
    .X(\u_cpu._0091_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1215_  (.A0(\u_cpu.ALU.ALUResult[2] ),
    .A1(\u_cpu.M_AXI_AWADDR[2] ),
    .S(\u_cpu._0586_ ),
    .X(\u_cpu._0595_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1216_  (.A(\u_cpu._0595_ ),
    .X(\u_cpu._0092_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1217_  (.A0(\u_cpu.ALU.ALUResult[3] ),
    .A1(\u_cpu.M_AXI_AWADDR[3] ),
    .S(\u_cpu._0586_ ),
    .X(\u_cpu._0596_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1218_  (.A(\u_cpu._0596_ ),
    .X(\u_cpu._0093_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1219_  (.A(\u_cpu._0520_ ),
    .X(\u_cpu._0597_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1220_  (.A0(\u_cpu.ALU.ALUResult[4] ),
    .A1(\u_cpu.M_AXI_AWADDR[4] ),
    .S(\u_cpu._0597_ ),
    .X(\u_cpu._0598_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1221_  (.A(\u_cpu._0598_ ),
    .X(\u_cpu._0094_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1222_  (.A0(\u_cpu.ALU.ALUResult[5] ),
    .A1(\u_cpu.M_AXI_AWADDR[5] ),
    .S(\u_cpu._0597_ ),
    .X(\u_cpu._0599_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1223_  (.A(\u_cpu._0599_ ),
    .X(\u_cpu._0095_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1224_  (.A0(\u_cpu.ALU.ALUResult[6] ),
    .A1(\u_cpu.M_AXI_AWADDR[6] ),
    .S(\u_cpu._0597_ ),
    .X(\u_cpu._0600_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1225_  (.A(\u_cpu._0600_ ),
    .X(\u_cpu._0096_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1226_  (.A0(\u_cpu.ALU.ALUResult[7] ),
    .A1(\u_cpu.M_AXI_AWADDR[7] ),
    .S(\u_cpu._0597_ ),
    .X(\u_cpu._0601_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1227_  (.A(\u_cpu._0601_ ),
    .X(\u_cpu._0097_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1228_  (.A0(\u_cpu.ALU.ALUResult[8] ),
    .A1(\u_cpu.M_AXI_AWADDR[8] ),
    .S(\u_cpu._0597_ ),
    .X(\u_cpu._0602_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1229_  (.A(\u_cpu._0602_ ),
    .X(\u_cpu._0098_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1230_  (.A0(\u_cpu.ALU.ALUResult[9] ),
    .A1(\u_cpu.M_AXI_AWADDR[9] ),
    .S(\u_cpu._0597_ ),
    .X(\u_cpu._0603_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1231_  (.A(\u_cpu._0603_ ),
    .X(\u_cpu._0099_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1232_  (.A0(\u_cpu.ALU.ALUResult[10] ),
    .A1(\u_cpu.M_AXI_AWADDR[10] ),
    .S(\u_cpu._0597_ ),
    .X(\u_cpu._0604_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1233_  (.A(\u_cpu._0604_ ),
    .X(\u_cpu._0100_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1234_  (.A0(\u_cpu.ALU.ALUResult[11] ),
    .A1(\u_cpu.M_AXI_AWADDR[11] ),
    .S(\u_cpu._0597_ ),
    .X(\u_cpu._0605_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1235_  (.A(\u_cpu._0605_ ),
    .X(\u_cpu._0101_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1236_  (.A0(\u_cpu.ALU.ALUResult[12] ),
    .A1(\u_cpu.M_AXI_AWADDR[12] ),
    .S(\u_cpu._0597_ ),
    .X(\u_cpu._0606_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1237_  (.A(\u_cpu._0606_ ),
    .X(\u_cpu._0102_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1238_  (.A0(\u_cpu.ALU.ALUResult[13] ),
    .A1(\u_cpu.M_AXI_AWADDR[13] ),
    .S(\u_cpu._0597_ ),
    .X(\u_cpu._0607_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1239_  (.A(\u_cpu._0607_ ),
    .X(\u_cpu._0103_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1240_  (.A(\u_cpu._0520_ ),
    .X(\u_cpu._0608_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1241_  (.A0(\u_cpu.ALU.ALUResult[14] ),
    .A1(\u_cpu.M_AXI_AWADDR[14] ),
    .S(\u_cpu._0608_ ),
    .X(\u_cpu._0609_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1242_  (.A(\u_cpu._0609_ ),
    .X(\u_cpu._0104_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1243_  (.A0(\u_cpu.ALU.ALUResult[15] ),
    .A1(\u_cpu.M_AXI_AWADDR[15] ),
    .S(\u_cpu._0608_ ),
    .X(\u_cpu._0610_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1244_  (.A(\u_cpu._0610_ ),
    .X(\u_cpu._0105_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1245_  (.A0(\u_cpu.ALU.ALUResult[16] ),
    .A1(\u_cpu.M_AXI_AWADDR[16] ),
    .S(\u_cpu._0608_ ),
    .X(\u_cpu._0611_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1246_  (.A(\u_cpu._0611_ ),
    .X(\u_cpu._0106_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1247_  (.A0(\u_cpu.ALU.ALUResult[17] ),
    .A1(\u_cpu.M_AXI_AWADDR[17] ),
    .S(\u_cpu._0608_ ),
    .X(\u_cpu._0612_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1248_  (.A(\u_cpu._0612_ ),
    .X(\u_cpu._0107_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1249_  (.A0(\u_cpu.ALU.ALUResult[18] ),
    .A1(\u_cpu.M_AXI_AWADDR[18] ),
    .S(\u_cpu._0608_ ),
    .X(\u_cpu._0613_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1250_  (.A(\u_cpu._0613_ ),
    .X(\u_cpu._0108_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1251_  (.A0(\u_cpu.ALU.ALUResult[19] ),
    .A1(\u_cpu.M_AXI_AWADDR[19] ),
    .S(\u_cpu._0608_ ),
    .X(\u_cpu._0614_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1252_  (.A(\u_cpu._0614_ ),
    .X(\u_cpu._0109_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1253_  (.A0(\u_cpu.ALU.ALUResult[20] ),
    .A1(\u_cpu.M_AXI_AWADDR[20] ),
    .S(\u_cpu._0608_ ),
    .X(\u_cpu._0615_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1254_  (.A(\u_cpu._0615_ ),
    .X(\u_cpu._0110_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1255_  (.A0(\u_cpu.ALU.ALUResult[21] ),
    .A1(\u_cpu.M_AXI_AWADDR[21] ),
    .S(\u_cpu._0608_ ),
    .X(\u_cpu._0616_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1256_  (.A(\u_cpu._0616_ ),
    .X(\u_cpu._0111_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1257_  (.A0(\u_cpu.ALU.ALUResult[22] ),
    .A1(\u_cpu.M_AXI_AWADDR[22] ),
    .S(\u_cpu._0608_ ),
    .X(\u_cpu._0617_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1258_  (.A(\u_cpu._0617_ ),
    .X(\u_cpu._0112_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1259_  (.A0(\u_cpu.ALU.ALUResult[23] ),
    .A1(\u_cpu.M_AXI_AWADDR[23] ),
    .S(\u_cpu._0608_ ),
    .X(\u_cpu._0618_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1260_  (.A(\u_cpu._0618_ ),
    .X(\u_cpu._0113_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1261_  (.A(\u_cpu._0519_ ),
    .X(\u_cpu._0619_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1262_  (.A0(\u_cpu.ALU.ALUResult[24] ),
    .A1(\u_cpu.M_AXI_AWADDR[24] ),
    .S(\u_cpu._0619_ ),
    .X(\u_cpu._0620_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1263_  (.A(\u_cpu._0620_ ),
    .X(\u_cpu._0114_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1264_  (.A0(\u_cpu.ALU.ALUResult[25] ),
    .A1(\u_cpu.M_AXI_AWADDR[25] ),
    .S(\u_cpu._0619_ ),
    .X(\u_cpu._0621_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1265_  (.A(\u_cpu._0621_ ),
    .X(\u_cpu._0115_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1266_  (.A0(\u_cpu.ALU.ALUResult[26] ),
    .A1(\u_cpu.M_AXI_AWADDR[26] ),
    .S(\u_cpu._0619_ ),
    .X(\u_cpu._0622_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1267_  (.A(\u_cpu._0622_ ),
    .X(\u_cpu._0116_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1268_  (.A0(\u_cpu.ALU.ALUResult[27] ),
    .A1(\u_cpu.M_AXI_AWADDR[27] ),
    .S(\u_cpu._0619_ ),
    .X(\u_cpu._0623_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1269_  (.A(\u_cpu._0623_ ),
    .X(\u_cpu._0117_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1270_  (.A0(\u_cpu.ALU.ALUResult[28] ),
    .A1(\u_cpu.M_AXI_AWADDR[28] ),
    .S(\u_cpu._0619_ ),
    .X(\u_cpu._0624_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1271_  (.A(\u_cpu._0624_ ),
    .X(\u_cpu._0118_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1272_  (.A0(\u_cpu.ALU.ALUResult[29] ),
    .A1(\u_cpu.M_AXI_AWADDR[29] ),
    .S(\u_cpu._0619_ ),
    .X(\u_cpu._0625_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1273_  (.A(\u_cpu._0625_ ),
    .X(\u_cpu._0119_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1274_  (.A0(\u_cpu.ALU.ALUResult[30] ),
    .A1(\u_cpu.M_AXI_AWADDR[30] ),
    .S(\u_cpu._0619_ ),
    .X(\u_cpu._0626_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1275_  (.A(\u_cpu._0626_ ),
    .X(\u_cpu._0120_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1276_  (.A0(\u_cpu.ALU.ALUResult[31] ),
    .A1(\u_cpu.M_AXI_AWADDR[31] ),
    .S(\u_cpu._0619_ ),
    .X(\u_cpu._0627_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1277_  (.A(\u_cpu._0627_ ),
    .X(\u_cpu._0121_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu._1278_  (.A(\u_cpu._0500_ ),
    .B(\u_cpu._0501_ ),
    .C(\u_cpu._0507_ ),
    .D(\u_cpu._0518_ ),
    .X(\u_cpu._0628_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1279_  (.A(\u_cpu._0628_ ),
    .X(\u_cpu._0629_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._1280_  (.A(\u_cpu.IMEM.a[2] ),
    .B(\u_cpu._0629_ ),
    .Y(\u_cpu._0630_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1281_  (.A(\u_cpu.IMEM.a[2] ),
    .B(\u_cpu._0510_ ),
    .C(\u_cpu._0518_ ),
    .X(\u_cpu._0631_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._1282_  (.A(\u_cpu._0630_ ),
    .B(\u_cpu._0631_ ),
    .Y(\u_cpu._0122_ ));
 sky130_fd_sc_hd__o22a_2 \u_cpu._1283_  (.A1(\u_cpu._0373_ ),
    .A2(\u_cpu._0521_ ),
    .B1(\u_cpu._0631_ ),
    .B2(\u_cpu.IMEM.a[3] ),
    .X(\u_cpu._0123_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1284_  (.A(\u_cpu.IMEM.a[3] ),
    .B(\u_cpu.IMEM.a[2] ),
    .C(\u_cpu._0629_ ),
    .X(\u_cpu._0632_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu._1285_  (.A(\u_cpu.IMEM.a[4] ),
    .B(\u_cpu._0632_ ),
    .X(\u_cpu._0124_ ));
 sky130_fd_sc_hd__o211a_2 \u_cpu._1286_  (.A1(\u_cpu._0370_ ),
    .A2(\u_cpu._0371_ ),
    .B1(\u_cpu._0629_ ),
    .C1(\u_cpu._0366_ ),
    .X(\u_cpu._0633_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu._1287_  (.A1(\u_cpu.IMEM.a[5] ),
    .A2(\u_cpu._0632_ ),
    .B1_N(\u_cpu._0633_ ),
    .X(\u_cpu._0125_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1288_  (.A(\u_cpu._0366_ ),
    .B(\u_cpu._0370_ ),
    .C(\u_cpu._0629_ ),
    .X(\u_cpu._0634_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu._1289_  (.A(\u_cpu.IMEM.a[6] ),
    .B(\u_cpu._0634_ ),
    .X(\u_cpu._0126_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1290_  (.A0(\u_cpu.IMEM.a[7] ),
    .A1(\u_cpu._0377_ ),
    .S(\u_cpu._0634_ ),
    .X(\u_cpu._0635_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1291_  (.A(\u_cpu._0635_ ),
    .X(\u_cpu._0127_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1292_  (.A(\u_cpu.IMEM.a[5] ),
    .B(\u_cpu.IMEM.a[4] ),
    .C(\u_cpu._0366_ ),
    .X(\u_cpu._0636_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1293_  (.A(\u_cpu._0375_ ),
    .B(\u_cpu._0629_ ),
    .C(\u_cpu._0636_ ),
    .X(\u_cpu._0637_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu._1294_  (.A(\u_cpu.IMEM.a[8] ),
    .B(\u_cpu._0637_ ),
    .X(\u_cpu._0128_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu._1295_  (.A1(\u_cpu._0386_ ),
    .A2(\u_cpu._0387_ ),
    .B1(\u_cpu._0637_ ),
    .X(\u_cpu._0638_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu._1296_  (.A1(\u_cpu.IMEM.a[9] ),
    .A2(\u_cpu._0637_ ),
    .B1_N(\u_cpu._0638_ ),
    .X(\u_cpu._0129_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._1297_  (.A(\u_cpu._0375_ ),
    .B(\u_cpu._0386_ ),
    .C(\u_cpu._0629_ ),
    .D(\u_cpu._0636_ ),
    .Y(\u_cpu._0639_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu._1298_  (.A(\u_cpu.IMEM.a[10] ),
    .B(\u_cpu._0639_ ),
    .Y(\u_cpu._0130_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._1299_  (.A(\u_cpu._0393_ ),
    .B(\u_cpu._0394_ ),
    .Y(\u_cpu._0640_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1300_  (.A0(\u_cpu._0640_ ),
    .A1(\u_cpu.IMEM.a[11] ),
    .S(\u_cpu._0639_ ),
    .X(\u_cpu._0641_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1301_  (.A(\u_cpu._0641_ ),
    .X(\u_cpu._0131_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._1302_  (.A(\u_cpu.IMEM.a[5] ),
    .B(\u_cpu.IMEM.a[4] ),
    .C(\u_cpu.IMEM.a[7] ),
    .D(\u_cpu.IMEM.a[6] ),
    .Y(\u_cpu._0642_ ));
 sky130_fd_sc_hd__or4_2 \u_cpu._1303_  (.A(\u_cpu._0373_ ),
    .B(\u_cpu._0383_ ),
    .C(\u_cpu._0398_ ),
    .D(\u_cpu._0642_ ),
    .X(\u_cpu._0643_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._1304_  (.A(\u_cpu._0619_ ),
    .B(\u_cpu._0643_ ),
    .Y(\u_cpu._0644_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu._1305_  (.A(\u_cpu.IMEM.a[12] ),
    .B(\u_cpu._0644_ ),
    .X(\u_cpu._0132_ ));
 sky130_fd_sc_hd__o21a_2 \u_cpu._1306_  (.A1(\u_cpu._0391_ ),
    .A2(\u_cpu._0392_ ),
    .B1(\u_cpu._0644_ ),
    .X(\u_cpu._0645_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu._1307_  (.A1(\u_cpu.IMEM.a[13] ),
    .A2(\u_cpu._0644_ ),
    .B1_N(\u_cpu._0645_ ),
    .X(\u_cpu._0133_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu._1308_  (.A(\u_cpu._0396_ ),
    .B(\u_cpu._0619_ ),
    .C(\u_cpu._0643_ ),
    .X(\u_cpu._0646_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu._1309_  (.A(\u_cpu.IMEM.a[14] ),
    .B(\u_cpu._0646_ ),
    .Y(\u_cpu._0134_ ));
 sky130_fd_sc_hd__nand2_2 \u_cpu._1310_  (.A(\u_cpu._0646_ ),
    .B(\u_cpu.IMEM.a[15] ),
    .Y(\u_cpu._0647_ ));
 sky130_fd_sc_hd__o31ai_2 \u_cpu._1311_  (.A1(\u_cpu._0381_ ),
    .A2(\u_cpu._0382_ ),
    .A3(\u_cpu._0646_ ),
    .B1(\u_cpu._0647_ ),
    .Y(\u_cpu._0135_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._1312_  (.A(\u_cpu.IMEM.a[11] ),
    .B(\u_cpu.IMEM.a[10] ),
    .C(\u_cpu.IMEM.a[13] ),
    .D(\u_cpu.IMEM.a[12] ),
    .Y(\u_cpu._0648_ ));
 sky130_fd_sc_hd__nor4_2 \u_cpu._1313_  (.A(\u_cpu._0373_ ),
    .B(\u_cpu._0383_ ),
    .C(\u_cpu._0642_ ),
    .D(\u_cpu._0648_ ),
    .Y(\u_cpu._0649_ ));
 sky130_fd_sc_hd__or3b_2 \u_cpu._1314_  (.A(\u_cpu._0389_ ),
    .B(\u_cpu._0520_ ),
    .C_N(\u_cpu._0649_ ),
    .X(\u_cpu._0650_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu._1315_  (.A(\u_cpu.IMEM.a[16] ),
    .B(\u_cpu._0650_ ),
    .Y(\u_cpu._0136_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1316_  (.A(\u_cpu.IMEM.a[15] ),
    .B(\u_cpu.IMEM.a[14] ),
    .C(\u_cpu._0649_ ),
    .X(\u_cpu._0651_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu._1317_  (.A(\u_cpu._0629_ ),
    .B(\u_cpu._0651_ ),
    .C(\u_cpu._0428_ ),
    .D(\u_cpu._0410_ ),
    .X(\u_cpu._0652_ ));
 sky130_fd_sc_hd__a21o_2 \u_cpu._1318_  (.A1(\u_cpu.IMEM.a[17] ),
    .A2(\u_cpu._0650_ ),
    .B1(\u_cpu._0652_ ),
    .X(\u_cpu._0137_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1319_  (.A(\u_cpu._0407_ ),
    .B(\u_cpu._0629_ ),
    .C(\u_cpu._0651_ ),
    .X(\u_cpu._0653_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu._1320_  (.A(\u_cpu.IMEM.a[18] ),
    .B(\u_cpu._0653_ ),
    .X(\u_cpu._0138_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1321_  (.A0(\u_cpu.IMEM.a[19] ),
    .A1(\u_cpu._0421_ ),
    .S(\u_cpu._0653_ ),
    .X(\u_cpu._0654_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1322_  (.A(\u_cpu._0654_ ),
    .X(\u_cpu._0139_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1323_  (.A(\u_cpu._0417_ ),
    .B(\u_cpu._0407_ ),
    .C(\u_cpu._0651_ ),
    .X(\u_cpu._0152_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu._1324_  (.A(\u_cpu._0505_ ),
    .B(\u_cpu._0507_ ),
    .C(\u_cpu._0518_ ),
    .D(\u_cpu._0152_ ),
    .X(\u_cpu._0153_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu._1325_  (.A(\u_cpu.IMEM.a[20] ),
    .B(\u_cpu._0153_ ),
    .X(\u_cpu._0140_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1326_  (.A0(\u_cpu.IMEM.a[21] ),
    .A1(\u_cpu._0420_ ),
    .S(\u_cpu._0153_ ),
    .X(\u_cpu._0154_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1327_  (.A(\u_cpu._0154_ ),
    .X(\u_cpu._0141_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1328_  (.A(\u_cpu._0416_ ),
    .B(\u_cpu._0628_ ),
    .C(\u_cpu._0152_ ),
    .X(\u_cpu._0155_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu._1329_  (.A(\u_cpu.IMEM.a[22] ),
    .B(\u_cpu._0155_ ),
    .X(\u_cpu._0142_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1330_  (.A0(\u_cpu.IMEM.a[23] ),
    .A1(\u_cpu._0413_ ),
    .S(\u_cpu._0155_ ),
    .X(\u_cpu._0156_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1331_  (.A(\u_cpu._0156_ ),
    .X(\u_cpu._0143_ ));
 sky130_fd_sc_hd__and4_2 \u_cpu._1332_  (.A(\u_cpu._0416_ ),
    .B(\u_cpu._0409_ ),
    .C(\u_cpu._0628_ ),
    .D(\u_cpu._0152_ ),
    .X(\u_cpu._0157_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu._1333_  (.A(\u_cpu.IMEM.a[24] ),
    .B(\u_cpu._0157_ ),
    .X(\u_cpu._0144_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1334_  (.A0(\u_cpu.IMEM.a[25] ),
    .A1(\u_cpu._0452_ ),
    .S(\u_cpu._0157_ ),
    .X(\u_cpu._0158_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1335_  (.A(\u_cpu._0158_ ),
    .X(\u_cpu._0145_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._1336_  (.A(\u_cpu._0382_ ),
    .B(\u_cpu._0417_ ),
    .C(\u_cpu._0407_ ),
    .D(\u_cpu._0649_ ),
    .Y(\u_cpu._0159_ ));
 sky130_fd_sc_hd__nand4_2 \u_cpu._1337_  (.A(\u_cpu.IMEM.a[25] ),
    .B(\u_cpu.IMEM.a[24] ),
    .C(\u_cpu._0416_ ),
    .D(\u_cpu._0409_ ),
    .Y(\u_cpu._0160_ ));
 sky130_fd_sc_hd__or3_2 \u_cpu._1338_  (.A(\u_cpu._0519_ ),
    .B(\u_cpu._0159_ ),
    .C(\u_cpu._0160_ ),
    .X(\u_cpu._0161_ ));
 sky130_fd_sc_hd__xnor2_2 \u_cpu._1339_  (.A(\u_cpu.IMEM.a[26] ),
    .B(\u_cpu._0161_ ),
    .Y(\u_cpu._0146_ ));
 sky130_fd_sc_hd__mux2_2 \u_cpu._1340_  (.A0(\u_cpu._0454_ ),
    .A1(\u_cpu.IMEM.a[27] ),
    .S(\u_cpu._0161_ ),
    .X(\u_cpu._0162_ ));
 sky130_fd_sc_hd__buf_1 \u_cpu._1341_  (.A(\u_cpu._0162_ ),
    .X(\u_cpu._0147_ ));
 sky130_fd_sc_hd__nor2_2 \u_cpu._1342_  (.A(\u_cpu._0159_ ),
    .B(\u_cpu._0160_ ),
    .Y(\u_cpu._0163_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1343_  (.A(\u_cpu.IMEM.a[27] ),
    .B(\u_cpu.IMEM.a[26] ),
    .C(\u_cpu._0163_ ),
    .X(\u_cpu._0164_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1344_  (.A(\u_cpu._0510_ ),
    .B(\u_cpu._0518_ ),
    .C(\u_cpu._0164_ ),
    .X(\u_cpu._0165_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu._1345_  (.A(\u_cpu.IMEM.a[28] ),
    .B(\u_cpu._0165_ ),
    .X(\u_cpu._0148_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu._1346_  (.A1(\u_cpu._0441_ ),
    .A2(\u_cpu._0442_ ),
    .B1(\u_cpu._0510_ ),
    .C1(\u_cpu._0518_ ),
    .D1(\u_cpu._0164_ ),
    .X(\u_cpu._0166_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu._1347_  (.A1(\u_cpu.IMEM.a[29] ),
    .A2(\u_cpu._0165_ ),
    .B1_N(\u_cpu._0166_ ),
    .X(\u_cpu._0149_ ));
 sky130_fd_sc_hd__and3_2 \u_cpu._1348_  (.A(\u_cpu._0442_ ),
    .B(\u_cpu._0629_ ),
    .C(\u_cpu._0164_ ),
    .X(\u_cpu._0167_ ));
 sky130_fd_sc_hd__xor2_2 \u_cpu._1349_  (.A(\u_cpu.IMEM.a[30] ),
    .B(\u_cpu._0167_ ),
    .X(\u_cpu._0150_ ));
 sky130_fd_sc_hd__o2111a_2 \u_cpu._1350_  (.A1(\u_cpu._0443_ ),
    .A2(\u_cpu._0444_ ),
    .B1(\u_cpu._0629_ ),
    .C1(\u_cpu._0164_ ),
    .D1(\u_cpu._0442_ ),
    .X(\u_cpu._0168_ ));
 sky130_fd_sc_hd__o21ba_2 \u_cpu._1351_  (.A1(\u_cpu.IMEM.a[31] ),
    .A2(\u_cpu._0167_ ),
    .B1_N(\u_cpu._0168_ ),
    .X(\u_cpu._0151_ ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1352_  (.CLK(clknet_leaf_66_wb_clk_i),
    .D(\u_cpu._0000_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[0] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1353_  (.CLK(clknet_leaf_66_wb_clk_i),
    .D(\u_cpu._0011_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[1] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1354_  (.CLK(clknet_leaf_66_wb_clk_i),
    .D(\u_cpu._0018_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[2] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1355_  (.CLK(clknet_leaf_65_wb_clk_i),
    .D(\u_cpu._0019_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[3] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1356_  (.CLK(clknet_leaf_66_wb_clk_i),
    .D(\u_cpu._0020_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[4] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1357_  (.CLK(clknet_leaf_65_wb_clk_i),
    .D(\u_cpu._0021_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[5] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1358_  (.CLK(clknet_leaf_65_wb_clk_i),
    .D(\u_cpu._0022_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[6] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1359_  (.CLK(clknet_leaf_61_wb_clk_i),
    .D(\u_cpu._0023_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[7] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1360_  (.CLK(clknet_leaf_61_wb_clk_i),
    .D(\u_cpu._0024_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[8] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1361_  (.CLK(clknet_leaf_61_wb_clk_i),
    .D(\u_cpu._0025_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[9] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1362_  (.CLK(clknet_leaf_61_wb_clk_i),
    .D(\u_cpu._0001_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[10] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1363_  (.CLK(clknet_leaf_61_wb_clk_i),
    .D(\u_cpu._0002_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[11] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1364_  (.CLK(clknet_leaf_61_wb_clk_i),
    .D(\u_cpu._0003_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[12] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1365_  (.CLK(clknet_leaf_61_wb_clk_i),
    .D(\u_cpu._0004_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[13] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1366_  (.CLK(clknet_leaf_61_wb_clk_i),
    .D(\u_cpu._0005_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[14] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1367_  (.CLK(clknet_leaf_61_wb_clk_i),
    .D(\u_cpu._0006_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[15] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1368_  (.CLK(clknet_leaf_61_wb_clk_i),
    .D(\u_cpu._0007_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[16] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1369_  (.CLK(clknet_leaf_62_wb_clk_i),
    .D(\u_cpu._0008_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[17] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1370_  (.CLK(clknet_leaf_62_wb_clk_i),
    .D(\u_cpu._0009_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[18] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1371_  (.CLK(clknet_leaf_65_wb_clk_i),
    .D(\u_cpu._0010_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[19] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1372_  (.CLK(clknet_leaf_65_wb_clk_i),
    .D(\u_cpu._0012_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[20] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1373_  (.CLK(clknet_leaf_65_wb_clk_i),
    .D(\u_cpu._0013_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[21] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1374_  (.CLK(clknet_leaf_65_wb_clk_i),
    .D(\u_cpu._0014_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[22] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1375_  (.CLK(clknet_leaf_65_wb_clk_i),
    .D(\u_cpu._0015_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[23] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1376_  (.CLK(clknet_leaf_65_wb_clk_i),
    .D(\u_cpu._0016_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[24] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1377_  (.CLK(clknet_leaf_64_wb_clk_i),
    .D(\u_cpu._0017_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.counter[25] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1378_  (.CLK(clknet_leaf_84_wb_clk_i),
    .D(\u_cpu._0026_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[0] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1379_  (.CLK(clknet_leaf_84_wb_clk_i),
    .D(\u_cpu._0027_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[1] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1380_  (.CLK(clknet_leaf_88_wb_clk_i),
    .D(\u_cpu._0028_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[2] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1381_  (.CLK(clknet_leaf_85_wb_clk_i),
    .D(\u_cpu._0029_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[3] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1382_  (.CLK(clknet_leaf_89_wb_clk_i),
    .D(\u_cpu._0030_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[4] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1383_  (.CLK(clknet_leaf_89_wb_clk_i),
    .D(\u_cpu._0031_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[5] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1384_  (.CLK(clknet_leaf_88_wb_clk_i),
    .D(\u_cpu._0032_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[6] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1385_  (.CLK(clknet_leaf_88_wb_clk_i),
    .D(\u_cpu._0033_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[7] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1386_  (.CLK(clknet_leaf_89_wb_clk_i),
    .D(\u_cpu._0034_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[8] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1387_  (.CLK(clknet_leaf_89_wb_clk_i),
    .D(\u_cpu._0035_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[9] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1388_  (.CLK(clknet_leaf_90_wb_clk_i),
    .D(\u_cpu._0036_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[10] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1389_  (.CLK(clknet_leaf_90_wb_clk_i),
    .D(\u_cpu._0037_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[11] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1390_  (.CLK(clknet_leaf_85_wb_clk_i),
    .D(\u_cpu._0038_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[12] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1391_  (.CLK(clknet_leaf_89_wb_clk_i),
    .D(\u_cpu._0039_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[13] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1392_  (.CLK(clknet_leaf_84_wb_clk_i),
    .D(\u_cpu._0040_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[14] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1393_  (.CLK(clknet_leaf_84_wb_clk_i),
    .D(\u_cpu._0041_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[15] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1394_  (.CLK(clknet_leaf_68_wb_clk_i),
    .D(\u_cpu._0042_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[16] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1395_  (.CLK(clknet_leaf_68_wb_clk_i),
    .D(\u_cpu._0043_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[17] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1396_  (.CLK(clknet_leaf_70_wb_clk_i),
    .D(\u_cpu._0044_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[18] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1397_  (.CLK(clknet_leaf_68_wb_clk_i),
    .D(\u_cpu._0045_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[19] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1398_  (.CLK(clknet_leaf_86_wb_clk_i),
    .D(\u_cpu._0046_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[20] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1399_  (.CLK(clknet_leaf_85_wb_clk_i),
    .D(\u_cpu._0047_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[21] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1400_  (.CLK(clknet_leaf_86_wb_clk_i),
    .D(\u_cpu._0048_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[22] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1401_  (.CLK(clknet_leaf_87_wb_clk_i),
    .D(\u_cpu._0049_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[23] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1402_  (.CLK(clknet_leaf_68_wb_clk_i),
    .D(\u_cpu._0050_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[24] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1403_  (.CLK(clknet_leaf_68_wb_clk_i),
    .D(\u_cpu._0051_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[25] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1404_  (.CLK(clknet_leaf_68_wb_clk_i),
    .D(\u_cpu._0052_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[26] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1405_  (.CLK(clknet_leaf_87_wb_clk_i),
    .D(\u_cpu._0053_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[27] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1406_  (.CLK(clknet_leaf_85_wb_clk_i),
    .D(\u_cpu._0054_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[28] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1407_  (.CLK(clknet_leaf_85_wb_clk_i),
    .D(\u_cpu._0055_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[29] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1408_  (.CLK(clknet_leaf_86_wb_clk_i),
    .D(\u_cpu._0056_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[30] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1409_  (.CLK(clknet_leaf_85_wb_clk_i),
    .D(\u_cpu._0057_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_WDATA[31] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1410_  (.CLK(clknet_leaf_20_wb_clk_i),
    .D(\u_cpu._0058_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1411_  (.CLK(clknet_leaf_20_wb_clk_i),
    .D(\u_cpu._0059_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.led[1] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1412_  (.CLK(clknet_leaf_17_wb_clk_i),
    .D(\u_cpu._0060_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.led[2] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1413_  (.CLK(clknet_leaf_19_wb_clk_i),
    .D(\u_cpu._0061_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.led[3] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1414_  (.CLK(clknet_leaf_21_wb_clk_i),
    .D(\u_cpu._0062_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.led[4] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1415_  (.CLK(clknet_leaf_20_wb_clk_i),
    .D(\u_cpu._0063_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.led[5] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1416_  (.CLK(clknet_leaf_17_wb_clk_i),
    .D(\u_cpu._0064_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.led[6] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1417_  (.CLK(clknet_leaf_17_wb_clk_i),
    .D(\u_cpu._0065_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.led[7] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1418_  (.CLK(clknet_leaf_17_wb_clk_i),
    .D(\u_cpu._0066_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.led[8] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1419_  (.CLK(clknet_leaf_19_wb_clk_i),
    .D(\u_cpu._0067_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.led[9] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1420_  (.CLK(clknet_leaf_22_wb_clk_i),
    .D(\u_cpu._0068_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[10] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1421_  (.CLK(clknet_leaf_20_wb_clk_i),
    .D(\u_cpu._0069_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[11] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1422_  (.CLK(clknet_leaf_19_wb_clk_i),
    .D(\u_cpu._0070_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[12] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1423_  (.CLK(clknet_leaf_19_wb_clk_i),
    .D(\u_cpu._0071_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[13] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1424_  (.CLK(clknet_leaf_22_wb_clk_i),
    .D(\u_cpu._0072_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[14] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1425_  (.CLK(clknet_leaf_22_wb_clk_i),
    .D(\u_cpu._0073_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[15] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1426_  (.CLK(clknet_leaf_23_wb_clk_i),
    .D(\u_cpu._0074_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[16] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1427_  (.CLK(clknet_leaf_22_wb_clk_i),
    .D(\u_cpu._0075_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[17] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1428_  (.CLK(clknet_leaf_24_wb_clk_i),
    .D(\u_cpu._0076_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[18] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1429_  (.CLK(clknet_leaf_24_wb_clk_i),
    .D(\u_cpu._0077_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[19] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1430_  (.CLK(clknet_leaf_22_wb_clk_i),
    .D(\u_cpu._0078_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[20] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1431_  (.CLK(clknet_leaf_22_wb_clk_i),
    .D(\u_cpu._0079_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[21] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1432_  (.CLK(clknet_leaf_23_wb_clk_i),
    .D(\u_cpu._0080_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[22] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1433_  (.CLK(clknet_leaf_23_wb_clk_i),
    .D(\u_cpu._0081_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[23] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1434_  (.CLK(clknet_leaf_23_wb_clk_i),
    .D(\u_cpu._0082_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[24] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1435_  (.CLK(clknet_leaf_23_wb_clk_i),
    .D(\u_cpu._0083_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[25] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1436_  (.CLK(clknet_leaf_25_wb_clk_i),
    .D(\u_cpu._0084_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[26] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1437_  (.CLK(clknet_leaf_25_wb_clk_i),
    .D(\u_cpu._0085_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[27] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1438_  (.CLK(clknet_leaf_23_wb_clk_i),
    .D(\u_cpu._0086_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[28] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1439_  (.CLK(clknet_leaf_24_wb_clk_i),
    .D(\u_cpu._0087_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[29] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1440_  (.CLK(clknet_leaf_25_wb_clk_i),
    .D(\u_cpu._0088_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[30] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1441_  (.CLK(clknet_leaf_25_wb_clk_i),
    .D(\u_cpu._0089_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.ALUResult_W_Reg[31] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1442_  (.CLK(clknet_leaf_25_wb_clk_i),
    .D(\u_cpu._0090_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[0] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1443_  (.CLK(clknet_leaf_17_wb_clk_i),
    .D(\u_cpu._0091_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[1] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1444_  (.CLK(clknet_leaf_17_wb_clk_i),
    .D(\u_cpu._0092_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[2] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1445_  (.CLK(clknet_leaf_19_wb_clk_i),
    .D(\u_cpu._0093_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[3] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1446_  (.CLK(clknet_leaf_19_wb_clk_i),
    .D(\u_cpu._0094_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[4] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1447_  (.CLK(clknet_leaf_20_wb_clk_i),
    .D(\u_cpu._0095_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[5] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1448_  (.CLK(clknet_leaf_17_wb_clk_i),
    .D(\u_cpu._0096_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[6] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1449_  (.CLK(clknet_leaf_17_wb_clk_i),
    .D(\u_cpu._0097_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[7] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1450_  (.CLK(clknet_leaf_16_wb_clk_i),
    .D(\u_cpu._0098_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[8] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1451_  (.CLK(clknet_leaf_18_wb_clk_i),
    .D(\u_cpu._0099_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[9] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1452_  (.CLK(clknet_leaf_22_wb_clk_i),
    .D(\u_cpu._0100_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[10] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1453_  (.CLK(clknet_leaf_21_wb_clk_i),
    .D(\u_cpu._0101_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[11] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1454_  (.CLK(clknet_leaf_19_wb_clk_i),
    .D(\u_cpu._0102_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[12] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1455_  (.CLK(clknet_leaf_18_wb_clk_i),
    .D(\u_cpu._0103_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[13] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1456_  (.CLK(clknet_leaf_22_wb_clk_i),
    .D(\u_cpu._0104_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[14] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1457_  (.CLK(clknet_leaf_24_wb_clk_i),
    .D(\u_cpu._0105_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[15] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1458_  (.CLK(clknet_leaf_23_wb_clk_i),
    .D(\u_cpu._0106_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[16] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1459_  (.CLK(clknet_leaf_23_wb_clk_i),
    .D(\u_cpu._0107_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[17] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1460_  (.CLK(clknet_leaf_24_wb_clk_i),
    .D(\u_cpu._0108_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[18] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1461_  (.CLK(clknet_leaf_24_wb_clk_i),
    .D(\u_cpu._0109_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[19] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1462_  (.CLK(clknet_leaf_22_wb_clk_i),
    .D(\u_cpu._0110_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[20] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1463_  (.CLK(clknet_leaf_23_wb_clk_i),
    .D(\u_cpu._0111_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[21] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1464_  (.CLK(clknet_leaf_25_wb_clk_i),
    .D(\u_cpu._0112_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[22] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1465_  (.CLK(clknet_leaf_24_wb_clk_i),
    .D(\u_cpu._0113_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[23] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1466_  (.CLK(clknet_leaf_25_wb_clk_i),
    .D(\u_cpu._0114_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[24] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1467_  (.CLK(clknet_leaf_25_wb_clk_i),
    .D(\u_cpu._0115_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[25] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1468_  (.CLK(clknet_leaf_25_wb_clk_i),
    .D(\u_cpu._0116_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[26] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1469_  (.CLK(clknet_leaf_25_wb_clk_i),
    .D(\u_cpu._0117_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[27] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1470_  (.CLK(clknet_leaf_23_wb_clk_i),
    .D(\u_cpu._0118_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[28] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1471_  (.CLK(clknet_leaf_26_wb_clk_i),
    .D(\u_cpu._0119_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[29] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1472_  (.CLK(clknet_leaf_26_wb_clk_i),
    .D(\u_cpu._0120_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[30] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1473_  (.CLK(clknet_leaf_25_wb_clk_i),
    .D(\u_cpu._0121_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.M_AXI_AWADDR[31] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1474_  (.CLK(clknet_leaf_66_wb_clk_i),
    .D(\u_cpu._0122_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[2] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1475_  (.CLK(clknet_leaf_66_wb_clk_i),
    .D(\u_cpu._0123_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[3] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1476_  (.CLK(clknet_leaf_66_wb_clk_i),
    .D(\u_cpu._0124_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[4] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1477_  (.CLK(clknet_leaf_66_wb_clk_i),
    .D(\u_cpu._0125_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[5] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1478_  (.CLK(clknet_leaf_67_wb_clk_i),
    .D(\u_cpu._0126_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[6] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1479_  (.CLK(clknet_leaf_67_wb_clk_i),
    .D(\u_cpu._0127_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[7] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1480_  (.CLK(clknet_leaf_67_wb_clk_i),
    .D(\u_cpu._0128_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[8] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1481_  (.CLK(clknet_leaf_67_wb_clk_i),
    .D(\u_cpu._0129_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[9] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1482_  (.CLK(clknet_leaf_66_wb_clk_i),
    .D(\u_cpu._0130_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[10] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1483_  (.CLK(clknet_leaf_66_wb_clk_i),
    .D(\u_cpu._0131_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[11] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1484_  (.CLK(clknet_leaf_65_wb_clk_i),
    .D(\u_cpu._0132_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[12] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1485_  (.CLK(clknet_leaf_64_wb_clk_i),
    .D(\u_cpu._0133_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[13] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1486_  (.CLK(clknet_leaf_67_wb_clk_i),
    .D(\u_cpu._0134_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[14] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1487_  (.CLK(clknet_leaf_67_wb_clk_i),
    .D(\u_cpu._0135_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[15] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1488_  (.CLK(clknet_leaf_67_wb_clk_i),
    .D(\u_cpu._0136_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[16] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1489_  (.CLK(clknet_leaf_67_wb_clk_i),
    .D(\u_cpu._0137_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[17] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1490_  (.CLK(clknet_leaf_67_wb_clk_i),
    .D(\u_cpu._0138_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[18] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1491_  (.CLK(clknet_leaf_64_wb_clk_i),
    .D(\u_cpu._0139_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[19] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1492_  (.CLK(clknet_leaf_64_wb_clk_i),
    .D(\u_cpu._0140_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[20] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1493_  (.CLK(clknet_leaf_64_wb_clk_i),
    .D(\u_cpu._0141_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[21] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1494_  (.CLK(clknet_leaf_67_wb_clk_i),
    .D(\u_cpu._0142_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[22] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1495_  (.CLK(clknet_leaf_67_wb_clk_i),
    .D(\u_cpu._0143_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[23] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1496_  (.CLK(clknet_leaf_64_wb_clk_i),
    .D(\u_cpu._0144_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[24] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1497_  (.CLK(clknet_leaf_64_wb_clk_i),
    .D(\u_cpu._0145_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[25] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1498_  (.CLK(clknet_leaf_63_wb_clk_i),
    .D(\u_cpu._0146_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[26] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1499_  (.CLK(clknet_leaf_64_wb_clk_i),
    .D(\u_cpu._0147_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[27] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1500_  (.CLK(clknet_leaf_62_wb_clk_i),
    .D(\u_cpu._0148_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[28] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1501_  (.CLK(clknet_leaf_64_wb_clk_i),
    .D(\u_cpu._0149_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[29] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1502_  (.CLK(clknet_leaf_63_wb_clk_i),
    .D(\u_cpu._0150_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[30] ));
 sky130_fd_sc_hd__dfrtp_2 \u_cpu._1503_  (.CLK(clknet_leaf_62_wb_clk_i),
    .D(\u_cpu._0151_ ),
    .RESET_B(\u_cpu.rst_n ),
    .Q(\u_cpu.IMEM.a[31] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1513_  (.LO(\u_cpu.REG_FILE.a3[0] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1514_  (.LO(\u_cpu.REG_FILE.a3[1] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1515_  (.LO(\u_cpu.REG_FILE.a3[2] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1516_  (.LO(\u_cpu.REG_FILE.a3[3] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1517_  (.LO(\u_cpu.REG_FILE.a3[4] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1518_  (.LO(\u_cpu.REG_FILE.wd3[0] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1519_  (.LO(\u_cpu.REG_FILE.wd3[1] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1520_  (.LO(\u_cpu.REG_FILE.wd3[2] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1521_  (.LO(\u_cpu.REG_FILE.wd3[3] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1522_  (.LO(\u_cpu.REG_FILE.wd3[4] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1523_  (.LO(\u_cpu.REG_FILE.wd3[5] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1524_  (.LO(\u_cpu.REG_FILE.wd3[6] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1525_  (.LO(\u_cpu.REG_FILE.wd3[7] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1526_  (.LO(\u_cpu.REG_FILE.wd3[8] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1527_  (.LO(\u_cpu.REG_FILE.wd3[9] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1528_  (.LO(\u_cpu.REG_FILE.wd3[10] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1529_  (.LO(\u_cpu.REG_FILE.wd3[11] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1530_  (.LO(\u_cpu.REG_FILE.wd3[12] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1531_  (.LO(\u_cpu.REG_FILE.wd3[13] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1532_  (.LO(\u_cpu.REG_FILE.wd3[14] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1533_  (.LO(\u_cpu.REG_FILE.wd3[15] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1534_  (.LO(\u_cpu.REG_FILE.wd3[16] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1535_  (.LO(\u_cpu.REG_FILE.wd3[17] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1536_  (.LO(\u_cpu.REG_FILE.wd3[18] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1537_  (.LO(\u_cpu.REG_FILE.wd3[19] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1538_  (.LO(\u_cpu.REG_FILE.wd3[20] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1539_  (.LO(\u_cpu.REG_FILE.wd3[21] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1540_  (.LO(\u_cpu.REG_FILE.wd3[22] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1541_  (.LO(\u_cpu.REG_FILE.wd3[23] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1542_  (.LO(\u_cpu.REG_FILE.wd3[24] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1543_  (.LO(\u_cpu.REG_FILE.wd3[25] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1544_  (.LO(\u_cpu.REG_FILE.wd3[26] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1545_  (.LO(\u_cpu.REG_FILE.wd3[27] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1546_  (.LO(\u_cpu.REG_FILE.wd3[28] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1547_  (.LO(\u_cpu.REG_FILE.wd3[29] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1548_  (.LO(\u_cpu.REG_FILE.wd3[30] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1549_  (.LO(\u_cpu.REG_FILE.wd3[31] ));
 sky130_fd_sc_hd__conb_1 \u_cpu._1550_  (.LO(\u_cpu.REG_FILE.we3 ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__decap_3 PHY_572 ();
 sky130_fd_sc_hd__decap_3 PHY_573 ();
 sky130_fd_sc_hd__decap_3 PHY_574 ();
 sky130_fd_sc_hd__decap_3 PHY_575 ();
 sky130_fd_sc_hd__decap_3 PHY_576 ();
 sky130_fd_sc_hd__decap_3 PHY_577 ();
 sky130_fd_sc_hd__decap_3 PHY_578 ();
 sky130_fd_sc_hd__decap_3 PHY_579 ();
 sky130_fd_sc_hd__decap_3 PHY_580 ();
 sky130_fd_sc_hd__decap_3 PHY_581 ();
 sky130_fd_sc_hd__decap_3 PHY_582 ();
 sky130_fd_sc_hd__decap_3 PHY_583 ();
 sky130_fd_sc_hd__decap_3 PHY_584 ();
 sky130_fd_sc_hd__decap_3 PHY_585 ();
 sky130_fd_sc_hd__decap_3 PHY_586 ();
 sky130_fd_sc_hd__decap_3 PHY_587 ();
 sky130_fd_sc_hd__decap_3 PHY_588 ();
 sky130_fd_sc_hd__decap_3 PHY_589 ();
 sky130_fd_sc_hd__decap_3 PHY_590 ();
 sky130_fd_sc_hd__decap_3 PHY_591 ();
 sky130_fd_sc_hd__decap_3 PHY_592 ();
 sky130_fd_sc_hd__decap_3 PHY_593 ();
 sky130_fd_sc_hd__decap_3 PHY_594 ();
 sky130_fd_sc_hd__decap_3 PHY_595 ();
 sky130_fd_sc_hd__decap_3 PHY_596 ();
 sky130_fd_sc_hd__decap_3 PHY_597 ();
 sky130_fd_sc_hd__decap_3 PHY_598 ();
 sky130_fd_sc_hd__decap_3 PHY_599 ();
 sky130_fd_sc_hd__decap_3 PHY_600 ();
 sky130_fd_sc_hd__decap_3 PHY_601 ();
 sky130_fd_sc_hd__decap_3 PHY_602 ();
 sky130_fd_sc_hd__decap_3 PHY_603 ();
 sky130_fd_sc_hd__decap_3 PHY_604 ();
 sky130_fd_sc_hd__decap_3 PHY_605 ();
 sky130_fd_sc_hd__decap_3 PHY_606 ();
 sky130_fd_sc_hd__decap_3 PHY_607 ();
 sky130_fd_sc_hd__decap_3 PHY_608 ();
 sky130_fd_sc_hd__decap_3 PHY_609 ();
 sky130_fd_sc_hd__decap_3 PHY_610 ();
 sky130_fd_sc_hd__decap_3 PHY_611 ();
 sky130_fd_sc_hd__decap_3 PHY_612 ();
 sky130_fd_sc_hd__decap_3 PHY_613 ();
 sky130_fd_sc_hd__decap_3 PHY_614 ();
 sky130_fd_sc_hd__decap_3 PHY_615 ();
 sky130_fd_sc_hd__decap_3 PHY_616 ();
 sky130_fd_sc_hd__decap_3 PHY_617 ();
 sky130_fd_sc_hd__decap_3 PHY_618 ();
 sky130_fd_sc_hd__decap_3 PHY_619 ();
 sky130_fd_sc_hd__decap_3 PHY_620 ();
 sky130_fd_sc_hd__decap_3 PHY_621 ();
 sky130_fd_sc_hd__decap_3 PHY_622 ();
 sky130_fd_sc_hd__decap_3 PHY_623 ();
 sky130_fd_sc_hd__decap_3 PHY_624 ();
 sky130_fd_sc_hd__decap_3 PHY_625 ();
 sky130_fd_sc_hd__decap_3 PHY_626 ();
 sky130_fd_sc_hd__decap_3 PHY_627 ();
 sky130_fd_sc_hd__decap_3 PHY_628 ();
 sky130_fd_sc_hd__decap_3 PHY_629 ();
 sky130_fd_sc_hd__decap_3 PHY_630 ();
 sky130_fd_sc_hd__decap_3 PHY_631 ();
 sky130_fd_sc_hd__decap_3 PHY_632 ();
 sky130_fd_sc_hd__decap_3 PHY_633 ();
 sky130_fd_sc_hd__decap_3 PHY_634 ();
 sky130_fd_sc_hd__decap_3 PHY_635 ();
 sky130_fd_sc_hd__decap_3 PHY_636 ();
 sky130_fd_sc_hd__decap_3 PHY_637 ();
 sky130_fd_sc_hd__decap_3 PHY_638 ();
 sky130_fd_sc_hd__decap_3 PHY_639 ();
 sky130_fd_sc_hd__decap_3 PHY_640 ();
 sky130_fd_sc_hd__decap_3 PHY_641 ();
 sky130_fd_sc_hd__decap_3 PHY_642 ();
 sky130_fd_sc_hd__decap_3 PHY_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11659 ();
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_37_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_39_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_40_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_41_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_42_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_43_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_44_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_45_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_46_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_47_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_48_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_49_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_50_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_51_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_52_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_53_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_54_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_55_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_56_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_57_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_58_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_59_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_60_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_61_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_62_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_63_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_64_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_65_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_66_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_67_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_68_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_69_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_70_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_71_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_72_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_73_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_74_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_75_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_76_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_77_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_78_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_79_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_80_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_81_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_82_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_83_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_84_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_85_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_86_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_87_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_88_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_89_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_90_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_91_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_92_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_93_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_94_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_95_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_96_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_97_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_98_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_99_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_100_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_101_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_102_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_103_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_104_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_105_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_106_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_107_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_108_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_109_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_110_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_111_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_112_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_113_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_114_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_115_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_116_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_117_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_118_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_119_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_120_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_121_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_122_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_123_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_124_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_125_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_126_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_127_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_128_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_129_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_7_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0__f_wb_clk_i (.A(clknet_3_0_0_wb_clk_i),
    .X(clknet_4_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1__f_wb_clk_i (.A(clknet_3_0_0_wb_clk_i),
    .X(clknet_4_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2__f_wb_clk_i (.A(clknet_3_1_0_wb_clk_i),
    .X(clknet_4_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3__f_wb_clk_i (.A(clknet_3_1_0_wb_clk_i),
    .X(clknet_4_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4__f_wb_clk_i (.A(clknet_3_2_0_wb_clk_i),
    .X(clknet_4_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5__f_wb_clk_i (.A(clknet_3_2_0_wb_clk_i),
    .X(clknet_4_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6__f_wb_clk_i (.A(clknet_3_3_0_wb_clk_i),
    .X(clknet_4_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7__f_wb_clk_i (.A(clknet_3_3_0_wb_clk_i),
    .X(clknet_4_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8__f_wb_clk_i (.A(clknet_3_4_0_wb_clk_i),
    .X(clknet_4_8__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9__f_wb_clk_i (.A(clknet_3_4_0_wb_clk_i),
    .X(clknet_4_9__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10__f_wb_clk_i (.A(clknet_3_5_0_wb_clk_i),
    .X(clknet_4_10__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11__f_wb_clk_i (.A(clknet_3_5_0_wb_clk_i),
    .X(clknet_4_11__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12__f_wb_clk_i (.A(clknet_3_6_0_wb_clk_i),
    .X(clknet_4_12__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13__f_wb_clk_i (.A(clknet_3_6_0_wb_clk_i),
    .X(clknet_4_13__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14__f_wb_clk_i (.A(clknet_3_7_0_wb_clk_i),
    .X(clknet_4_14__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15__f_wb_clk_i (.A(clknet_3_7_0_wb_clk_i),
    .X(clknet_4_15__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\u_cpu.ALU.ALUResult[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\u_cpu.ALU.ALUResult[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\u_cpu.ALU.Product_Wallace[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\u_cpu.ALU.SrcA[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\u_cpu.ALU.SrcA[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\u_cpu.ALU.SrcA[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\u_cpu.ALU.SrcA[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\u_cpu.ALU.SrcA[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\u_cpu.ALU.SrcA[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\u_cpu.ALU.SrcA[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\u_cpu.ALU.SrcA[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\u_cpu.ALU.SrcA[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\u_cpu.ALU.SrcA[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\u_cpu.ALU.SrcB[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\u_cpu.ALU.SrcB[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\u_cpu.ALU.SrcB[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(\u_cpu.ALU.SrcB[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\u_cpu.ALU.SrcB[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\u_cpu.ALU.SrcB[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\u_cpu.ALU.SrcB[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\u_cpu.ALU.SrcB[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(\u_cpu.ALU.SrcB[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(\u_cpu.ALU.SrcB[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(\u_cpu.ALU.u_wallace._0272_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(\u_cpu.ALU.u_wallace._1333_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(\u_cpu.ALU.u_wallace._4450_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(\u_cpu.ALU.u_wallace._4450_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(\u_cpu.ALU.u_wallace._4554_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(\u_cpu.ALU.u_wallace._4662_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(\u_cpu.IMEM._0042_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(\u_cpu.IMEM._0113_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(\u_cpu.IMEM._0158_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(\u_cpu.IMEM._0262_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(\u_cpu.IMEM._0315_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(\u_cpu.IMEM._0321_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(\u_cpu.IMEM._0321_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(\u_cpu.IMEM._0351_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(\u_cpu.IMEM._0407_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(\u_cpu.IMEM._0450_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(\u_cpu.IMEM._0633_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(\u_cpu.IMEM.rd[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(\u_cpu.REG_FILE._01031_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(\u_cpu.REG_FILE._01032_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(\u_cpu.REG_FILE._01060_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(\u_cpu.REG_FILE._01106_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(\u_cpu.REG_FILE._01106_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(\u_cpu.REG_FILE._01106_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(\u_cpu.REG_FILE._01120_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(\u_cpu.REG_FILE._01125_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(\u_cpu.REG_FILE._01148_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(\u_cpu.REG_FILE._01151_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(\u_cpu.REG_FILE._01258_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(\u_cpu.REG_FILE._01258_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(\u_cpu.REG_FILE._01258_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(\u_cpu.REG_FILE._01258_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(\u_cpu.REG_FILE._01305_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(\u_cpu.REG_FILE._01305_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(\u_cpu.REG_FILE._01305_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(\u_cpu.REG_FILE._01305_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(\u_cpu.REG_FILE._01340_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(\u_cpu.REG_FILE._01340_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(\u_cpu.REG_FILE._01340_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(\u_cpu.REG_FILE._01340_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(\u_cpu.REG_FILE._01382_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(\u_cpu.REG_FILE._01611_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(\u_cpu.REG_FILE._01712_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(\u_cpu.REG_FILE._01811_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(\u_cpu.REG_FILE._01863_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(\u_cpu.REG_FILE._01962_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(\u_cpu.REG_FILE._02062_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(\u_cpu.REG_FILE._02580_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(\u_cpu.REG_FILE._02721_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(\u_cpu.REG_FILE._02754_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(\u_cpu.REG_FILE._02754_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(\u_cpu.REG_FILE._02793_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(\u_cpu.REG_FILE._02816_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(\u_cpu.REG_FILE._02816_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(\u_cpu.REG_FILE._02832_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(\u_cpu.REG_FILE._02838_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(\u_cpu.REG_FILE._02838_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(\u_cpu.REG_FILE._02838_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(\u_cpu.REG_FILE._02838_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(\u_cpu.REG_FILE._02838_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(\u_cpu.REG_FILE._02859_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(\u_cpu.REG_FILE._02867_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(\u_cpu.REG_FILE._02880_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(\u_cpu.REG_FILE._02880_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(\u_cpu.REG_FILE._02931_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(\u_cpu.REG_FILE._02931_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(\u_cpu.REG_FILE._02931_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(\u_cpu.REG_FILE._02945_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(\u_cpu.REG_FILE._02953_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(\u_cpu.REG_FILE._02970_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(\u_cpu.REG_FILE._02970_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(\u_cpu.REG_FILE._02970_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(\u_cpu.REG_FILE._02970_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(\u_cpu.REG_FILE._02970_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(\u_cpu.REG_FILE._02983_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(\u_cpu.REG_FILE._02983_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(\u_cpu.REG_FILE._02983_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(\u_cpu.REG_FILE._02983_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(\u_cpu.REG_FILE._02983_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(\u_cpu.REG_FILE._02986_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(\u_cpu.REG_FILE._02986_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(\u_cpu.REG_FILE._03050_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(\u_cpu.REG_FILE._03050_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(\u_cpu.REG_FILE._03050_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(\u_cpu.REG_FILE._03050_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(\u_cpu.REG_FILE._03060_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(\u_cpu.REG_FILE._03143_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(\u_cpu.REG_FILE._03143_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(\u_cpu.REG_FILE._03201_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(\u_cpu.REG_FILE._03204_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(\u_cpu.REG_FILE._03351_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(\u_cpu.REG_FILE._03537_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(\u_cpu.REG_FILE._03697_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(\u_cpu.REG_FILE._03743_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(\u_cpu.REG_FILE._03743_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(\u_cpu.REG_FILE._03743_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(\u_cpu.REG_FILE._03743_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(\u_cpu.REG_FILE._03787_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(\u_cpu.REG_FILE._03879_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(\u_cpu.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(\u_cpu.rst_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(\u_cpu.rst_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(\u_cpu.rst_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(clknet_leaf_39_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(\u_cpu.ALU.ALUResult[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(\u_cpu.ALU.SrcA[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(\u_cpu.ALU.SrcA[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(\u_cpu.ALU.SrcA[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(\u_cpu.ALU.u_wallace._0578_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(\u_cpu.ALU.u_wallace._4698_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(\u_cpu.IMEM._0080_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(\u_cpu.IMEM._0167_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(\u_cpu.IMEM._0351_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(\u_cpu.REG_FILE._01029_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(\u_cpu.REG_FILE._01029_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(\u_cpu.REG_FILE._01029_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(\u_cpu.REG_FILE._01029_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(\u_cpu.REG_FILE._01032_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(\u_cpu.REG_FILE._01125_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(\u_cpu.REG_FILE._01125_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(\u_cpu.REG_FILE._01125_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(\u_cpu.REG_FILE._01148_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(\u_cpu.REG_FILE._01148_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(\u_cpu.REG_FILE._01148_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(\u_cpu.REG_FILE._01148_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(\u_cpu.REG_FILE._01148_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(\u_cpu.REG_FILE._01148_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(\u_cpu.REG_FILE._01148_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(\u_cpu.REG_FILE._01382_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(\u_cpu.REG_FILE._01382_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(\u_cpu.REG_FILE._01382_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(\u_cpu.REG_FILE._01550_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(\u_cpu.REG_FILE._01550_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(\u_cpu.REG_FILE._01553_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(\u_cpu.REG_FILE._01553_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(\u_cpu.REG_FILE._02788_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(\u_cpu.REG_FILE._02804_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(\u_cpu.REG_FILE._02826_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(\u_cpu.REG_FILE._02880_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(\u_cpu.REG_FILE._02880_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(\u_cpu.REG_FILE._02880_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(\u_cpu.REG_FILE._02970_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(\u_cpu.REG_FILE._03024_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(\u_cpu.REG_FILE._03125_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(\u_cpu.REG_FILE._03133_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(\u_cpu.REG_FILE._03133_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(\u_cpu.REG_FILE._03331_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(\u_cpu.REG_FILE._03331_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(\u_cpu.REG_FILE._03351_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(\u_cpu.REG_FILE._04283_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(\u_cpu.rst_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(\u_cpu.rst_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(\u_cpu.rst_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(\u_cpu.ALU.u_wallace._1070_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(\u_cpu.ALU.u_wallace._1070_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(\u_cpu.ALU.u_wallace._1070_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(\u_cpu.REG_FILE._01032_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(\u_cpu.REG_FILE._02853_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(\u_cpu.REG_FILE._02853_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(\u_cpu.REG_FILE._02986_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(\u_cpu.REG_FILE._02986_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(\u_cpu.rst_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(\u_cpu.rst_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(\u_cpu.rst_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(\u_cpu.REG_FILE._01032_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(\u_cpu.rst_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(\u_cpu.rst_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(\u_cpu.REG_FILE._01032_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(\u_cpu.rst_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(\u_cpu.rst_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(\u_cpu.rst_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(\u_cpu.REG_FILE._01032_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(\u_cpu.rst_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(\u_cpu.rst_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(\u_cpu.rst_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(\u_cpu.REG_FILE._01032_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(\u_cpu.REG_FILE._01032_ ));
endmodule
